`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QL+s4GDNDZ7Z3MXm3H+iAQdEkAcUlnKxsXQATs2uQrpUrsT4ifW1jaOw59WEB11k
kp0zatMh8sOdaYVF1oFgDf88iTJxR+6MTwMLULfj/F7cb0eVHrIfW172i/XexEie
h0qWQps99dU3lYFrLHyJzUGj9IcwEI3JMr83sdk02eSiIQgjfoAny+4KutLxoV7t
Vdv6Oml16IW4jhcz8AHZABBM4t694LjBGmXjkLO7Leqa8GK07UuuHOqwnZCdI9gp
6XNSbuZK44IWNsTOh32XRPgZkVZixSTTv68L2v2pq4uvaw82Mwewt+f+vuIPLz60
JWW97c3ZA7SiFDeDavTWwdvXoULaN1qk1Tl65Le86KU/rZ8+nqq9hmuNS0E2AWyn
ViuxhpVQT5Rb/I899H8mVig7IdRn0wqKJOeEXGVJD1DNB6uQdqn1OtkgFRRZdpyM
HhI5GWYRQJMNgVNc9mz/HWJBFZ6eV0XujvYXaojWwalhmv6XyiTFG/oV2YNoMFox
RUcTDMDKFF5sylmcARVZvRp9I47YDb5RvlwdQNsQBGmSh6RNP2sEGKPPxJJz46gX
5livBDnIzBsGs1e9Hqs3O9vthEJbfzaCJCvZ/fQnQynZAl9T73AtNBwyI23jxFjS
4w97vGnP6qD24C/dJn/zGW681EOMa0EuLoJgq0ITPXVn6vkAXxxWTrbyFqMI1J6T
KnubshztCmsUh1DkZXRW43eP+r0A8+oYWVFZjxw9IrgCVtD0urPRHIWH7v8f7mHa
iek8c5Ih3MW87NIOqf6fgpKx7pbU6C0OOq9Os3bs8iInQvWVfSBCarOOE/fWvu6R
TLmSVigWSThYqkFxIoQsb+Kbx8eH2fj71IYgDLeTVyw2qoCVUCI9KacF9bSLxRtb
XjWYFpA0d4fDzC/ATleNwlOUaGV4Vv+Rnfw07LoKyWn9wdWbqa+XiaJIXzNytHSF
xZ0Tw1Ye+lAD+OF2/JiuXIwF2cIxKKd/6eYEoc3eQH0BlKu/NaosBQLTuyZc8sVo
qwwElEwXC/VOoEN2sW9Xo6XwdfqIg+L3ZvFmUES7KoNapZwCwuJ6JxwfmBFu+AY4
xIElNw0MFz1iVWJRzNDjygP0p9rnIg8oh/MEJt0Qb/9uPkOG57khWCbfHBXlKO53
VkaB0BH407nxzsQAdGMn2gae6RE7uO003UoOsf+Er6bpglBvoFd4Jpi8kVMxwsYW
O/orZo1GMmsW0sBamSRsWBFDXmvbYChjQ+Vs9T5RdDsWElB7NSJxztU/51FYmn4M
WTfwTlvhXryGfRN05fo/g2rEBIWJNy5jN4xdTPKNzJn/8frrnU7ikSmuNqO4i/la
zIwFK3qa88SfpYDbBY3s5dXydyp/w1Jvi+sVDTxtvfQfx6ESthqk4JipHbnmdRZi
Dzkj80HMrAc+9LRs6rCK+3uQZiIGqzfeq283tWwa8lciYNUoGfgyT2rfm4RY7Hz0
HTWZcileiymYLI7ZOUQN4TJgf5qllDX/cQUclPs5DTel8qsDz+NZM2mI3zsUTZuw
GoaZSL3LHANNmLQiu9txkuBViXlbNpbDrirI3F8zxf8=
`protect END_PROTECTED
