`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oxQFCzHE8soNXubkM+8aHHmgz6IrA4GOvX7qpyX6i8uscEgDeVIA13Vev3uwW9g/
CKl0KHkzfKLReMm2sw8R43FMrv+uLVIh9DzoSPeTptQk17lkQaVzT83dRq/uCKkQ
vWuLmV4iKLmhbaecUOZEhyMPyWfAr3DlNPH+BJgn8FaO2Et08YvEE7Oq2+JhAQ1A
gGve12zTyvu4bBYV2CABlrfc6De0vLPg9dbDAn3JaAJF8U+MlZRGqw8b8H3ltMXn
eYvHSOQpno9CXIoNbOjLSy8v6Nv9BH2T8TwAmxKuK25dDpcqcmv5NOcnXVg62Apd
XCdRhNH8urxGY+YmGtP3oamgj0wcABe9lwpk0lARiDgEiYfQrzZe1cAPLfcAMu1B
pmlPWKcISg/6XiYTsQqkAChw3WhKs86aAjOuIBozXu9+aRf+aXMgAeo9NnvNuC1X
wziaStkKAfEPywPqwY446LNz6dqxr2O9u0l4yo/o/Pp9Ij8yOr8w379ba7/xpS39
p2K7k+d5hKG4mNPmzhp9AhL9ZRXIXGspzkhFOByDgMxFizGf7Q9qCBZkz5uExaAQ
D+HNzxR2wBYCg9KoKfd4VhU1gQLle2Yq/+YuEWlRNyPgKEp+nCrk/zYgGE8H/BSD
86x4qxhrUnyfPckkwh8sLkjKwldwH5xIkjWv7T+0hXihMeeuWg+pjnlp61F86ioR
wf4zl3p2GZSXmQbvPmqThH9FOcGxeE1M/rUthEyvdcTTQ/upeqnMXTu66jdjd3OS
TtQy5LbMxBEBPlD4Uiv3qd7/vR78QP4nkj02EYBcrHuRbjHwFjTdswgLvLtAofmx
sSnQh1id4rylAumJsiA7Z+GX27MPYQV2Je+aGdJ8/+FAoEZS7hrAMuxv5CGzede8
nDElPdqLAjkO8j929r91fq3e1n7O7lBDyVBzVkg369abHOkmJFYs8sUrykiy81ZN
/8uzrRZhX2d8WJfP36M+BX6zR91VowRZ5xdwiPuz2JMUEtsMUocTEFpxl8lqE5Yh
JXMVZDpN6Jr6zXIg71WzIPZaMAoFkeooptZkFg1xoMhUosmQo9xNmKCEm8AT7hsx
j5syWxRP/PLber16JWuyhwijKGoly3K2WulTGC7UxBg1x1JzN9f/MyEjqnpf2Ypk
NJM/lnP0K7cyNDZlHdMacaHQXUfABIHRnGG3s48XQfemfcLbWxR9gR06Zk5x2Q62
puPq0xSz2vDqIexPRrFUAwplZkCPo4f8sRiBad/gBxh5raFIriJpdwiq4YqjnKog
ktjBjX3xum9+jVnhxTG2AVnvw8T9edwzffm/a1ck8flbJXbU30rWZ4YsA2vjenxH
Q7fZdnZ8wvEXsKJ93vfXOMPurfOwSWt0XFRsILOPAIWiFEbpakUUNEw5uDgOHDvw
4JrORijlCC/w31MLAeJFFTqMcCxbpt6riFwiFSrk0h2Bo8MZd4TRa1CFGe6rdO0h
etsNjtRHt1QyRNmxDQgmBoM2lmFs+oRT8meCekWv3H+rCiV/HdgSfN3q99FC1RND
9JDPde5sCzKOb3TnnZdR6vfTWhlvX7vhcX2++85EBMngkdMhpwypqnO8vZO1i8jc
7lLB+EiG6McE1BhK3N7hakJ060ygv1yUti1HeyDj9CQ=
`protect END_PROTECTED
