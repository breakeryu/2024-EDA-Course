`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tA8AafLJ4oZ1PJXYlsQATbpviF7sunlU7ffZtmBX+h7bvVLmpWqGCVNVz1azpuHZ
m8+yCipt1BPcfpRe97wL/3XswyL1tJ0xxRFFyt3CXL60gwYOCBtGDz227wdzLJPO
SxNogKcvFchm83NHmB39ArOmlHh78bj0x4LOFrHXnJ9Su9bgNmQYZ0rTP6l1Tuqn
nzS44UnJq5/rDBGbTOPDx0YjMyhgRwvvox4mc/bDyGLHz6A9rIjezRi8ZhGa8BRS
nmU9pF7Gzp+T3Rf9zG/qdKfWJ/icZx/U4AShf6Df0/GrRG1KlXg0+JSyLXSojiVj
gO8mkoBORN5eIbbqh0FnmdBr+6YsXtIlkH7z/LpTWn47I7k/1i4lJy5BzqG2v3jV
zQ6FCckaGEvtyH2GM+kzk+ratYIDK3Eo/YjaL6bp3o1vNJN0pj/4VpquMSB7kHPe
MSFWV2rUuMKiqsSjs9QfaoZS+othzYSEKC/go1F77+do2T4AnB3d1M5XDGAIHB2L
0QSBQ5XWSzp133xGgNrlhfVeXFddXRrVRBAZTuboabvyHTJgH0oUFmY0642spn6H
2YzZIi6U9fWGylUd03JwDXWwTM9DryYUlfxI2JO/3buo+Q/3htMbn5WqqoFUslmn
xLDCyf6BHs2ID8I8DKSD3q/WPFzntJABhqQyfhUIshFPdMsWpdzVXOjQQB+wI9Rq
8eAVCuxalcb/zHkg+UfcSnH6o2e5mpuFxu8f+XzdiMKMtEmElw+aPRIkpGYKuMOh
HjT5ztZGkjcEyxlRcjxqwDbco4oIAXFp+E6HuiBeZxLsIna9QvcyhKIfWcVcME7R
rL72JT+uFTkjhg+01MLByEpA/UjBzh/XZ+3V1J63ul5oCBYaYf6spKMlYL9V4fzB
GbSq8B9gcJ1Ec2vgVtkaVeFxxTknBHbyeRbugEwxZzmiicAIcjyVKBgR5f5wuXvm
W5R9OBXLlSC0TKWNhy1TifqrjjUUcFC7urXXRAmB/W68OMkkm+3Ew0ff6gUZ4TLf
tYosgBn7FFiqyy2qFsB+4dYa27pCGEUZXgURbc6CUkOteMbv1BeARXxHcv1JAV8z
dqs2qbz/1nXt0vg0g9ww/zE19SUJWVvPsQl4hiIccf4bNpjHjug/2IsCyxXV2EZU
ifyyNAPE7SuUbF8PfqCnQlRCnq8TwanlE/yiNjQHp8Tp6dYeB5Omqi4CmmBCY7TO
/Am/UOl+q3EhirJfw2fVrNKaBGL0+Rugpe7Lo1mmMwzsmQK0f4D/47BnQZq7zBOh
HvnYBGfW24VhtDhL6pFV1QjO0DLOexojieVtGYiOV8B9IgTkEnpFIReW06dQLnjK
k0oGzX45tMauL+3eXJYoMYTaLtfLaqtb7yRQr7j8AVvce9Ym4gEshVIHkeAStOu7
+1MnFhuFY3zyppi/c/o7kh6caQ4srvymlToOWE4fxu7UfogqrEKm9/IrPGBSCNWt
SbkU+tTdjUsMjaw3kW1upAyGE7Hbh1+/xmMl2wj7j26ziW6QZQbCR+qdLwat3r5S
OAuILTv1Vrrr60ZRAp8WzKtHEwk6YMcC6H/V5Xe4zRXdhZyKYAzM/9+B3MeWMFDw
OG2xlBX6xkkGfIW02NNGbEHZDZByifKkyAhayuw2gi6Zm4V1Ap4PdidNwSVLfBH+
QFKMbdNSvJNKlmWlTTtaJd88ILr/9eV2PjV2yDzHHwT1xhjoRTqAphtAS+BLqZ96
rpmfhGCcfZV4hd5wnlOuho9rErDyWZ9XAZNaXlWqc+35kvH6oTa3W9dilBdlqlsk
BUM/ftkCdl/UYgCwBe313D1KZOHgpscBuCgtLssmIVHpKjoAYfGj383lH406WJdJ
7YJof75XpD1t0eQuNDftF/Z0fMQqV/EpziEujt8mNJs9ukID8Fpgc5iMFi+ZfuM3
P0H0H1c1261817j02iIzm5Upj5lU8/59uMN3FvYVwpn9Vc/3Gqmyw0B0MKEKUm/g
sSiRx6Hmfuez/d9GdDIl/bh/vqV/g/jlZs0sBe9jKQiwbVDG5hT7NNgMg+JJNWlr
T22F6taE7xms0b3YDagQOB6RG+HzmNnI0XztKiPJqCfhSZ6IpwEzVHZmRb4fcV1t
AXqohNSgulGLsnJ40A8I+whBF8Siwrais9GzwwaUIornyCnoWP/2OvHdhy3JBlBF
ZHPqCgKcZFjs64jt0U5djhgwx4egXmAjits2JakjLYoeNNy2dnWH/iZR5Lmi/Y/e
r4Oi0ROE3m8UHYe4xu9HVhIslCYo1/q70s5yRCIvm8BaBPrzNy9HIK658dH7pWvm
egrjsi7IOxg4s5XZC+jjXutDABL1FmHTdc+6ctkeqbgcTAPjLTKlO0kir+7uYJkp
2mPwDSL5YNMBDKfNgpitVoDd4J6wTTR9Emfz0ZrAYdurBHCGdTCgx8NNwLb4l57v
+QV+Rxi0JVpP0LNhNgQtMavXYP2jsJQ0J+CzX31m5DuoMMgj2npJ4ZYOolcS3gtf
Us80pm6NxykgyspgswFJMZ+g7t2OZ9fJTStz/i9f1oceW/Y6I1sHAGDsCoDLDubf
U4n3sUgiugj5hPyKNFVbkn/EdeF0GcGADHmu/Z9TEVzey07mmLqykmf3RC1lz0Qf
qHTfePKi4L7OSRnd/Mgk021ybQ+Ux4UH3wciyUzMlOwVNMiwAI4mZCI4zt00/Nma
JhJo7nb3OiR1qgb6rhnTNJqd0VzShzfx04eQ/erpylnYA/Ly+WT+8yMsP7J0yxoQ
B4LeYm2D4K1nR4Zp+M9EmNUyU2DvvB4RPsxZxvYPTeKPAxkHrJc4OEaokWCU96wj
BE6TYc6zOWPnOazZN+sHniHveSmP8IMRA08iWWHmn1en+DIqb7gL8wNUXva287Us
sbWNFGIp+23ZjI+xf+1RTrejDbd5IIckoAEkVDZxBMZUgI/NYOnE+GZeMvsSbhTs
fqyF/ro0duYyVciCVjt1DWveOr7c9ZbXcVCtZU90Kh/TdJsfr/D01fEMl5QIyNeQ
zw9kA9XfuePJUx0WjvOktFbczijgzvK5vnq4HYHIPninEr2YtMypGyOYKL7tu+BC
TEMxSbeDrmY2Rc/Qa9qMkdl1yyoAjjnG0tZ4WxZa9Shpx84UX8UAYmtEZdw9gYvG
UInutJtSpyhTa8/83rwpORUxfuyknY/DEWVJ5L1RMti0axhdwB2U6Gyp1an6HMv9
mKn9PzzljI/KYh2rtPKiL0pWzco9144p4XEkNzLNjXQGxlICIccnIjZ4DbLwlXTJ
PCgYgu42vBxRe6uwf8Fg7hnkepAQkzPzBxzIuvPvcxQpK8JnhGEThGuokGImw/eL
dNBpUCEHoroS/Pxk45w2K8lPtnHyRiu2psQDtg1HxDyb2QASk1H5GWloffNA2MN/
R6eg6zIYenGM/qGn0fGzju+HoQp/xnDL8546oWoyHdzAoe7CSDYgrxsKToIZEpSd
Z8NTjnFsdJHSzycwQ4xKKW1zA5RkAqJ7Y9kLD1KgTUU65Zez7DEiNeCqfwj5T4fo
JfHho035xqFajVH0IPFBCvmKfVfuWFlpcDP9TxbBVSSlUAWAYn91zJ08AeLJUUQf
TsGlLG0GRgTavz1u5uth+vflHNTpSk+t0HqtgyIHB/ZNfwcFhaGMLMU5/J9aZqo3
yHe/7arSCc0aCNchB+h6OI2sWL2LAeMs/fXSmoFoPTZZ6j3LiOtgPFJtzVA0eMQj
SYTyfNyuoAuABfu7vLHMow==
`protect END_PROTECTED
