`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sXThJlcHmoHoBA0AYxxUeTD4LjqMKZpbt9LhGMaQk/kONFSuYdUrN6PVZ0b9x/zG
c3TlYHcaIsrKd6WFJv6C8Js6sFpzFbKcOnJGTX2Lvy9R7jf0IFDf/x73hftzOQn/
PU2ZBzCuYWWLNDuuhlslv6jqX8gXNrnqRGMjplkYFAPyjYXWdk19ioMHugWEnAWF
`protect END_PROTECTED
