`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdy3pX8qXCae5RK30uHh+ETM//wuSMLcmdiKb5luWzgYyE+EIYzPaLy8v+wkIoxI
4KdtFYlT4K0B4r2tB+D5v9Ch3/t+rnVRZ7WDWUzl5JJ1nN5qDobXRYxVrAdXoeNp
F5GKU0iEBbxpSPeEdezFpFiwvi9/gPxXzJAVJVVJTodcB7Ja3LAglPBsKi9dTCxi
2nMz++kq+CJpGWs521D6v1d2qRcWq4d92QBT21KI9qB+o78Ot3p2UYMmkVsyODIQ
Ra1uX96JTMt8blwYWtDP3PlmNm718B3j+7YCcDBgwNTbp+xS9rFJRC1WDAdP1yDR
uodTCC7RCSmSyJfVEKYVt4Tp715tncDP+xhwFVjkh8y2vfpO/iAsJkABqopbxUBA
Mw85xFx4gn0BbPhCjEgb4Wrf/KSKzKVr+qf1lFlgn++0Rp12HAWap+O48S+VKtq5
cuMUWOIG8xkeuqcjzLNg/Fl5IfEBZXAh5EmrYyjYdI3qyzl39pg9rAlkC5j47Rlt
1p8OkueYnLSDhiZP06sNAiVWr1UfzrlcG0WIv4+UTugtUkloCl2/w8zf8C6EKZtx
AaTp4OcokarM9IMgyhGPVDk6KqvqdwpOtQnpN8FeFeQc3LAkxsjFSHvT1e3tdD5V
ADVa4IgD1P8VQdJHn9w/xxAu4pF9LWk1Z1VF048lu8AzmlywYMotF6bOzQzd4lJO
+i1cPcjRBz34MQqXyKs+sfixhRsIEVzWNVeznR/3jM4=
`protect END_PROTECTED
