`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/QCK21jTeA1l6n+cAvcXeNKGswNsf/4QF3n80+wL70T4TorPWC+klGyB/cjnOgR
AkKlhP6pudCnAt1VKoh//NJ3paCl/1xwDDigqV/6tP/3qgvxhLRUxg1Z4EZD9T1f
rcPwMNM87UJ5MumL0wtZZEV4B0Ol+Skn7zC0nWXaqTvTS8ZxPLbLPOEeDhau58A5
NoMMYXIuee395sq854gvf36vLlfTpdlRx2x+OvcMOoY8EPGb4tlvE2dhmG5vQUmb
QVKGMnBggmCYQv9rZAqhU8xShW2OhR7IJQCeUTMk0C2ko53OuUasIi8ZaKCZpqrg
MNtqSnJMcrlpaYzzQ+aYPSbkezjHqKphsqSbEz48dmqu1ZfPV1kiqyo8NHRuun6K
O8RCVhAGKW5eTljP/ThOzUZ03aqxyKc4jvOVQjR5JDSPu5/QEuifY4O/EUWd8Ahe
XD+KmhPM4RgR6ylg4roLzBxLw4KML1mYdZtxJWtwSiOylUqBQxvDBo9kMSWCpZDT
TaZYK3TBQPPwCScEEQn8hpWYDxyDaSi7D1pgGOA66tjuWfcwSoXx9gUG07+EzeZ4
c/9V+q0oTumIA+tVme/8OzCctv8AeVKHUB4f3VlfXxjbqsJt9YwG/oKGCrjth0xJ
xIzak6s5flXkcDYtKU8vq8yirUZkMt9pOaLyHHw6/PLQNu7pUqA5jqBk8jr+mbWC
3MwoG7C/RbHRt4P/2VlFIV2Zp4iYLgvM/gCBnBC3UaV3Q+s6AH4O0Yw5O/JJewE5
Lw7NLTeeGXUpg3ihAZ9RJwu7kMWPl3oFaR8pjEHAPsrA6UuKQxZWkd5ILTaMBUHy
`protect END_PROTECTED
