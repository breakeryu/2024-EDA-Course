`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jCUWjEnmZQ2kh6Y3c9G5qkew0momflaLXEZOSUwhPL5rryrSmY4byX37dXEKyrmW
GSEG6ObYxZpdTZadfbvWY0TnWlUgGWC2VOfwTOCBkZ6C9bNGy9tCOAZwIZWlAz2h
pGJNlFl7oPJ7C/7Vc0D5tn7GMKNjfsaAw9LI3kK5kZ4=
`protect END_PROTECTED
