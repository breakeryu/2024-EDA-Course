`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3VdNxp+SOxoDGjSvxQDjTBdxiiSGjaMvu+ekAXKC3L5EdFEKp+8xHyWuajq8eovI
V5CeLy9VpPj4ksgmG6u3R/keP5g+oFsKAut+b6pNzrbm9EbOD3Q7BcrjUqez0yTm
KkPVft2dPsVPZIuTNnz+rG0aUpxU4S6ydHPitA0JHHwf3QQn5XXIJ5zyQPLmXhrc
UmhawMXAHzADYp9OlqROQBAYzZHmZlDG35r8MCm1rMv/3PL1CrLOOe37fsqJk84H
5D+hpOIA8No5xpS/AhQ+i8jd2eZ4VcQWC+SB2Oa21vZ/VhCExr1oFTF7zWQWmT1k
qVahMT5hhqneP5a5X/Yk3pXZb7g0eamP68FgqLvpe/0ZhtUytzZObz60An56MM47
2nmkaGrCTqHN4zZ4Jop555fkaFGplWVnq28EFcGVrW1V7aDyPbbjA0g31qnoOSlm
hNQXR2OMYqHQBVu5WsLHc6+Hnt/c1NBVeMrD3VYZvpzriWDCKVUQruCVgsWmhNAU
9ZlBAl1xW2BIDmkZj84/AVPCM2/clbdNKK+pfJM/wekTFecQewJUaB4gLpfpv0GR
rkdcX1ahaPkvoUqML6/15uEJnoY4q0pPRSsfkCEckVnmuaPf7Xz5ReOH9+egEx+b
nOY2vkjoox9dbTxCBC7Op88fTGDo4TlYAXaL3CSAcmxdsbhY6KtlcdLcdTLXd8Nl
Br3GwLYAjUIrPe+ma7HGAo9Cw5skgMqOLwBSU7orypWdjDTvlzek7kOCh3zC1YAP
cL2Nv1rL0kdnHdqCOJEQNaow4fj3jbfwcc+q9iJ57Q8PQxOLK7iIZV0zk3WSi4xf
UcunX3hzNeVb9Brp29oibF7f0Mv0ao7pgzYQs2cBWtHfHgfO2bOlnQX2eNCJmUqK
RpvsnAJK+M29fWhfokxYS/CPp2HiXquP2AAs4NWf01jXVCN/XxufOA6GyfasMpg+
YSnwk+BtbQ1FhpB9B5uuBbVxgwNYSLjMKbCXMUSULwTHW8R8M8Wqlb5gPDVJu+z+
wDBZ+jSPcmiupNCVBuIFQkPC5rE4BIeVfHo/20T2cBYwAPho9Wtb89TlvypDA/+z
lre0XYzXQHoFag12j9xr1CBF/vZfjRR+8HcB5hgAZqjs1ASm+TlifMzodE3XyyRV
Nr08MAxbNrgq0e0leGPdqj5y6BUmdEMeFRhYi30UoRKA3+HCqbeOOLFLB3BuvHzh
V5ut+VsOJpZj1H/7zXGJ4g/o7RRYbqLGly0PUXYPhHg+L7E9h3NhTfHF73HYM9p/
1IJLiEln4/cA20lmXri05OP/hTmr+858+wr6cVIctNWBOAZDhSwjt2g8I4w2uMiV
8nE2stVAJBKZ+iZlm6SE7MRLmIkcv/GPXl7TyYBE3ZRGbUuesmi5PBGaePbcbGff
fDaiSEMZEv1k535mi2/YeNnM4kg8MD+YnBTJ7vD4RWjSonr+C2QgtMV1PbeKHJHd
maArVAhkmWNR261z5jK4eB5opZSlVGvrOY/ntK5/+BnhQPlXe+OvGy1OVEh6oH5O
yFqjEhby8srJ5aYpYma0rNu+WMqgxHnP86Xqtt93Sm4vPD5f6JNriL2iMfBNaBis
+/TVMbgluGrMtspx9zo5L+m2xSC6HAivLyQ1uNgzVJ4an/lQ2jjQctxCMwxcL2Ls
4PScnzokjhQYgRwL2xFAysB51LxCJcgCHH/O5X1wZQSjD3mq5Ywe/vPa0Ov2m9Wy
pVhBf9t+RP6ZdiPr5xZr6pZM1eO+iZAx/bJhhbUhcVgDay9ERrfFW8CR/fvzr2ne
CBVJeOVBkPARFRg3VTuBOcOc2SobEeOTdBcLjHa4iHlcfoDyXmKtdf7JFioB0ltw
JB4yU6Hif5Qk6RpYWwK+lw2qllwkmnz1iMuMKLQzclP4QGHQt5boqcjjR7dH0o/N
0Dc0/pM4JgTgCT8J+TwSoOY2QlR7UAH4bHWFhoiAW9aYiHbXMDh/qKtbJ1m7Z+tH
60G7pTJAZWVyTq10DJ9uB1zZx4F3MTDeZuu/fgt7GMt2Hn/Mh4aBXuwMceDhmVIq
1lsiIwf9RKQVnQEK5CZA3VEf1SHhWkLdufUNljoKR90YAMrZeZus0gP06HNx6Zk4
G2lbqio8xuhCLog85YLCYcImLegXR+dyR9Ooo6HJOlpTb6ixnLmvInwEXsVFILE/
nHsE1NhQBMLbNMcWEQYREwTvStCZvpJx5vyhntSaPDk=
`protect END_PROTECTED
