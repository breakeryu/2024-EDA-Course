`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XOOXDNwQZ0o55OA2OyTf17+2TObQx/QDte2IKXt33v4mZkk1iqkOrLSptpVm9hjS
Z+T6wTrJVd9P18JlcU8z8iSiwKdmdloLE26g4dAdmg0fXo/Ay7n6FYe7l+ZLnJzF
HpTtrvKZc9Wv7tW/ztGNaokVi121CY6o2gXoDgpWr/IZDL9r2DKNPzWdY+lv+gO9
eJ4CYQX/nXM5NGwfQzBb855yKMCCOk2mAPiGRT4RaC4c0tfuNu9hpQHrailkJtlv
U+jcnVbwupoaTzzpbcZRXBu8JRZVdY+FLEenjXzAj5D/Vp91tLm55DRUsAXVCt8u
ovT0VDmC0NdulSvgmuW3A2oOC0J4gK3YCDh0L/xWnvtMy378exct9pYNp3R3Qw0M
L4w+4zTf0wIUYIDt21vbyvZ/lSRkICNfTte0eFootaYJlDU+Y5KMARcNqixDKVoY
SXtEHR5CEaZ5uyYMjnLsdFVMWszQJXoTXWGyhtjUlNW9FfyEfcuuP5Wl6WMWDmvC
1Pm1ltErnRzxPojs7e6/9RNvxLXZAcdERSconudU7jRYpOwxY2WdXhpuVqYBH1hd
BuyzQJsgJi8GBtnVqZm1TVYTdJptgauCQGcVekZCCV7HbIigWg2Iz2lfC6ii3UBi
T5++YKfuOw0xYdFyJinFYFGloIpnFfULrjvnkK2a4kE3NvvQzNhyBlGzP4EVIXvD
f1PbgINmGgdE9oGi6GXZyHpEOj76xdHLbdJH+NoSEseMc2ZezE3xugz4N/qN4a3x
34N45mf7kqQwgJjtf78uzGeX9eeVuswfNDjE3jr7Ni3ThlJ2nFdHxiayggyvq8jZ
fD32zbiwwFBsMBExEuQFNQ==
`protect END_PROTECTED
