`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQnxKf2E+Qhmk/LlFymzNl50783eeYatp6tqdUgZNt0Ebzauvq491SLB699G+Tx2
2DiTfdoCFKP8NWxVOPkRJh1clP3c08a/vxkLksb1X9YVJNYwWXYIkOb2g2e065GY
yLNohVUFc3coaWseIeX6BcHCI0H4N8BpNBX8MPRves0CclMcsVzWjHJj4qS5jw4m
05MlLrkA9MYFK9d5zsfT93Vc8EXEcIQSRKhvu/oLj1QteE3nw6erVcRhNnNqL6pl
hxEQX0xuqRvi3zojRzs9mXuqjX1KkLk6ctoLuQojBtGVKWTF8oIselcHS9ee1Y0M
v1KWrZ+cIdqIJuihoO/YP59TCfhXjOjLQzfxpuY07D4JqvENc7+Jgh5qaW9umiB1
T65MQrETHdW+HLpW0cORoDgXrz851UmImXDuc+hbq5ShAe47cgWZDLs65E3l9Feq
wZZkEg5UDAEqhTUUEuVicBMlAd5H1V5slPbskB1BupKMuUSmU+CwaaiY2PxgMEJh
A6MaKj+eVa/Y2T/brOSRDJHTEk8MZOhjxSUxz8AFMcSUwDk1L7SUW/zPXzRlLSDv
8wa/IeCZPukgkfpYK+nGxdMsJFlqZ2YlxB5hXQyoQRb9ksoxevI2gsgGmZsuYkbB
NpGfLaBlsPyg4kdiQQlcJ6QiqHrMP8nYv1VZPQuxaUO9P2q0mCY32bkn4nSZUt8L
BmyucbyGoXrzMPSb58N80P/P3rsIu0PwKq3iI4amIhtcU6KC6wA9KUBJ/vBIoavL
vD2vD34S42AUks8v0h5972gQo2salqGgFpuUx7DibHFtQ6+zgAkMIEWtq00On850
fOhUTRXROvLRqIh7vZ1bb7FmR//GHeP619C6jzNlZBdzwQszdyRyWq18AO33j/xc
Zb1OrxlXlGHKV84lY1BKvXxsy5WY4kCA8aR8LU0+5HDBObJYYjST3xJKHHtL/O4u
PHzKco4UNd8HefE68lwe1S/YZ5NxGp6UFgmsaQyyESoCPyYR++YSb/rUe83wYnyn
zo+Q+pHgmsqh/865XnDARza+pnC7RtrixZXly66CijmA1s66M88vJwWm5yVOa7sf
z/4g1lDEamyeOu4zImQjgUW18tf0+ZkTCSYOw7BzokDsOiGlhdHTdwUlSXu+K6nU
AKFqfTPch4gET9KjvyFPytb6F4iOTwkbuv3y5tfBLWv5+6Z4OUx9F7dvkseYcUHo
xGbWAkmkORG4Av0ODHwBvioYVC687iyahHv1sDgrHofN5zcv0hQIlRudSot+mULs
T6J9I57/0CAIoq6cQK488vwSRQKpKy9SdWK/0m3WJtKEnhkHoQu9XhbA1UMln4k7
FYg16/QSJU46L87f2MHXlqi8scdjIv84Lf49NPgQVqslgdrEfGDzO5Z8Do4d/u//
ODhnoLfYtiFBj+BehXlHY/sbNLl65ojWSS12O0riz8PCRGnrGsoIg8skOqWPcmX2
kWgTV8buEv905v4L1RmuUT9KG/VVXB1a9pIFI/iqRGHtGKlMM4yunbqqMChpJSOa
pM3B8DofGMYUq2q8dpHdo0po20ufibL2bDySh54R1DzUtlijz94QqmqVO/fsSX8F
/+J2o0qIm8WJlROHYRqPacG0zqmIoV8z/F8xE/Ap44Kw2yurs0WZdQAn+WAg7OzP
a/Z/TanEyuXq/iBy63xZtwFhMhHzfVkwbfK8t4H3k6DNJke0KK8xJuEYKk1/Jz2E
tWkvEXyPRZJRtSNkd8ho6zOkhgC6HXiGdfFx22LIVvFIbLyZ32SeaMEUz0vqdkLL
soTH+VRIUpKdyfYHp7P9h2Te2Bo4nLhHr0BVdtnYadZvVUkeF+AgojDqFmcZH5jF
Qt8SybHyUHW1n95M6xwzpLCCU2DhdZRA/PvgNWR5v86wDxKFDANhR/Q2qG9AzIx8
wSo/WK2JLR0HeN4EZjcsE3gcfLDAZDXVo4apAK8S2a1cAllosUD3IVpVqR6GqUN3
VNpGAlB3j41xRq8RSkx4aZUkiQQnRKbm8IL0CDA6ZRRwsOvnrXSwQPcbj5wdeeIF
4MY4ILfNz76YcMHrsUUZaRRg84R7juq3ke1BIRikaIg/eHBtcr6lTwjoJ11z9Wps
1MKLq1kBQ/dso8+4L2gyljgNYVd/J5JFJ/wTovBlRpuGaLy0OojMmHPURRbgfTAu
M8vFB3OE4MgWl/WYero+a1irFlvMV8N/v8G31x9ynQ2Nr2HiB+pbQ+8Z+2Q1LnJ3
JZZermxPE0edieYxP3Dl0CykuM3NtqSaDj49ZToJ+1vhXzBlf75zz0efwfTg6oiJ
izojY6hfOti2mP3LueMcNiA72pMzFceLpWaYZy7mkrWIEKc0ITNbDXSVvpxSSWQo
lAV8k5XH8SMvUgdKhSb/7vcRwCqJZeE64wvadOO7tbS2pPTwRc3OIY17VD7J6d4f
cUV2R9TUwaazrfQ+bQTQkj+VSncxm3Bw7iu2IoLl+qIeER8tRrFEN+ywAgWv1qbf
oOyNjKUhYd6wmkXF3JwwqmxT/vc2HhNpBNOu3vBbpvxsFbvysyk4KM3cnuKZFo1c
YoPfkinrgbqEsoaBAntq10ROhXGhbedLMAE3rqXnDHGFIuJGr9Tg57G0IzSjWkBE
ejK90ZhtkacEec81Pz3yodMqUtT9yr5FCDavZHEEzimjnkDHlS9rUAcf4AGmXlbU
Q7xFGxK161woH1XdW1h2zsnZ7mX4X1c47R97D0jnDdfE3k3xZK2ctkJSqB9LwKxf
nfqego9p3XyDieWrgDqid8VUMP+xvE5mEYDAVWa97CnbDXbaHEOgTefzn8Fgdjro
a90fqrYn6579RwwzZu9HGk7YhPZIMFECU0mtnM48L0K/Yqq2elplnJ3KSeE7a/rX
b06FEKGoJ0FPH7kAOIe8OL9/m4BZ6x9tzlIRiqrfF8UVFeRpBOUd5skIO7Z9omRF
oN2kYdScXx78h3TLpWYT/3Z0boFfI+QT1nJMVdDrVypEs9LGprF4f5IYH3au/yYc
gK4Oe20QYzIPuIHJOFgjZvxlsBkGIiWIUG5EsKpC+qgA2b64XNAguKfWid1sF+j/
202MOmzppEsuKKkCR01ABFkkaU8QAkHPa3bRQt3F52rPts5Lc8gxXfe9vkJ4LCkv
ksW4pKAePccdJfiKF1pcIviywJfbE9xxfJm0XYq1Da+eBrF2Z+cP6gDSLz3MrnDZ
QwvhaAfymXD/SRJtwzpOxGnsKRm5bJtlfRh79LTBzURHh58Z08KKUjtvMYU9ldFq
2YptvKoSK9tdOfvBZ2fd9P+9mYz+9lzivys0FOQ7UdAyoSgAU/Q3gAKWOa1cFPAt
d7cZ7+pooMqfahWjtGJzTQZZRxYDX5wR2MSesRE9JMajfcrKBGBSe+G8ER5YQrY+
FL8VTV3KRqsI9wSCdDdxDO5FLFjQPGcaxoYQNbPnyF6XQG4LezDRXzu1zeBf2nwg
IAYXLQ86YaF3lkDrWo/nkFq4sQOiejN6xu54QgkpDPl7k8wScI43IHRDDxSrAIMg
0Ur3F29mvXUAIa9WxxM3derSi4Zaz4/souRz+lNYWTuommypl17QMTULu6DTGHnG
QGMTVDu+okxMyCpjc5TEor9i3XzXXEvqf+1AKAebx4Ipb68+claCf2hDgbz6aG+H
/M/ytwWnU1VWSWw2cTVO0A==
`protect END_PROTECTED
