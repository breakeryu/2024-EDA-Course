`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x6Hml5UnN0WH1Ie5WF9enhl2s3jHtOzSxB/Z5pAzIKkHwbqyu8J7LNivVEjZcHrP
HF7XDnKlp+ZUIZ7LqdeFGc1nb7B8veoRzuTxVWOoq+y1AES42dZzpISl76XDXov9
63I+H0Km0r16hF3Jo0DPSI5987cAryYwSkJB4aLc+P3JaKh0ENU69Z9bhvc0CKr+
Zlzg2oBq0GBT8b3t7cgGbUC/j6FItLfhLLhf/rDCxgFV2WpSEv0xq6P3ytCxnmDT
frqOqDPeoUhFiCLrCzLWIoOumo+r+eSjrcGSaP4gOh2pwsoTop1WT6BOdrAjmr3F
Ig8sU3unqD9Xsl+d+wVdyCA6GAxrt2CQHflR1M6VgoY+RGlP/Kjq4Ph3L/pz9G5p
tjgHlAvrZfJEnkSRd4FLSU0JnAnfbn102Bf+yGtFYq57cZCslxRT6jMUVYoQng6Z
xWboWmcVuqH2hjJ1PdcwYSEKpyqdj+aW3ckpn/JzJJDdKYDTIL04mTgTOGDVReKM
mNM/y9IWmDP0OK+lxhhy0lU6mKOghoBka82bolkEvaMijo3EfaS91+jmGkzYyy5M
AHCmSwIStl+6hmPrHLn02ukQn8R0lxHpK7jc40kwWa4c6U6Vv37ZZSpi7IcnsC27
pBOFptW315HWFMwe32vic13YN2hjHkibY+i9gahnCf5CGvAZH6/KbNcB93/PfHGk
25vVoHtDQP0D7PFy+zrIZGWFkjc2djm6lJGOaoGHQo8m8GthR+CmWgZ+L2w6RF4O
KX+H7xDWjbvl6404dEbOSl8bDhWm98lR0HAVFC/yp9X1hmia/pMXAVbVH80XaTEN
lmPebC0SCiGlgnrH1vAoEQ==
`protect END_PROTECTED
