`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uSb0Ue0hhvBJr/siaUKFDmGb8BZevOMAqYFOnumNHyOtuU/wn0ShtyvijRbF48Q
I04ikJP1qDcL3EixOc0zjPRl0mL1wF2kGR28Lj8DXb3Q7aFRA4eeaeqmESBhq8ea
313XCBMRKUcyuKgZ8QdmLpp/zG8bbIev6eGV+ah00sRbPfo9ZRefJ184d1u2sRUs
X+EmKvzcMF4BzHlB3VX40p9H83k3rmQpJCEN/LP4mEu3lW4rF1FtPkWA5La3E3Nx
XNnlZ3nmgCx1V4eYUWRrl4NGm1H9HMpFJgLHjP+rg8z1Cf13t8M5vuULDWwNCtHP
6aQ2tRdubVCzHeFSp1rdtE+cFkiwsEA0LrRKYm1+WnTuXzkIuISm7nooMq+AZs/3
/w9DjlTCT/xpILuE5CVB0D71eCqdjvsunpcScKAIEtEo4raUrsAwGAQT7HVLPW6y
SVyO/QfJrCoI8mywkqTTV38SazQMni5H8xCZGaX+W7/JxlzmXmdvqceuEHUeSEmg
8HRLoyMxbOwdOkNcZaqwGMHUfgZi4vXb/VTiBrwW9XnoFc8FeuWd57eFZvc6evnC
hWM3XjBOffEJaijUq0St48m6BKpR6F1QUZYZ9VZkN1+JYlAfbuiaoNRWZKU+rp4R
XH0HtRD4mi9n9iTV2gvPy0blQOVGMsFLQkybXoNXpdfYArlsfGbD9l2PEKZZgRjm
oaf5AN6cdglKQdg7dx9ARLWm1s9bGNRJCWEURwgCDZgzbHeuadYSn0MuUI7Jn3Sg
pjif1GAIB1wGjwlhYGn7kS7PRtvDkukWhlzNS7qw9lcBLWUPRaDwIrvN+K7yHig3
EctLllZca1bGumxK5UMuxzK2i3Ebzx5ScAxWtQVfgwo3FGVFpZ2xpwVzw+cvyfAV
4TjqqN2erKrtNie2Uqwb/yj+BYPFxcE4FxF2C5Mua+W9IL1oXSnUOudnzP/VdakC
SkWMLh+GhFs/l38BU+zrUFQfovcFEaa+SvIn6nN/QKKI4kYy5BBiTuT9Qrv3C95+
XTC2h8eCLiVNaDBlNkXVpIh3PBhDJTSGrrbJ0kMbYv3FnoQJFX3lPFz/OR5G/dvw
W0+/4ub7tYc/fnqKXuURWN+b22hdIOEEztalVJ1s1fhmRFY7GXAgBTIRywvJgp6i
HVNWy57ew73ws3IaeEg2O3MZr8i9I6Vv+3HhFMnGSpf7K+wrlvzF7eJdUbjdQBpo
Epan69CLe5ju69pSgNAdaMjnU0c8XhQ3iidbKdWtoJPfcbd6wXpPaZRJYVOQluIK
oDKeVfFy0TtzvfB//YJ8oUEA1IdQ8hg4DK039beZn+sfegx3TjoS2VqxdXRkaurM
lftnTArEOSOe2U1BZbKNQf8GXaWs9NoAYGFeM0pTkstHvpaTlTP/xNffvmKZP4fH
cZFuacrxP9AF8hANKOtByHh4a+BiQOXKvGUbA/bGifH6y5+ufwn38yewB5hmgTkf
CmE9JMCZ2lMKgRpHfZE/fz1UkkzXrDUTj9n77QN5oAt1LqwUyLxYbxSghUm581sy
qV4/b5QkkBdVnhwkf0ZS7QsSEbU0UzdBkVSgPmVj64KSrsJNUC6cHDfUkwgx6Rds
0CdWjiVE0dGGG+BpMJFIEn6oPeRZZU/RrSubCl77le/97lWDcnKyI9CQ9dUXB8U5
QCnXnmclwcTRG0loJI0CuIr+J+aVnUVrT2Zb3/Hk/XclcXIQy49W3kB+bzuWdpTD
iT/NoKIIvQaIMVu3e7MN+fhG0T8qE/Y9qoYU62PLQLqpMnA6McJ29CO3/DohtbzF
Qi2+Ez/UaX6q3sPAHYpOC7UB6pdzpBddvNxurG2aDKLIEec25cTdwOYdGyvf1hVz
ehZ/24TSkHeNnEahvM28/kodx9r1WLpBm+VcWE9lX5g2xzNn2qa8X8pFhhq72NbU
fG3m1NAUGU9GE5G0FvEmM4zBBfDaDA0fUCZkkaxmGJL9nxyNT4UV9O9VY98KdmwC
XwlKwyqCMKDz6Ak3cYlay9IIx0ROtAlILqmyQ6INefMXHM9s2GIF6XjqL7L9E/b6
TkBjncRcqUYOrbUenVg6i87lH5e6/WBLi9Kr4AcAu7d8FJ6+d5NYFvOtATrJXlEB
2TDOwvIi7byFWztirTvLsEKk763SyKlDd8g0DFpcyeN0zfjLTdaiFJfxlodFPg7+
V14o1UxqUfaYkeJbHTSFnxMmZ33cqCmZoK1OxP7XetLGjNVyoW2N+GGLdkNbvRM4
zZVs+OIeCilZcmTDM07fpbRW+Aomso/UXw8R5mDZ9u2EMyeTciNRmXSlQxZfzD6C
k+FbG2MJxiDEDLGhQJTiAPMXbxea+kDiFWu1gCXmTGgVEVBT4dM4MQPjSo00/LDo
vRBOzGN83kRuM+C+2t05mNfAB9rQgaE3sp4Uncg6ZlZlTIsIUpWzRVmr7K1zNgfV
C62wEl58QKxwSy+okpk9r0jBgpXNy9QJAC3R5JvJw5fcn5Neg9EF9DHTVzq3wG3M
Qlf9U5IzaogSltLuiPxxngmS1Vllqg4oBemVHYdn40ZluqfonUH4G2Gagb9gU+DQ
G8kGg9khUZ40p1VyxuCX/IU/EkQxLpu4Lfm9g05bvQxPSccuddtd4wcD0f+9Q+uT
OGUVvv2XlLWN/ooeRX5FOHjeSohxDRGbfaDRUcI3Xw+5R6WMKHRiHchauuV3RW56
1dOsgYJb63e8v01r/2Mgl0k6vBD10woaKgaUqVN7p+WKNviq/WCPhVT2dslEseqk
/Bt13fOPyQvuzhdoNZpDLFhiKrf8QbZh5cHBOzPizyQPJG9QyRkdYEp1ZNG9N14/
IAdQ0UgHi9MBx/gpyN4fx/lI/m8TkhSBt6sj8M/hAAY3UZaz/3Kx+/owETIEHiUl
XHOvNFYfOaQv3kqKe0qfrH7EFjzT5HJrCRyeudF/mBeOkMCYuBH/1jKrrJmWAgdq
/17VJzU9nJPFGwZBvah2bFYqDzsw/Jk1UNcSvrCMKBKV83h3HiKc+xBuGa+EVLMU
YiK6SjOS+4rVTPUGWdoowbV3CX+138/K1a7xdPVWF8a9tOuVkp9GX+0yyAv57MIx
uXHXcK7PEKIoNhJ8ZRMhIS73KYfK5QqFSUU0FZSG7rbKVpg7UZlphEcPgzXf3XQK
ky4LPzkjXuebgRHyez6T48Y7S05uh6Jd19maJCIu7QQ4ZSsXbiE7GCeoTtwTb4On
s9YQUcDvM85dF4SbRMlTzp+NZ5rZHMhH6vSjr8b6XGmCRpRJN0yx/aN4D1nMzuZr
Ylzqlj7qPhc4Ba/akHJml2lOcm6Z1DZ8gQnsanT0k6uWvMCcA+gaRZPhSp/LRbct
eU+mS7PTsE79OoDGVr5wjE3tC1FejhyIHZ+12Ro7TjXjv9qqvj9dlojQXUrkNrz2
184IrqREBdkmhNvGv2+ShDScQQJYEgfPAnvtEtmlpu5tpM5yHxPs3F4viJgLfJwn
eYMr3PMWOwontdHl6AKkVwSkbPriktj3IWy5VW4kfOfeq8kFaeAXzXAveOygTZdi
iqcTzC8OR3T5FoyKYeBcJjTd9SXhNKdvNFQd1Ec0bKe++odKB3NSZGW/p+D5TaNG
7ORN2vax4OBDiA3ovR2oBeGJNJOL29/aYHNW7i2qY6T/IpSvRaZD4HxjRo+BlYhC
XxA3/GwT3UUXuuN1AlKRiTvLv5oIWwp/jr3fMldA5woh7W8qY7QtGLrXz94oPNGl
fDt5LqG018Y51hATh9v5J75q4hsCOCny5RISJ8yFoPb0zx+TfeazbNungRtCUXP3
3Or3bAjvQ2VXAKyfBUoUA5NKPcKuwBedZhNdJTWvktNgdAxmJEnmmnFSMvYxZKDF
tGYJsElQp8MJEWahr5J3zwfVtvWA84Yn1bauxRE6K2A18WTTOo6TUFvi3hmQuje/
fnUseyAyVyej8hq3d7m3XbExPzmS6KHSuug5OwLMD/j7/ImA2RXD37XPtv3F9uSP
ajDxmQ9pdCW2DChxOnxctlVon87ZBl2Iydw6OWXwrVTSamOkz+PntnA2DXIJ9k4H
HjNWJ+78K9te8gavlTQh8Uq6HT4bEm7pC3mYcZhs2VvpZVxTfHK2AkWuVXbzH7jl
EY9D+xx81kL2SLsR9QpRmqbjP3wWavMMWkheGm884KYFl4L6b0w17qttQLlTbcGi
6KoyW2NjKjNxzNCcVsh+sZsmGIL7RzOzqO+uCBnOHUPYGqQ8LAQQolowhtnENKLU
muUSylFILOFY2kM9Q3xt/+yO79CC930r21jafSufp6c5j2v96xRh06cREJK7zW4X
goUZ3mfGEDA0Ltd/ZPIluBSbCyYIzx/Vs9s+mrbNGBJLA8GwO4IQFrSZXzk8HyK3
UG4P/yMUpDg3iy5hUPFlR/g9of4bp9HJma2jFPYK+NbqEcrMZIAWu1giu39vh9Xx
vMqy7DVaFl4w31WbfLwRMk7k3B+y7Sgi969sO+WyZVzP4YMO/WiZoOANgL/OPpO9
3GpHF3UjXVbf3OBYHWZrMdyHmpUB2ZP3x4oEEEeFtl1eiF2MnuxRMndgI8bLymYJ
kkwptlqgJQCeHt4QVe4Qa+M1KRunecTjsJ5jMryYJC2WZW8fkJho0h0nfIzMaqp/
3lCdS5HOPQtLv7APG6ws1c81cm87DZx1dMHLp4bkHJzVqWPNwFn+PsmEOuJh22xo
OfWbbim4A6Zdsd+SwVBEehGrjNg4/wUg2cnmcdbvS6OIz7mP5dZvDCFpWI9WoWjf
J1SY1dAIXFyC/4E8jEqrIacjHfDHHnicBzWOQhLHEttRSR5XPLOS2Y6bo7Mjw4Uw
PACpbfsxkS90uejUlnT8MUtN1OktKWG11AEiUVa2HhtyIRZNiv0AZbw7NpJmf8ZU
2EKdfOqXcU6NGkxzPXV5/hcSrnuwF2n79fYvxCLz2QED44KkEtIURu+vcUoPYTzU
1bKmf8DPufps/Ftt+33yMT7TeSYCepwx9pMWO6Yy/6cA+S71pgK4eYabhIiNu1R4
7bxEXh5NPQbNrAfImRRdkb3Mz6yqlhqFK3pAIX86hNjnji+wa9MBVKIkvtweiC5R
OlPMVqNU0gTvnMZBdElkdRDeHPxUBKnLicu1G1Xoty7ZUO69AuqoxaZtu0VFALV2
SInn91sNg7jJ3Ok5AeUuIsxwqer4nCVDDcNwcmN6US3uLM9fbltzmVDOWWooph0V
jSA4JL2XvQwOuhs1vSSrlrainbsRoC/wvmalPSpwr2OxA10QcN6Vcwz9C/oH9EUN
22JqKtINyoLdnc8nvSYrc4ptpPF+8O8KnILuOZo+IdZyln3h6/D4e6g9ooCEEk+r
J7/VIYlHBS5d78Tq2tR8+kJUE0ctW/pV3mHLh2n/YvcvARfMK4KVuYXCkE87+WbX
QT+uQ1Kbo2/dexEqJ05L+oyaD4pUrybf/0B09WqZRurT2/MvZdrrWZ0ts03bl9P+
i3qP6EbbeDZFubf8x+xF5fH72yrJzqg4FkN0Ce7rB60fYp8mZh9oHLz3GDYvvvqz
BaJMxlzS2+FA3IBks6uXhwCN9hQxJJkARrXitYmtESf9mVlqrNBFszPCpWMXcqEI
aFoezulI9PcUrG+TfzQ6WcjdTvzCCxuX9nfhAh8kvyicTyrsG2h1/w+EYxw7gZpv
lz35wLgT+47fY3GR2y/Tt3UfneCiMlA7U6ORVVU6+tWp7FMCmw6kpe6nc76BTkS7
IRdXT9OQ6Seh6pP02otzhsq9mAS+aq/Brq2q8nEnQcZcQ3up6edN83/7uliP4NsS
Z7hhOPox2jo6wxgVDTXYuSj+xkXF04FjcwuHNfnbD10yFot0GUV3STn1O5grDPDh
B6Pmb+G5XSDnkXgPvHmprtG1W+6rE0i4ztI5ADkpmEX3Hzjke80ylxyLIrTc+xeX
E2aq5Iw3mhXYevskju8pY+9aBGjHsS6VquOwp2u4Ba4CZYcT2UlKRw+4Xst9QWqY
mhif8udaLcYeDjWrYY4ZMgjtmSfw8pHakVyGnPsoRifwbf83nGGLtKZW78avFJu3
/zO5Nb/LkOEsboJAD0yb2twEN5fflT0+XqhR54zNS8OS+jawww/69UUtikgnmq5R
SLoMOwkrGg+bqga0lkpxFC3HUNKZlOHT2VXpUTRZZ9Gw9ETakKYmnM3PcSmxrzH8
6elyggxY6WE955OrkaNxPzPmkQR+63wmCTSrEFxNLGkH1l20zpOwuvw39c4arZQa
ll1MVI0UO9BJs1235PE2P7ctPKmCmaEjvsim/UbgcoBAahVjOIz+sC+U6siSCxNN
KdJerzydDdNeIKtLaQ5NgtDx2GDe92zm4x2zeJigvH4sr69ILODbI02wuDUjr9pz
MElCsM8l7NloItH2Km07CmZa7aAxvD+cXa8X2UnBEMJ109Dd1/zpN9ZsLTBQCGpU
gsvP4+13qUl6lrhr6YyXEnSz696wmmyRatRz3T9RZUbKu63UEzOG3zbjddYrc9PU
eTme/6sBCqgt7ttZMO449VbP3CEb3x9EHBIaqPFAzaYkTDlR8xpzv58+LttzgvXm
+JM6dkCCZsKhtFi7FClVjM0NqXPBk5ZEtjThoAbKBrGHXroPTAVS6EXo92v4tHuF
ygE8Eflrd58qpXx+vy1LU+mBXRYk4qfSYWpuZOCaTDBMCp7VtNipDlB9QxmDPL0D
E1PIlTnLjQBbJlkLK/3nclRAFWj4xCDyLXUlLjfet3Njx2X0syRVHF5jcbMXj4lM
9rwLdERU9CptGPVx1Ex1M41Xd66lXgqD1DOHr6PXJFlrqydRewsfXnPgsOk4hqMG
1rLLuuXJlEVLEK00xoiRvH1jfeSL1lFa0T7RCH30iXrkhgthTDQRU7XkgKeY/vAU
JPJvkUV1c/BeqeAAMawTdh1blBi1r6uxZRoYVnJQEMxJQp4guYd/kEFWKJGrsH4A
5pcNumL4FCywLhHoI338GryRRY4IVoeG/pBsJjCxvh7BCkjynJ71DUDjdLMHwnIo
C5WSNO5jjKNPrm34rcEgemvjENUnaBlua00vHBK7qSjNQQELi90NYeA3ur5iwv3y
UeZ88/ovW+TU/n+rvJIDuSTCUA6v52r17IlE5kUUsDTWUPYrMoGgmTXwcRpFAqio
roGVRDuRxT+O2zPDgsti4N6moMNEJmGsZ4TNS+AEqP0il6DURwyG0An6DDlKjhAt
zgcoIP0IcppmvhnkpQR8LrKOh1MazSr1URLctFMhwx2akLQEcvs6pwQ0FWruaJo/
elf/7HdiGvOU8R69zUprLxGqtJqTWyfzYJZ0NtSggO/bw7LWWkYqce6z3vzrmkJb
PvEJt1k5DknFPxl+3Pt/NOnjDi3vj9xA/QdEi6FgSr5O8oyS+8sNIXjEHzS2ykaN
YmUDR2HYxp2Bq0eME60JuznhW9pIXZ5txvGgyhOUEo58ys9eudiEh7d232D8SViu
8ySfbbNvg+ebZzk/yD2VtSQVXUfjyCj1/2q9c2WVS8RSg3JPI10s8i4qlG5xhDPQ
m+2hQ7GgcmyZamZ8+MiNdOX3pwfmL2RWFYqCLEUEitQC3jb2KkMGMisUkNRxFFTG
vA9jzrLkuef7jet9Hyk5KWyT9AbDqhf6nW8PlPNYDzvoddeRINbAnYIKgnnDc+aV
PL5+z4jMDlJCJNPAxCflqdxpTgkgCvFH9DJAV0rJkuq1Xh2OqO0+sAGP7Le9+Qfo
G231KIXITnzRdMHs5it9L6VaibxyIs5N1SmCmcSjHxiZuByqgSmL137zbDMFnOHo
LeQzSNLnO7BYNKfapFoqPcFTu73vlxqGsKxTgf1zLs+dbWe4aFOCwXGJMnvcImEX
HAyiQN1hgJlTso3VfPKZZfov45xiTbxf+uCU62NfdNT2hrC7rhPyaGcEcDPx4pQQ
o/mzFQlsvlVkcW647E0196eIkPJSdF3WnJnfo+QRhMhReIXygr6NOD6M4JBlsyR9
Gvcwve+XmtcE4wX7xSqhI83xmetlnKg3tOe7JHyG/+ue+vkI4Tbpf5Ap6iGvJjhr
JpVqUU1t+O11G4LXTjB6xwILGF8efW/TEUd5DTtqQDIBlLxm9BMrkcakrRv3jGPq
uljBmE1VFUy1eacDlrJzBTFUNHAErDkzjdKIgZQ//RzNhThFNdyVylMvYsRaJdMz
wP3xgpdA2yrAePLJa8Qs8clcsYk41W9HcFwM039nrklQY2TprkfcPAnNrgTkG2cx
vn/XG1PaL87PQhfWX/Rd2jpIyBlj9j24BipjGtgoKDf97cp5CVKMzIs01/nxwcIT
QCKS3W7Tzc+0bSvuSv9GFUtaWVa6qY3aSv7Iq9TS1LQ/Q4qvyief+6Di4LcstUg2
7+VKOujcqYJrbMPvDKm4gl73j449nN4gtX+4dQSHSHrqIY0do0pInuYXuxxDLnFF
Axvr/AiWKlyvlI49K/33uLwlmt7aB3zjuH5vI7pIRFpJZrALUOlP21xUopMgg03u
bKlpKA0eQS/myPIH4aM6fe303tfeE2y9c+XGhcY+69Nm6MC+enevxIAHX2LVFSav
yU8fGrR1T+x3q8LzEXmgSzKOa6UDvcQ65ZnJxr1uD15QcliQibGOvPfdwTIiDbAG
bd+LlePY7IWbn+0Sm1QF6d1yWbti1j9oBDD4CNbb/TgY8Xuxp8+3ju4nf3Vfb3kD
wPskON7KwYOO9G7Q4kOknkYfYTMLrDNNUYr4pF4QpBe9qWyPF4EDOIrm/cRgIkim
f9WFDEPVEMVaaqLgnTib9PND6iGKNcJqGnZ3eZtJywLh2DHd7JMnkuZkwS677/7H
Gok8O0QwsFZUybgf2bXqL+3SdeT3KS3gu9OdD5a/OId+XItFuCWQphrM71I7biUG
7l0X1aHf/KORmEY5Cd9F2RoiTnvtflhja95NUUE5P654/HzOAydx9Ufox2PioXXm
VK+1GC7e/YaTnT6kT6+xxskJnAJYgWyEzewqf8KSvy488aPNOMS1Fnmu8AWLTsN9
o0kjMnuHl/6AJC2HuqS4i6BefAr20q5qV7xIj04Hi6AG1qPGiShGm3hU13+9kLcP
5ywQruDphHmai767Zj/7VQEvwyGLCzpgV+Zfof7Lj+4uERvR8EvzPjy25zg3ZEpk
t4o7UsZyLpJPD5hBXrioubGtE48lo4WiKRl2sxgNrRo0Lb/g+C2MM6Ot41Sta2QN
Y81QpKJJzVHf+X6Q7Lw2oMhQcUlBLQCfhGhQjBdx6k+hxwV4xCCewOv9Q6WGNG56
7c1PqOlCpvcDmEQDBN6GjmguANRzwTYZW7TnGr8QHEhVX3SQAfZN9d825SN6JFwI
sX0eFSCx46hdWaduRB6iJJ2+ZsGLi6lZeUJy//vqJ9bJDCFrEtUVRchtjo9CpMEJ
nIKdfCtWSemlNDPDu6VEKpRJOi9/EREhgP4mEWfSyM06GeTy6TM6QcDRyX4HaEtf
NiS0zw0Zzy5uK9LJNH9SeNBuiN8ZOnJyHjgNsKGiyQ8+D3Jd95Aksl3bsnTvrIgd
YXx5Cx5GTQTQv4OmxM0OO7WVUg49+/f18a1g9r3w7NDNLtucrsFrvDmXFRuwnjO0
PzER3h2+YrQ2OmQa6zPniGOGTED3j9dEnwes2GTYUEUwfuYwLzEV0J+AVabcre6v
Da2YyaKmoUVxKx2qw9G3wMiO2a8UGaSm96SmkxFA0shVITsjJME5z+33P6oodnvS
kNUqvTdrSDEU2yFJpAjxt0UWwO4soxjnUiLUofpG2PkRvKCBezj731obMomY1IqS
SKSoF+OgcKb56LCXHqeZUL1cz9ORtod2tcyxJnpEQYrXjQ75NPNjiGlD7aFspasL
3VM1cDfnfM/f/WGHaSUZjw2VqtHam4XPu42or0DhuxOBMo4zFy/eMGnbvxcgKQ2g
Qt3RHFGaA5p52NJyZtYgsy43Nzr7DmN7d+MXXzbk8umTsp7n9tEKNu/cEMsjVbt0
ojZzms3RfpaaQ8ucTARtq416N8mGBvb6z1p/egPvJvHCzOXwZBqXXTt6XI/LBaiG
96JXqbUXLwASadn2fNgv17ukzceL5KWVu0/CW8vmAXMGeTlLbK2BC1VdeUnH0ze5
0Ab1qwUdl1mignYWE8y/s5Sxe3A3f8rxyJOJbyw4SaTUhwUoy2d0Zu4++kas74c8
M/5z3tMwklwoI4Ir+lIT6Euww+hEngOUo8TXzGIfQJxQ7GXCHOYTvC/sltqaBCwf
56fKFDpuqtMpW+yQBB8+q0icl4WPp4vu922WmRcWqneohfaBFFDBqyOXzIypExJ0
nDmLoa/OLiJJ+1MTt/33CsRPRNHxAwGpI6wo5zkFoyMBhBb6iDrH33sqr1Nmtlin
KWAXNskJfa9EejV9g62O9QlMKh5XVLo4oYvfI+hvOCR/gTbxjCl8rb2rC7CXwgJY
pc/60G402AzfhpS1R7rjH9HXC+9YqDUzC0Gy0trDP8dkr53H2lYy5Ig0RmxByu2w
O7vX0u/awnR5+9XNq3b3yNiq95m8uAvWHf5OKXwfyr3PTIP0n/sNlncMMpkU1Deb
JW+vN6VL/zUJtW6sZ4scnKOjRyObzp2Jz5Xf79sx7ZSSL47wJuKmSX+sjFDYBwR9
EnFp9zAJr0mmFMMkvQuge8MGsM9qg5T4piaRiX8RvarNJrIfKJbqQsjoLKlrMg1y
tml5VYI79EXAMi91WAWxfjtq5iJzyAX+X2P9394d+NjbEn1CnT/quXexdVHbo+uM
7uSt2nRs9rs6RGKNVS+KNCZz7S0O/Mk3DBebJ7N/6U5/YtkB4vpU90I6VlwdOrPL
4YVTQYmhYmTfyyZEeTA9XHL/Ce5eDkbO9gzjizX894Ss8QaCK33ZlSyB2x8AuTQB
aKjLCmQlcXlxD93EXewO7YqQOpG+JxZk/4TOo5loJpLriy69Ka+Wj6mUh6LKWav5
Mn8WBM/rT6618RNA4uDSYL4LhrdRLMyjtIqelEzG1v6l/iRoV06+q7Vb13zCXkTn
Zz0igXRhO4fvaiIVf0iHxBuocK8pZCMIUqgEbjpaXGnZxB/C0VZoGaEgnJspVb82
t34rNeUvAhSEdl+TZdl7HdEOxE48B/iZuOjBU0kkp77NDa2wKR7tp9G1aWMSf0Cr
QYYS4BPmJj3AT5y2YJosBcUvRNcHo8Zj9ZWxYyfKp6L/KdVizOzrSM1w/Oe60tdm
OrPq5zhZUdfifottXLa1G7LQg1NGfWpBXL9XZnPP85pagR8tdili1dXZ9HBoFoVW
52PPOt/237d31HtC4u4+ecu0ejy38J5x8xO9xV1/xeDh1lTvjUBo4eEwLEYsHgz3
qchM1Qh2IflTfHEsdRXrBNSIWh+xJfbxycYJ3/zLCDjE5y6RU3f8xxpbA31MZ+P1
IGGi3QDkkVYAQu/expr8aneVMLHVulboEmEbuVP556u2pAqkpOyUhbLNv6KfV0+r
gycA9heBFoIGKtamv8mgyIxGUpWF7fPvtf+JoRlG54kDBW49rti0Fv5viU+Mr7C+
EMF5iaE6JUxJ8uyfBGHRu51RKk/BPq/B4BoIqtsw+XtYdlSeI7CzPDxyy1t3Mg7V
teIi/nRegjfLb0d2oxQuanxJRBmHecg58XzQN+c1c3a5WKSIECTfDZ6/A3naEA36
EZXaHxy7ja3fPI8t0nKFwMsBodkfnJz3PXsfCjPTuURjBWhnDUJfr5lmjt16+j0U
xrxLfYaoEZ3eKfNhkKSafLAYpZl2hVSex2LTBFKh69XFDJwHMhq2JGFG6disSaNG
35oXf8EnG7z2jJBKkD9QYs9nn4aq0813WClrTS7ApPKCxpK1UyzfSAY3uECQMVSj
rcnuJiA6kx7j56QEwJ77dmuDFLS2ylPTS5OOgMAPHovxr12eG+O4Mn+Yq01ni3iV
jQnhzqtp2DLi8yxI6/+a0TDtyuDBs71s2+aQo2QPUwFVseRZmIOTD+Od+8X1EUaJ
SA2No5LbZ1KyBqtF8wqL8/6shOpg0T5sMyR/ZibSKv84hjQ3eZCSm6l/g6UOL+7N
Z3ZJjrrPxxppaeWCzD+pfKOySLGoDPI3iYT1+Aalj1z5FMbpBiLRrTmXMhFlnT+S
1HGdegfRe2vOf/ModCPeb2ZwgH77paKB0FbebgtnmmMkABodmxVHOmyDyX6CqZlW
qyMBczlS89rBB/qI+PgwBcLGQPl5EuIfddj5qUxraBlUCB2z0VqvLp3KuCOoK2du
84XxtbHE511IXlFickHkFGOe7YKvopHIG67hMLLItQNiFGc+PBHG7f0GWAa5tNEv
bHFeDDBZE8cCavQAWa8aB/cZWuqDh82k3LGIQPIOFrk68w79P5/lOJW9dbSaHjDU
Kl/I5Ur/scEqniXem6XorVCweMmXZvDw2pxRjSWVPKIj1BH6Ny3a+SMoxI8SUrG7
t8xv6X2XaJwMMD1DjYNUw/t+2BPN5gIDA3Vqaho02//lZDieILLe3CjkEJK141t1
ls1g1RGnoMrF7HkEJj+LaOtHh5DVf+dFJC44/NWi3rxVUt2jP63hwcDykVVzrFjK
RlBbNFlPRJKeJsYFxDHeeV8QR3N/LoMPbzp5M70KVMG2RCmN03SusBFs+1BExrrO
0u3urvGW2OPnuOrBfHa537xS30DpQ/TRz5MxLTCWN6F8cV9ImTmevf063G+ao5LP
/TaO59fRucOIol458W85IsFLeHxeB6xCeH43xApCCriCuJoX83Gx9OjmniQ9xTqN
MZOqHAln99iWCG0jyXXwn1wyGMGTC8V8sSX/9Vj7mZ49wAI/TYCUEzZC52EM1z/U
DGXC51IfCwHmx4eEKZs0euN6dZ/3z+ZONTLwk3uyzf7yhzE+ULIOq+uWRjt1WI8O
234sisbFW4RDldbjoeNzkcnx95NKdb57OWGVm0fxbMNl2lUPq+yGgoS4cLf+/hxx
UMr+NtPAl1oc1/+Z87D91FoSpVDKEK2FZvbWCjeh5waQFr3gsDgeKA9lqYs/Y0eL
VkLiFIqLs9WWRIB3l+6XNQS+wPH1vVniOvly8OXSJPbxX1dvdVNXx1KV1M83VPaM
N00P8J+f1JiSBlWk89eMQRhH9BqAfdUIjirpVgsLye2N0zPrg8irgcgTVz/kGBso
HWHvPYlFun8Ag1MMqe6jaZWqb7ZemyqfbP8Z9R+sBGZAuBrq6JaxRovdAXsLrN89
Bm2Q+RL3e1v4kg8LMHS/Sq0tdBM8LhEArMvcvBD57hDDXazDJJpw1WKy8bvC/hXV
ucks6Vcv9cAJqNeiGnQu/qk8sVyhHCh/lNuJ2GFeW8yWt227LbawknpG1zV4p0Z0
aD5VJJ1T3zqs+f1on6ISUnyndXZNtd2u2eIOARL2cAf5pQoFpksDfHRxEHapHM2v
VilBU7ZuLVRGVFVU4rXnjVa3Z/1fcaINNnEUfn+PfZDIhB6VO8fz03mVri7Isq/7
fd7UImILKOdiQTek6Jnck62+ioqbo0a/t7nWg/WE14YNRRfG8/Ihzeh4xbQQrOhH
zOlp2Wz1QIsqTn4wm+88Pf4URtFbBMukZO7+hS11x+9plXv779IdoC9DZUpwXpQx
x6Lgjsw1ZM1RUa4VdACwWU/kMKn3PY1bGIHIiHOGD8aozTUBKuvuFF7//xWjNZ+H
eqrrdItyvORdG4h3hcU267T27Vfu2XOMU9d2NvXXypk1euK1sBOVBqeMGyOmpKVM
Lk5W8wqRkgnkNAjlcOo5kpGMM8+2rOT21kLnYY/JRp4GG84vDHgJqVPFtWiCFip5
xYLphP7imlTaewV9xrhGZ6n1Mh7Jq7RCYXOoW2K5p83TzgsqMN/Wf26n437zYu7g
cb/Vue/8fqEyuj38+MnCyhn6BmdVB0Yh7HkPRNPTgLdXQ/tcrOaulHp//uDP+vnV
gA8bLdxGvrQcj5PIctEE97/P+KkoTLiDMfKawM666xl0R43+RsbzwetZn597B88V
U4mtaIVB7vZQIg9g1y7jgZaRLeB8HBBgdfPhVRDWO6SNbdhtsVf4bg+IUXsLQlsc
hHkMUPHHp/QzLLCW7/4JJf8RAi38ub0TtZ+ci3WHhFRRDABbeG7rbMOI/ZYOk72p
YKm0a7AVRtIYehuCGlmfNzwSh3+3qu0ueQeFRi00eL0RT5R0J7j1WBUgiXmbfV5L
h20BVJjwk3YDCJqFTlF6yk/QLawCejgY2Bzbc82x+YTijScYoNAW3Fwp3ZyKxk7l
O2AcAp0GunWNddFcKrb+YSpzWAvPFAqugqvtxq82/byUKuiYSTUDKppw2ngQYM6g
VzS5UmT77VNEatoHuXMj2QCiPlicNQk6D1N9q3KTDfNCV1WjI0OY5k6K/2dkryqO
BlEZQ3z9PiOIZmsL0I5cVzKUFU4G3IVhHVMzTdhox7RHU0OR7xeUhbdChsJbNMvy
R6USGfhOOLCspX5N5LhYEjYbT9VLxcy7C1Ovrt9Jbxr6GIkwgeJbs2cAFlBqskMP
8HZZa4t0AkmcjY8Zge7CKphgfEwUJytQk+PsVAwZ1l2qEnRpsdE6ucLnwdf4YzCb
7RMSYXecDjGEmc0MVtyl4H2GRdDT6eQ+nhrIx5YS6rNGz5RZnaA6+mopCLY/Sy3E
aWYGe6DwvHFyEU7XwGKrR3/vL32S1pJGYp+IrFmqmXD4c368whphMQc9Hv7hqWL+
OrxSMlUi7kZ8QRkEnG6VsVJxD1EBXkU7eNKemw8hae13ODEzVtZd6JI4AOknSzaX
eVEq7jmvHqfXwLISc7moSKcINiqqa+wwYRPrzuI+xMIEZdyV3syHoTKEk+lZgMfB
MK1hI2+wDhy7iJ1IGuQe3gU+HAiKETB5FIbhE/6qKqyTrpSru6P7lZm2bRgmPdkf
4w/jLXUhfvinsnnVj2XnOzyDJVw8J7V1Wi9N6AnW4NslqSjfKkhlsF2q6W8JNQ9P
NKMm9PPdPPJZnDbDpnzFxnuHOIDDJL33NP5ZdMDCsI8idtvWi31Qs7LH3Pi1GCB8
ocWp/rTDfg5isq5vh6An3ERq/o1bbtPlVoNwkX/hTq5h+gWQv+X2UPkwilMYkcqS
gRJOe0sKX1Gtxh3F3It7Wvj9clbMrnIL+Ioqu6BGRsp31FAiTd3iNz8LwT8twMAJ
MyOjHzWbU43A9W4ddspRXUdqQBF5nnTlQ4+fl6GfOb1K1YfDZMf26jAmLq7ThIzY
n0YxqS9IbIXRCXjTAeevst6eaiU/6nxTK5fNu4OWf7i5OUJPNge+RlGEy4z2iAEZ
sI1vc2S8//K9EL4/qUjq9m58G+B5p5XO1HKX8K8iilNRMoSOwEKgHdrEWZujBoUM
zT2AKVrE/Bzr9Cg9K5+A7poSn/UCdu1/d93kmzTfw+nFmd229welnuwdG8HbgjFz
tqdPcfNvxakgGIuHtLa2elYe81lLZz3zDHGjYCQ1+N5zt3Nq7yNQGKO9kQX2Kgqo
AMhJA4tfZcy+CiCvW/Ey3urEi+CXHQYpZwXNlevyHTayi8Nu8UGavF5CUKffRpqv
aHjFc2ukVQ89iBulS3Aa/LCE0HNN0n3HucncYq0tQ8dm3FIEiNKLkT6Mxy4S/sRe
j7Yvk4DpafLnlag4PGhiaxe746pgo2S9oB87TqLR9A0X3nLAhZxCv1ZvR6/bAPl8
zJhljbzkdmTvxjTCMiS68DtbiX4/3ubfZrAHLk9qI04cdXOcalpCRp45ug78ceQ0
+lk1Q39FJaltKw8LBroS2/Q5Lf6nqUpv8cLe2HjNo3oKbgDbGZ1mQDr61vI17+yF
M0rBDJ9D54L2slIn6I53BS66MV2BS6pN5rn2ZFnXMi4FRS4QFTtezjcKMggkgFfS
YLCwd4Ni/7mtPb8dOvilBGdWCsqI3hnuKeHq2AOwLwlvlbG/UD3jIoDr0qsHbmmx
ByF720zgcYsbf632D8wV8ZDH3OPmdrUhcpm3SllbXmIQsxUORtLHIGDXZlmNTpgG
A2eLWZskSJhqJTJPMIyJTygrgSKUpp1BD/I1caQlFh0zNZ3CRBJRhzIsmfa/4t09
RfLa6u6Nvx9OPfECQSS8+c0lHyxAmAnV7tBfJt8IlNQGw5nUt0/zjIjWBA61aWuj
Mpi5fFq3U42zmKVH051vEX6SZ4l7VidNuX7JRfm3l5WWyDbZQNEnQeYFsmoPUtFz
/viR5l0A6ul+QvZaGc7xmW8vyWJOhpT/4MkM/EAIak5doG66hEnb9Q67K9MjoOkB
0Y8UdRitw1zdVsbtKk220UsVN6r5b8rcOMSPMgC4DARHw/aXYYP04c0fIppnr9xn
2fa6uS/SWhdMn2sQJz88CxNigmLEYEvCqfIpaAjqKv/dItfqsNVb3d97wfb0+Q73
icGMZI0PawTNiStckD3VhiMKsGqMSl8rUpq5cMORDwbA5YTTOJ3JeorYWs/W9vhx
WYmeny77O+Czja7+6mh0GGnF/w16+4sB76k6LoZrC3RpJetsZO81dlnsCoR4HXdf
pskhiLbhjKBafTbxZ9O3OWGNKvNBAwV8W4f6Wxq82HLLdULfbTQlMap+xXqAelrE
hLYy1nxFTz/bX1tQC0PMfiFgh5lUJeKK9SyBaxvPpz9wOg7t372KyMAOdVEwGqxf
rLyCqkbZa8glcTZ3rV/s+O0jVJorPET7Pg4/mKDdkeWcemaYtGAYDvpZ+mM+aOxO
4zIPOAJ7qL9sG/m7LhrCY4dKk2oaE0JVTvneEEgNNLWcip1OQJOo9SkZO4PLweFx
hg7GdCsd9RP0TB5cIXMcYmuGG62C4aZfyqIQYApze7oGd7+aEA1WymY04yX2yd3Y
qcQiHpmv1dZeu3IovbNO0aEHmDgwI4D0Yd2/FF0mXMWd3ms9gWaEe/UOo0hjILuY
874sPbvCC3hw6ONkghieykc815yfcHHWEz+D3bplhVpxin/rHNU8ZjqmOFDnYttt
Z/w2iu3QXvjrlp+W09WVkHhXMD9jrh26UwkBVQ74+OSz36cas0yewv/r8shDM4Kw
mmZq3TEWl8VzTIs5+r6/8bofUBnH6nUUu2p1UYURVRewgbvjtp4bngfEWIdMs8wy
amObCmLbOwzedoSUGKTGl5vTocZUoWUgpBz3Bz+KFF4X3h03UoYF1oESjODAE1kD
O0QMatI220eWCCKzLeArrAoUOkVfsSi9XkcGkPwccTRHqKdvJksfN1dEx4Hv+7CF
ax+b5kv4cvIDeNRpLkd6V3hlB9JoOHihXVtPxJOCaX8+7iVfxlkFtKDS1gzCCLX1
h/Iuv6Bu0uhwZ5fIt4oZGBGrvSlRDBDTHumjXdU4opHn+Yx7dawzGV0Xgk+S5PoE
/PEq+/crSvvLgx7NOdLfPZkI+p5nac7hWfwv4m/zRILrt1amvRKxF//Nw/iw1MpN
U0wypYwm9JQaTvNwJhOiIE8uYEfLbtrlGxO9QoSUnGigWQQmCKHxkwu9JuFbQ8sJ
suy6VmRYxz3lRguHe6BCGb8wDCiGBtgw+v8P5haqM38xCawwzl3DI+u/402NrDXE
uhOWLuG7wXA2OV8db4sP0Aj7BQbp3II+xef0FnFoKfb/tazWYQ56p9qcCdQ4DvHX
H8nm+HQWTYdEE4x7qVPsgHtbsKeBlt3jlhAoV/Y00xwqBu0/ZdtmvKQKDqna4kFI
wCc8+etporFzs8aWZZgzCCBGFzlpU49JpUDB/CurASf+tdwiTUtRsM98Tg/93XZv
DprmgdsUdvllocQ92qjumUU/gHggh+rvnuf4GerInKNWPbqxFh3B/xAwzRpCnZrP
1WXjBi7UkTY3uv1AEjCkNTqlk8w0f0qMV99VttTmylr27T3c0iv8NIsLLfBGL+rv
1OUUNHTDah94LYEkFYrhU6eNLX1rW5PnEwh//5U6pwfo00pOnVVMDP2FCsNxMgYg
i9EdX/X+rSi++UPYRx69kQHM4gPpvTMOqznrf2rRUwU7xe4IIZ9t3MnznqtdqWo6
dZuE3CNeaeOt3wi3zWi+1ilsUTrqd1vxMvGmLfyKw465g4cNxMPmvfG2dmo/BZJ+
ZIFNZ5gJxH5mlI9LFhCv50W1NE0F5PQi88V77ILxTzaUoVE0U065zlR9vCVtXQBy
/X+G+AM78i07qBBcUDgZR2rP0FPlHOKwaIZcq9uD5ZGGSySL6HG5phNFEnEontBf
BEsxm0EU1NZrzT9S4iGBoqrghE+DDEIlrLMk3sKUaEkqytrJrnZx7uB/TDFS8heh
cYo58n4Z8K0B87mBQX+eBLzTn29L+pOq9Qp+1QFIkXHXRumarfw2JIoDzPzkJSjd
8esIX5kFNJD4XmIngsLBbvA59D/J2ND6yU/3i1fCOeX20uxB6FpNnHTZW7yAuUw0
Nu+ZLcbHPXROaOziVWeWBUvLkbuaJf4a6S/liX1B1mNZidXHddtxW0NA3Vvh3k6t
ynBKytqSXPkxgJb+kfSBZJdGPKTNDvqba/cYaIJRnWlD5bIC6ujgE9j9YfDwlbik
/V65lhcIhM/ZpsmM7B9+6dk6lqzAAKzdV8jdg+5IVRqB+X6hOiOYlsr1hLG4i9rp
D4N6HLo+CB/yPjrx/dg3nEEHCIkS+cx6rOUH5th9kn1HFAiqaN8+mTFN6PPgDE0m
HI+oVjqp7GpZsHh5FvoLcCxAQWM4vyrAzOmx9PVunbVqTEKeaP/Ng4uvc30piqbs
ZU4QQQZvuvbFiLixqSD5ax1Xa4RKyQWFi2V/UJEKiaENfDGUtsBM9A1xierGtdDx
64TFyUXnSe2mxNpCG7fx05vLZbEUuQiO2EE3V0jcrbkDe9GNO2ulugfYWE8cn8Jl
tmCEAV702h3fGZvaBn7azi45VLMf8IKeZgr1XuZXSQwPZUn7RkTUlS9rdo5MPrzn
/ypQu9es4T30fGEaiiURSqn/GDMp+w3zSruSuwPqwyx5NqBT5VEyAwdwu2Eygd5A
RJU0PiBFv6WVrnnV/Q94xpSN4/aOWkYFxRMYM50kqcMXTfsK5de8PKxNm9OYsedh
9uqjig50q4OiFwoBlMpFe6hPxEbVa/uvrYWrksDLpfZkePC7H71A9W4Op0xhLaZR
OBZE9TypebSiUgQtedsBXKqdd8de38xEclCABjec+5nkIbc9GumswKfPq5jVAXBg
1tX8IINIagiTHqZLkwWDJkm5AFARWoW7Oax1vuhgoVQjglJyTLjIxRY1pQwAOT9G
EOnmxQ8eTTo/0lWP2a2iF+I5owj1e94C9rybHKisLnjnUQNgap49m6FG26H8SUmf
pHRbGQuOYgYlLq2u1PNWvgVrQQ67CQVJfhcqoY4Lz0eZ4t/DjVecGfY8/Sepe45v
nAebQkYAfCx7tFXzNWQyGvq2JuyV1hx8RzJjTmzSV8wtZ8gPeZGigmca7sZhLWgz
tsEybjHQFZmeM3fOKpEiOEGLdClz8V1VDT2tcymXJ9mWqVHKGWk8CX2WpWWWlT5c
zKmUFHOz3AVTdYExhGO30JAPEUzbFWdJ6HmOrxSdoPG/ks9OQaAfpaBi2UZs24Id
3SAS/wYSyy7ySxj55Ak0UTx29rxAMwKcVOtFAQ7Vc2jiWh+MMBtYe+EFp8MK8Wzp
RNMMjQkjELCN6tn6c1KwK9L03Pt5iX3CO5mefx7BlZ7heS0oRtX6rj0CNUeJiBiH
+M8HX7g35+hygISp416alx2oYhqdFPkw5Rd589BU97lMZILxmhIZNLn+5uvhgTJh
Cl3FImeCqy39b7joM8jNH96wGpBh7Y7QxElNRPvq2gdfMannHaY/0TJJL2Ma4B6n
M3+Ot8TXqOurjXP8QscRJWuauVshH8YQ7t7xuMcpZZHo8dPmn3jUTL1VCn5iTMYB
W+CxScV7ahT70n2QIcjnWw7ng537S0l9ZgiM2+u3oUd9w9EKxr0UpdKIm3d1ccBu
Z8mwW28MjK9roGDMH2vXFGMu7QFye8yTaor7b6/44mnKWdGI5O1PhEXqg8y3vdOp
W9X60ANixopxaqPdGEPfkINmmAkTTSojWgsJEme9Uo7Ox0YFc9PidksP5V1SJ3WQ
0VGrH68PZMieLmk/6ZXPKjEQ3S/IMD1F+KSVUjcJkHJZjJb/ZoaaCo3rSScfMwQD
A2lR8AmLhuloCVtBPVyimOzwZqOSSslGdlije70W5jeOREk9IGhQQrvnG6egKQuq
SxBlSE/zXDTIaS9YUMpAOv4y943hkKlzLR1V9goqppBCNoBxrdyay8xLv8qUP4dc
RypJvcXoNMSrXVwG1X5LrgcXzbONFgwz2Olo6OJHdiWDHT/lfG2gxiO66kc/Zqyn
4jDaRCHRCDbhINoeuYjDIXYJ5TdoAy5VHL5DS5xwSxUY6ViYer93JBOBc9nL5J7C
Yt4ftv3PUU0JkE9tWO1Z2o+Fezoa99JgnFkphSY4DiB9xWp5/CLBGumHA2PpnglE
7vlNe+I/DwebtmyJWbebrZBrmEHpawfKjaaG7luMFpsgTBodzV9RxdWGINhoXr26
e1AWQNF3+ORUh0mtDEzCXWEoNs7imKpTAEsoeQfsOZDZcrCnLzIq7cQxf4hSjhl7
mQ4FQZym+6gcUzMvC95pj99sw+zyNQ1rwO6a3XhCic2OjPAStzYA1t6fhDeyynAU
+lk9EaOHvjngLOTFfb0kJW+MnwyFy4I4KPCGzcOG9hfxDD1r994jLOfcrMQnYkAy
l1jfJGYfUpYgiTilNzIPZiJARGS41HqPnYTyWg98dm8KlEfaBVhzbgAaUgksiz0o
wKhaliuZoqUZpkwwZTJATrMkOFTDX4rVXy9KkXUq8II1u/uurpahreBhZkAPDPAy
BZ1z0RfqSuXUPXCL54TqtMGcXjtzO/C5nzEFwcYPBDQ5AdVsDGA8iO1Cab6uqip1
VduBNT6j5aBVjxErAPY6L+vxEVWB4uMNrB2Py0kv0DCMPOxxcQHb+bTYskDa8t1a
Hmqzh77IQa0xXH6yTn809KjaDmUu2TgUPhFDvRXUDtNox2Lnw0FRFPuwDfKKj0JE
D1W4ONyqD4nclOb2rtAYrCQ2OMfij/31HB0jYmdiIDxuXFynStAQwiwKFQq5FaLF
GOo3HLJnLqR0A8XiIx2Y7vnhUCbKAMuPQT3IS9QycRqmCJg1VQFiiP5cGGTzeNcM
29OBlCwVwtHcWsdJFoI0nhV8j1CtwzkcZMeYMlIril13lDfZXsMqRSOS4qL+Rqsz
JY4k/+m0Vm2F2X+cBSEYEnTLo9jcd+Rs8CLhBHR4tcsqIGQBJyV5+Hu2F1f0waba
IWuoeR2gVzCFJhquGV2DAKrcmzBcFYzUJPeo/xLTJkv36fYmuEbSdF0swHbbm8JD
3fhL7vZNwq3a6MeYaoclyp8QMh47HT8Uys1tN7/sSZBv2q349Gi81y0wBQIiupEZ
IQnBXppnhR+xEZewco1reE8pI8If4tfQ9ZmJk/GBr5sNqVE/C2yx1P+t9ia9hYZh
GLtq4cGQ5I7FTEI/+NKSFSFE4EijidMPvvB+1r13OISU7+IA/51wvTqMd8zxkTdc
VCzOm0otzOcPXafH4EYoF7nsjUl6v9qJjR2vyQTmJLLMn2ES0COE651/zh1TIUoY
Qg0i4WicE+EUtmeEmwKqsNxJyJgNEjPR2aYKBxStYjBW7jwvNAqbjjVItVslD8ZS
ePKmVDNxUPU67f3KAPLrQOHh19P3cFaZkos/NqThTZp4CIPT9wDdAa/aI2hI6FuL
zrtPfzq3jnGUu/Ixzjfzx2w9HjzsnqFRHk/JYm2Z46I3TFizeP1o6ydmjefucGDl
bLz0jzMXLfrEBEhvm9qVl7S53fyKe4yzXV40IMPCSgml9qIvpu0LAjBHj1Xo+Pvg
rPinjSwPlmLP2Vc1jFi6ce/THyAz2W4hQ3Ef3/vdaqEfa4yJYx/9qPNydwVJKRv+
qdpdMajQDYnMmAvnV/DXapsaMNme0b2wn3dD2uqmOmBP3NMfcLyJY1YY98Z6zzGZ
0PWtsd0Gu+3ykVCBZyZdR+OR4Ss31+USooSwShBX9X10VxB504kF99zzHEhTdJk1
dJoSdW3yFt4S5uZOvDZRF4w6OeyVYISEnDvGg3kQHe7fqPn2skpfhYxohVPFz+Yd
H8MRmnhMr0dBMuUG54fgGdOgrBltfy07JAD7v+G74wNEojo9q3c4b3cMerY9yJWK
Ku2ZgrcBTMgjCfmPrzdxuW+DyqoxY9vTPccsrnGD2NClfa3RFmNhL3C869hdJSAn
JPB1hYY59IIwxTtDy9dsl7Ob1jC4AeN7+5FC9W/cxX+Cwrmk5Z/ci1EAJ3SIB7T7
9GhNdY7XFqwq3WO1rmulk78apWpm8UkibugvRU3DZ9F1/cQbwF2hbLsy4GmZ7fIz
Uk1pxqG2u6/i8aLJJCWgg4yWUG/ZPHgq9Dynakkros35vWI1gY5eLCc7K+2z81yP
YO1T0BANCLKRz00Ham5XK0cWj+4cdq6RQnhXaweGvOQTz4xPqfWvQ4NZY5nYhf+x
ToMa1GYRASxni9kf+SJFO+lxL9id4rGFtUuKNtZEfVQt1S9U8Dq1pVYeYEn81Nxc
GmXGhYCaD7Cq9WpZJmqJgEqfKD6DvLKHBifVpLSKVDWOUzW3cnPAkgmnZEss6k3z
b0vi+GDpeoRbGCILmPFifRjGNsRTXDQFNSc/JE+/T45VyYbKksiR67z7Q2AgN+AS
Ea+UL6/N4UDIVucXTEpUpQsVX49WjEheDV/cq7EgfIVCz54Ui8cuHoQzQSMfNuC6
QjYcNxMFsyTUlo6Q0da9AU52TRtmo/KrjroYcU8dbt/i8F7mh2PWiakd7RwBIB9l
v0lGIxChtEGL9AVfl8HULavVFm0v0XlB2F78sr02JOYddeiv+QNnLKZsTkWOvecV
61JFQuRW8l/3huMUhIeFiZ8n0hp6Yfbs72qOoGfYBvMlMr/3mYyFEXxwXJB85HaW
59rh6eUKpz/YaRbjD0DZeQRO/EofybWmEY+RuYKCHhjfSNmnZtjwGQ9wW29KM2ZW
5MZu+jsfqPXIoFGDToNJccBIYSPf0kr63L9/TG23y6n3ytTvNzLQVr20F/KNsIq2
3Z8NC+gQboGVlDG7Rt5Xep64dXQBsUuIHGL/DXi2EEF2Q7zg/Wnn1DDOHzKNUh8T
KbvhEtr2dGxkfuOsmS3WJfVDW5KIvrbPgwjJ7Cv1xAJI2ZRci9rOFbDK3KA90xQQ
vnnHsPkk04x1bXBSN6SU2fiRF26LyparNR6B7JaH5fV2vb/9zX8CWc7mPRo+FMjb
JhmyBvClD7BBOYTZ+wWx53adQoZpy/5ZiqOWXqpUrH8reuUDCUXRIJVx4ToYLBEO
0HFmEZH8zvLP6JFr9ZhzF9LewUtoYh2mrgRuxTXPZg5PnQk237VWOYSFImXWsK9g
iv+gvTytxwY/HGXrsc6je7i8yPH5gd2VFDvxPam+mj1aSG/3p6tR0qBppk7dqyMo
K6kSMQlTSPzkHZ0cSzOJkRobNOxgwebLocYTW9KeVe44s7/bnkDbsOOndLofOsHT
bXBsvfktcJHxpSt8lO4TAsoNkiSHi1x/M3DaeIINT7/CmqSks6YOAXTN447HNEen
QgfVswCrqn+VuE/Qn4RPby2Z6cfghSTlm2bdM3hV2/d9gbvC3tZRblq+J7L6z6/A
kbqCqGh8lBNUCbtHeXKveOZXYkPNGuotOcuCftOPrcSC85ajUejsZkH3sNevXOBS
sCcuBlVl5RfMTkJthcqSNnnBfSucRHKR7SakMLaOwSXSoReazqnFTYxpGgyTcQcn
3cXzEerNvlHdfOoBqdtZvp8EAhabGxu9KOB0q/iq//2hsdHMrwBrAnteSFFaGAST
RT+rroUFBATnHCCVtwM9PETJfkZPvVdMmoXn1V6Qf4mJS+uAgO2AyeMIxH9dDYVw
sWim0gpQf+PHVwvDqLmPDn6w26nKzhBNi2Q0wD4OoZXvsZcPec7mYHeSbMNqnRet
IUb+eI0Fy9CTgAZsM7V66GbhvKFNFQBHieumdq4vUHFnA0z+u+0z8isNmSZL8pSv
sHXItbVIODs9pKMbiziqiDKQcBnzgTfxKH5VdWCGVdofMaIFNECagKQfxfYoOUJ8
qAU+BjnBWp7IEO606RlmNbguhgXw1vSDXJT/mYr/pJCwCxNYx9RkCEOosdIyw7zU
b15Le+Wsy8VAXQDgMAcuFruCuOnlrdnsyWnQVNctwdBH39s4ZTeJm+O03t5eTr1L
HgEELA+DxelUFqivB1AidEvdYKwTAQqJA8ViCApgCZulKnwNZ3CiuN4DFtwqxHxf
/XjEWro1aLGk5D9QXd97uSFdPXmRhk6mOBzlVq95HRMeBo3nMcla0AazlprzmFCd
AaXLoYjhaHAY58lJDYW7cyCh4ZWot9X5b3ne/s2DKl2tfitWra4xNsmlpCm9Wwkv
CPXcmNSmmeVhZDnnRKSf/FZGHa18wgwLpI9UE0iKKgOn4vFM1sJ19tQ22BzYsxY6
s+bWm3b58JpBJlFXVKDKaxjbJI2YpfE7QcX6ertfM00e1KAM17CWoTAMH+p+HLDF
G11OnMwzqS9zonTuU1D+3Tl/oOZ2fnyqQIOE9Hazaiiy2bqrsgbRVB15ei9ZDx9A
EbqS0PW8wwRZlN1X+8rhtqI76bJlWjTphQLcB2N+IwLxncFE1dr4bHFFvjnvwJYS
NhQ6hZAsM8U7GRDsqjinMSMkC6x5Prx0sVO9E28xEpvjPPc6D3pPaufDlYbMTzGD
svy6Fm/EmyrgzqQsimWX4edJ5aXst+u/MHpGrm7KUrqtQJ/M94TtaYwFyaHNTEst
YOGSuVPTF8R+BMLwsr2O8nNi0+yw6+AST+VSewJSDWaaB2WfmLkgFH45dAo4Q3jd
26/GYMDmr8OoSFOAJSg54RsHJx9lCtZUynU9f8xqWay+g/CnonkOLCJ1PgreXTP5
bF95QbPL+btp8Lud0Gqa/5Tb5nTCrs1MYPq6T9Yr5V2in8dySGG6Mq+3N59fKtce
anMLM0lPQBG3elSFd61dZylK+H3Q/ux13PHQ1Liz7+OgZDkQ9mTBc8KudAKm/yuK
K+arwUsFFXyt/BOWDdDelOv7OLbhl/BncuRmBUii0ktOQmCAsdtWSyuGoj+CFiw6
H8VEImxV8CNQuzlbSuZXUlHxebxkvedKtV3ASwg9MeiHRXujR6Z7gepUAi8/e3iy
91vKKU71T7hmcG/3WePRN7STB7L8kgFXn+KLv7yqzK5kn645Nl18Lsr/pykCUVQz
rWAwjdChTd2hwcnzgQ9ioRbWkd+0dMm1OfUMLE/e94vdTQRF+0YVq7oRpCBA9Lve
Be8tnKHGGpUqDPNOqG/A/70xUslU/gf6zh5PF/Tq3e5nATpF+eNzOAdCWuPINjvc
kD9pUX42Hpr/08qokKvmEqS5qLTOciwKgoRgtsyjb2Tsm1edcaGZaGHAw/hE0t7R
OI0thAwdPAZKt0M7C9DBUfk2bJL1nNzfWKKnbFOqr1AJMLykybXYhauo7oVCzFLK
22Tj9v5V5seqIe2nt9Jlge9IyLE90v0xrhf38BQq6hDCMYZDEOG5nCSqTDb1aYsF
0VjUIgHuHEgXUMj4SjkzqxFbRyMnIXhAbrDWsRsBPLFZI6nwlYfplCbhTP5YeDvM
72AqU4tyuJXy22Yg4onHH9Wjd79hyCGnWqyAAKargJ7+958cXYzDeoFlVu1or+9n
IZIhJM+xxya7mYTD1VjDS5EPPYBoX9GIwRpwzON/1pgzEmXH5JJAqpqf0xrhUqRx
Owqoo+MSiJd+KXy3aLoHemoXgQNbynFXndt7fP7dmI/t3vy1tsR6JATzc0rg22Xt
dnW1MsKkTglXLHT02D8zn9ymntBsuZrHtIb71LW2QXvvFYYFUddWoaZFtL0GSOlK
g2blj6CUiN9GnP2iy3nrRE3iZz9SU8lbZU6Q9dSi197QQAgazk5FQkuw2+93+v0U
Yy4s1UXRIlw1/qV9YzUUiX8v9OJ0a/XV+LGX1EFae60oR07Ubl5mMo9/zWNnzO25
d8lDjHlQQQPXWRckWj3+nDz13aVnVQj7V6i27ov7OmRYgwXnFMHVBZ/6gLBM/G+p
YWpxY3mn5Os/c/tzpVSVPcoUY6oFxd/vPaMqZe8rr6YLBRkAzK/qExd+G4h3mMLO
6NIfITOD4Ii2Cy5aKLHsL018TFlhM/vYBz6xHHszrHF3AUhwZ9NOAJJ3FG8ruyQi
crA8gMrXt8MrwoGoEALL4A3mRLwp+AEa77hl9iqFBQbLWgZLUU15uVQkxiip10oZ
TGAC5E0OowR9EipJbj9fgG0vBpnOchyy6JztFm2YwflA6JX+MS5yy/zboK9ZKBHR
VP1nQkgVgP9c4a/Q0Djjtsz7aGfIEsAfKJsHH3GhopvPXzv5m1y+I4a4HSrfW1BO
PYdN0kuP+KIAbQ+/ipemk6qDcaw0dT1KiavRQmqwYI5pcGcsKgslO27G6MjYaIuE
C+5uifGLJ2/2w6XBbjwVYeBwI++JsGGfiouGhz4idJGw4txlttaOO1zQ7U6VNd2o
JrDW7BKoF5PqDEH+R38agh2R6hA50wdtopaE//qBtoYDwDqaOzT5er6HDE75NRYg
p4GNrkig1YB2BY10ZByy1UnvDtbjlwljufiFI/oY3tsqGD502qQShePorTSavBKW
pns+euSH7UKRdZHWFuMz1EAb199wJtMZesM6mHucWaaroWaAzGpnT84qdL0fKO1f
YJd9PMHRxp79USmin/S6NRd3tMI2RzOtcrF3KY9oDmDvx36g1+cARW3ufGew6cHC
u5G34c7sfLpbvBrWAU3E04Kwinsj7LURPhgfkhs+P2uHO/9wn8Tvu6Ec3cWsjo55
Zz4cvronusArlu8YWdfKaCTo1rzT0RGykVd2CiCgrpBZAN6bgr7KkwwGXpscarqp
wIJi5ZNo/qUi/0oAWVfda+0Y+SCREGyjwYO8xWz4a2p7IhvR5aJMRzrBdzQz1XL3
JeHQec7IoR1ZxZP1HdiN3d4JODoopaEQ4idOZRnQ3FeLP9ku9YRDKQrRiCe3i44b
rJNSZKU1xLzqTPBCqwBwju7yLpe4JhXu11f/s+u2EvRcGkxkQ2NmAV7+ThDnH1hS
lL1hUPfLOx55neBa3tFxxdI4AzpifPS6FjiR6QNQvm6UJQSf7lC1bfbprxbuHChQ
iQC/ZEVOdM6gmVlsuriiOhf1ShVuEuVwQhIzB6KCEHl2hMbHQe7VffQ9+hB4UuGt
NMEcD3VG+YlTFYoX7tNexIHCFiAMkyp3dOb7fB+MYZEEsve1PmDacXFW567rbYDx
aKIqnQYX7z6NgV1hYwpts67BEIdC/VNpCUmC2k9jDndPJvh5Q6Xuh87p5prkjavq
WpDgnAGacTB45voKyLJOkH+7R/JPp4epmFMa/sBBXl4Bfs5bxZzDxIIUnRBwTkx8
gCuWGI7bO4u4V2gl9dkb+GwupW6TvL0w+mxZtZ7jltQDcoY4DWk/hduD3q4LF1Vj
8KFQ2XFznSEhc8wSYDDtGTyPlRTTU50OR1IsZPKryStLx6CK4ewxLMgISklRMwGy
uxtA7ATKC4ybyai9a+gAKXjhuDYycy2IjdUKX3pWiAB2oVdYjzwyDtkZu2SGqk7H
O9tWUpNwjk61aAKN2UpcSzr8WLq86jIP3V1bmyZj06eOm7QTnBW1p8bFs5Dgp9m0
gZe1ahkBFVUwD/VDokD79ISdL/Tl4MDx+nehV0vCI3Q3EW0FVsOcJD7WBMhOgV3h
vmxhNh93q26tRspsZAXBFc3nWY/e93X9qPS/OquHqLSDYXK3UOsR3eiBgE9X3HvL
u7pjUbKDA2wvjeMwygHztwBQhY6AlI6+as679F1d/HNcb1eowNMttLzsmn1c95gw
oSL934/PUqIOADIzGI7J4jRZiSOMMHCw3pu1u2v/zwRse3E/kZiPMeB+oM68bvaR
fMAYnVqbO5KRU+BEYrCFdZfyDwPUMig6saBFk3z6mydz+2n3rx9/TEJj/KRBb2Sv
m4htbPfcNue9EOCAr0y2SzSQXB9BQv9Z43ZjcfPzTB0YCOFwxeO1UFxY0AdaCsRn
ag1t1p4jhOONodInSzRh1uqYG0kUGVz6ZMOVX0ROIDUNYEqLFkdjC2GShFqwuifp
On/XudWYmZfK3YKw+AuNFQWAMV4JoxxB7El0jq9Lb6/Me0G+R+dIE7kGFTUyPL8w
+0hSZrCYLhxBtOjfVUUtXqznnoMOKi3Ik90YZZ+WRkfTb79NvktboliOrtDfn6pG
NDHRLgcd7BT9kQHzN/lWi1IhOrG+rBeJRLGa5Vgb2MHfJZLFVxXyd6ouMVwxat8v
zc1ZdECCJ1ouDecZgmmfcTdtWr2MioNOV5siqawaYKOXfg33VvuL+aBLqQTAxMIR
z7D8uFoQvlYhlbqH0jZwJqz6zO87STP5PTnsxiD0L60X248sl+BwjU0YY0oapGBR
U/blvybSWa2LgLbqpWT3Qtc5Dpc3a3DFKGb4qal6lBJLOkyxQVDo7OkSfzbDXHzQ
tfaF8JADP8aeJPbVaZ6goHlRJc080sq6oO2J7vXAYcq8gLXCxy7mfDQ9a8cu1ifX
SdyUJ2t7sUfZJ/E/khKglp8wiKwA54/uAtzTsN9h3wdOKROKzFDtLkA5YGWGC1XZ
Qk6pMcEbGEXi84pB35ccx4vVKxb1tAQp252mn5odmA5Z+mPV4JDk3Dke9lXjlITX
zjCcikA72baRG5VnJ0oy3QDo1H8fBzpOEXbZgm5xF0vE2XnOZozGAk87I0N3zVEa
ASIO6d+5ACPPYqKdGPJ6/JIxqEhGQu2gZpNe9q+WdSYrHoi4fEftrGeqBp5L1Oo5
S4gl3wTnA64NfA/8Ylb2QcsCwCNrrmkp6hieJ9tNjqTes0ENFu/QdM2mvYL6dKjK
r48p3/p9E9CA5Fw3hW872XPfEXL7C4jLWpWWYeQM5xEu7UlQLbO2C8B4t/9J3MZM
KNpAQrojvh/xAk1bqn/Q9/tbSiXdiZJbvO6IHkdstFofd5P9He8om3KpiwBU0Ye7
+tGdjpDPMt1ZC+PC93CNX4nTXI2dQCU7Tismum7M8UlkuvBk9rvjmRknTHSnbzKp
KdnyIXgJrqK4kEsYct/d4hPFoZyyceDelbBdq403ZpLRsCD6u2FCH8f0Gg/yf1+c
VWGAX+kZPY70JRaEcfssIicGUJEM+q5AZ6Vu3sM2fL4k5KRiRtJVEs1FIZOQlvgO
RD0nFFKS8Ij7wrgbWVjR46OY6oUWpfYzFivGegC95HJRnN9s2WJnta4U6YfVmQQ3
fu18MaQ2+mVBWnkgaav1y4h6ohIjGRQGq10LJ6aogKMdAOPw5w5ow5BVe8rL6Jxv
Q5WabUv6grY7ne0bGj1uZGhHNjhR4TUu2pCMRJH+nsu1A4QE8G9ijS+IeyE8kEzE
H22RS78yKVGpgogkx2TRa4s5wpn3xLnW5oRSGIlZEb4b+J16CgoSWqsej2J94/rx
+/sZkJjKPQay2bLKgVOBVpuN5K+bf2wpBv4m22lA0cLy7EdfCgXJH8c+eqrAbIcw
ceXeOVtTs02hSOTtknVHvmF8aB1Qdw+FveREUMsso6owrQvHc8/vxGJuOtbvTXrs
XNsxGwW85OQDZt2iwXVSlsaRaLqOEW3KeA94qu6ZHE+flLOxaubGC28ps+Jyx3tz
b8XfIIc53jqO4wVxwPkxwvguxp11yaaP4bOxjJMyHP5sAwNrawTSpSlv3MG7B3xs
G8wzjaESPgIi2ebVtWzJth1L93tCxrJDUYLXzL7uhgNKSSleVbkTTZKGfYLJ0EXl
u3duZbmptc59lPIeYtMFEaj6oQyf+nKYEfyg2iIuRNOYr1PVGFN7Jjp4olC4jd6g
VZkbSj/gkesKzAGoonZ78CU8G2qnR+lylQzoNevKClzCifkGtdvDocc2f4Eq7nYh
Wm0wktw4fg6RcHVoMde5ziqjR22yyrbKHzAzgU6zbLl0Q8lIrAi1vgemMkgaPKs1
CwTVQXfG+i1pBnuDAaUgyf/+IPhKx6tXvHx1h5dirFOjGBkGVz5FgSnaTcGPoAVa
6BCkxr944W/pEcZtCZc18UXTV9ZDn21Hm543dmPADcyNtLhhGCmDJT72Bqk5Uwdc
Un10ZRYXMCqd4J7v5FmiEd1dkR7GhK9MCIu11hFFvLyUNAg0d25n7/Z92mvTbywZ
9xM7JANO3Hh999E/KzTiWl/6rH/GBCnyYgwpcirLlI38gu8TgqpMKfySxxIZQndF
3UVevkw08BNl6VzQuC6nr/0sJXOvUsZqO1oc+0Rl79Sy/qqPVi8YN2ZGpYeBdEXW
//RXzxtW6YFYst39ELDFtJfPMWeBmhtn+uJNeU/AN6F5PLWf3lIi00yWfk97klcb
wmKN8jPpOCH1v0kOIgstWGmSrJi+QYRLbuaJeYKGfRM+bq7e5u/LOx+my3Cu/fwD
QruxMbkyocgHdi6322iy0uKtiYolpwXVaCl/YAuu9CTRGB+69AeKRXAc2XTKG9Wa
v7VzJfomVd5xQGD9pEH03t5ijkxlH7KQ7aBjhpdpbYE4y9fymsR2DBg2dQKcNYEN
iw3MVfBbARlj9UzbNttCpgmxqdW3L30XxiCFdo8zzNsJNwFScD4tybR/ig/K9EEK
WzAFsVI5eNM1HSvCeglc9V6ofScY6prrBqb9fdcgQcworgka05N166SIMn31erZ+
eK4KpNXtaSeY+S73FV67mPuo5eddDqnfrOK6TNp0yPV0yXyi2AcZe+NbRu6ijKU3
iO6BLPxiEbLtvL+11ILqSTkMtwMKRV6sR7+4jVkW7wFoIeRCOsL/7QTdV29JDMpE
RHnn5DruU2ooo3jIMoEAzO29i8FiJY5TszZVudh9dxEfxNC2wunrkacZUxUdDJnA
vvL0J6LUyNOSGd5wdt7YoXBNJZwB+Yzgc5grrtL7260Jx25rzrPDanL71pUbPDhN
zaQ0kN2uZjSVTcweGXABR1g9ZQyzay09iVfNTmkaKANW8b4cpw5Si9JG+iqSEZpI
ajzDymECRgxj9U5jtcJOa1IfCn0syTcWdMN41YualtNa670T4Mh1/wOz4FludwdS
Rj4aUVQOdmyPKJvmsUoqPj2cRJQjuFZp4LB2MPuv4cRi92yrrSesGdAZbp+xI2mG
vYhwgPqWj64MuODMrHfebHSEQWI1vqEBU3d/sjO3wS9niXur3/mUyZww+Q2p9zQr
FehbsJt31Gmc1t/N2db7Cew/inXD8YHX2/kvAoPhmh/Ar2ss6U8BbNiKFNmClyjE
sPWCi89KBuGWxNpCvpaipD6chvTZ4ecwLMnzt9WsAFIkQ5gxYyMe1u3Eh2ueroSF
KgVE8nNN8xxSK9iEfOPS3xpxs4McBayggaKxoq9b6mXaPZXZXOxdY77dDcR4ixMu
rm4v70KJ7fCaxwR81S81t+B6zPpBEmX45/XHmyMoHYidNtipbUpwQg299bOJluG2
hLvteZKZ1vwt8PDWSeSylcRFzf1zENH9K6oPlShWxPN/A6RBoGgOqUrxbXigip8S
p3LmJiK2m7OQUx7AgyC3eC4h/34Yzpabx+b/7jD7lKEIX4rIHjEWLtDlMsaXv8Pg
0AHKTUnGCKgW21ie8T3jQ/VP38nx+tVLWCGSxWuqIie66ZJI0tBpp4zhw1uptO3/
6cTg0hu0Xov+p2472RWJiRYz25JXjCCPiVl5kTu5h/cEzjezoBw0MoUwMoCS2Xyq
E9rDVX7AF3ge7ub3kT9sRXX/126XgjlPI5IPRSpS7Rc9RUSNT8+39R0Ve3FtRuH8
z0XftM+80rs4dgCYAuRyPPc0XXxe2IR+vPorLsRiM9ESOKP0URxsm7Q5TrZnDTDX
5hChowY229S2OAAtPQ1b8Mw581pNQgd4vhY7LvU6DqAPMJTi5/O9fqlP1Tf83hy+
aZOuKBzf23NlpQaiXL0i/whnEeB0sGN0S2bOTI1RRh/+TBQbFvJKCjQrN6Ulmea8
58DZwNAVIgCrCLiSVnU2d46yy4zb+1MnU2NthzxiDP2GU8IWxQmnryi+iwIKGCze
mDy6V75A6oqtw5xN4iUz443U2Or2r0mBqX71MDEHsuGuSmSNOOq8gk1x6TkHXqsj
slNwkSGTyzOgxNF6xzlkSVlSN1W5I9/yNmZJH3G0VAdhDjoxPdqQ0AlEuedzHsMR
L08C53gJPwedAjpLk4Q6WMTNZYwo35GOpw/hMc3Ho7M6yQTGzl5cVGxlpcWFsFl8
fpbqi+yfw/fq4df8jmjscqwvi0POqyqT+qasVjUmNbh20k814ipYlWSK8G9KEzl8
Sy25RiEA9HdvFnDWkhZ+Ds0SDDhN3At3vwSJxCLH6JfJYUdXYmPYD1dWFVExnUA3
/Xqks3NCLPCzEsNwSJ36ZOiGGMm69zzv3RbkDZQfgG1D0hbfOl8Ej92OivJ+XYAT
194rMS9fJ+qgR02GwiTpKfSmEZa1U9Z3l9kSWn5Av/bOqor/nki5wnyo/lIxDKxr
6SPd/3occ+8FLLbC+6FoJalEhZ5O4cJkAzD91AqfEbM0DQ/JOlvjG9raGkCo5gA/
ygs+R7f+iLIkAU91OkNDKpIUC+py+wW2BVluhE+s9SMylFiO6ggn2LVmR1w9abpk
POCmXNMXQHTtGrw8NxRSfzoyu/AJPLxHMlL+E5NI0ufWqXlRKN92EL/SeFBuSbNS
wRXTNHLrbjabmlSZmzY97Ik/sNgAbSzuChIu0+5I1/0N2OLUvYxPnl8LPcl1U9qn
6qcJOgnA9ADC816NqymHSHXytf13LHSqc6xEoqtPtm6tz6DXsf/btmA1O+OgLNsd
4e2Pn74oZO6LVo9EaFm9tOtVKBhow7H+KKx/XXmd2HuIQgke/czJioWCwft53Vao
ZGACpFrBgw/+bZ9fVS1nHeuxbLQUQ042GLu2GEGXgoGD/W5T5AXJhSbOMvUEFAI+
iW5/J0O/uQBbaKuk5gs/8YWzoDSlmi8w1uufLQDNTASkCJ1HDAKUr7fXcbqzEUUQ
Tml2DFnvpn8hFI2Ob0muJ9KlBnGf6G7X9SLmFXhTIMPvZS5Gu8YExQpZtLIdsvxP
1KgugsDDiAzRnUtB7NSDCPG7tMhqf4MGFh8PJvmsYnjJgUgsZPUDB7DnAymNZleC
l+PikykxqT/iiv1fm5JOqrbyEGRJlkodQZPyQRYQkTMwwsH4sD1JJTNicvknyA2n
yv9vBX54Q0pN77pZ0bgArcNFQl3FsaI+DHy198Jb7wG+02IxuZjScNzVzWFL5vvu
15OhzSqrdgGHxNv5KLzJMlUoxGV1bIrAySqN9qHOEQyK7isEt3EVwQa5+hc2LazD
w6yvaxcD4mO5pL+RIN2triTbiHV+4TvK4SsTeBzyVjKlAs6blhkSO+AhdLluT6Ah
O0fGKwe4PEDqbeHfLyoTRGIc1PLHhumk92bCKJ25d62RvUYjAyIwfRkWEISUSMEU
9kimREX+I0glsRTBV1Kvk59XE6mS276OrZlS+4tgcgztQZT44ecUfxehVEQo3krz
eNZ8fjC1nk3wEjiU4+Q8bVbZtDyFHqZgtzsPDb6OIyvqzbR+wx3cWZetSo8Z5Kve
VgEiT4DxPAqHgXAEPjwj/nKdX3Oneb1Vjj7tS5BxeVRsK8dFqdMagH4Sg91mWRtS
elM4DMt6AxzDfgvQYVZrT29u68FuNLW2XXQaDwStthuJo43dOGLg5uzXqfO1vYhk
RThPAR49ba+7Sr0wZil50RBFL6z6ruenfPenSnVpE82p9NBksJjz3RNpyeiU9f30
XpC5q1HuA2sdywGUeTxEHsdEuxVlXGdSZZ0FOTKksFIk5KII8A3uwNduwwDb9uOM
r1jITdZ6/Y44oACNc8d80N/CVtFnDxGcoOd6X+86fUIcHy3N+oPhAyK+EUI+hEGM
6Nx9hNXv9SvCgzA6KVUlFmcSYtTUWSAluxXPMIQwGyi+SiF5g7W4LWPPPVhgJ+Rq
37dHClHoy08VC888rzLZy58sHykrh5wvOU/hMv4B4t3zXnUcGINpWrUtAKmiYl+E
hHWRHHWqtYp+1DgqLM7cHPpc09Diuwmo0rutNKqOe5ez6z/qXaN7ibcK+T29Zw71
1Y0Pokiw7ScTM5qHwtYtTnRKvsFmv51hHCbCQnyK+kOeu2S9bWw0dM3UZAhen9Hi
fsqEr7fAM1n7Xwa6BlNctEicap0r2PSWTpHfYnH+2HL7uXN5JPtmw1LNFgrSKN0I
Ex8wIP3uphmHly6PBNOTOItK4SOs+SuGBwIurwLIXR6+0amfARh50G+dFckNeKMu
iW6Yh1zo0Qj7lqRK/ZaKcg7BhMDuRE/u2H0agTI39KtPUrunm0kutVjV/WZGiDJs
+WtVWuXaPH9OhFz5AZsrhwCr0oH4imJjELCgScwfUDVQ4L/7QWEVNmUEkCJKbMEk
17reALCOSyur3mUO3DM/eO/fo2p72epj/8jSXwsfmXdmkQrpK57NfEKadoAfScvr
SxhJsH2HRE39iVjsFEkUIPXKVBJne0dXNVOtTaHOCfS2OElznb8KpUJEh0TutC8G
a/Q/AcN2DOaznP0GvduXPcVgmoQjMkRIJUZuHa092vyMZ0gd/DTt1VTlgjnXVPfp
PFvE57LtTNxLEyhZlLM9vK6By+kPe6MjsbA9cbUqHk36bs5lH1ETlF0hLEuF/OGA
V0flOS0oNiN58g0Ee4V0t9MSrpicf2DGkzy7JlqwwibGgHOp8SUCWhKt/GenejJF
dRnXhGG1cmWbP3O368QkxN5OKFIIwDWOvX2FGCEpZxA22QAulRATS1eX349fQiUm
laJOREvlPVGGKiREU6WOBZgl29MH2LpfHbAwcCA7Lr8JA5x08dWnxNG3nmx0OTbw
CiOV76rnViu8X2k91Q2D3qWqOeiKW+dtL2cVLCtm+M/vbYcx73VxvTOHvocV5Fj5
viCY9gQLUQSDJfos6C7Qgy3usQDVTCa2o1lI3TFFMK804VlN1q+h37xTFHXm+DF3
pls/OJzpiKD7VvK3NMp2+SP1Fad6233fKQZkR2REjv4IztJEb0+SsAXv83+clevC
gIIjRdJl5guoWt6gAGMis6eCpFV9ZmxLXXP9uvgFdhWDYlVvAHDN/KVqkTmZDTVm
FzCxG2e8xmjghDyMcNLyhwGUC6+w2B2Y13bWHHRkNceN7qz1U7Cpzb5ZZG/x8wSu
bE5FHy9eLmOBzYCYXJibRXWr3bM/jnYKfT0DrWYTZycnpT+8xZlW4hgrVQtEiNi0
YwLbu/0U3bl4z5sEVrJOVq9dkYDljZ1MLY1aVJt80sFVQmHYuA0Ab9v60zMLLHY5
4gVsnVP9oWSe6nc/dfTRLnxA7qA/1mvt/vNbYBQicij2yXRQilIvNpGe4d4Q+M0K
kBpJTXEqJnH7ODtLHJcM6jDbNgdBbNFIBW/6iotFlruas9BQ38pEYwSnMyemecrG
6e7xZJBuPZu0BUKiuFwAMbvMHfuoAfKTBcFvpGKo0wseSswA9We+jIzEBHuUanhT
mU1Etb2oI71hai9x5/KkpjSNQjvy3EA0ciQ9YB5nLILpZoPca4c1cdy0C+dJVsZR
XE8eOOkWRjPNIG8KgYk4MatcMXXIVcuV1fQiJKaYpH51byM4Wz67THHSfWP3SGMG
+jOaAwnD2OKZ0Px1UZRB6EDjtTSzIIOG8MNc8dt9O2WCwrVyN/FkxV/QdfpPcMNV
J3BcRvj0OISabqKKR6irIK7mwHOfBuOSnbXNO0dAwhGAlXazhknMy254ZsBBJbcs
JO7XWM1C2N8Mbmi9NryfyZc9rBmYZseHWPrfVK3jEShxz1eYZckAf4o/2r4EjsPD
0mzoxlN4MKPiGn2KJ53cmx5lP9ykG68M7IY2oZNPIXGXhmKdFfRln40NvsJJi89q
bGlXenKkkuilByI3OqJfS+yNhWUE/l4pAE2LbyN3W5UGlr3DikM1wmcpKsX6GyQF
3Y19UVyBuAS8Tss0MH9WR2Vst1OiygQrRrEOXI1YUxwTjkQfTuuedbxpX8WmTmWP
Ee6Ng5banpsop0QliYsQXeE39jvNvFIrSQVaxaTbKtUSw274Yf+8+2LBb/Em7G9S
PSEx6XaRcUq3ZPDB8YcJp6iC2hGZJpO+RvylwuDkvRIl+wptYCWKZPXi8CENREdK
9XdrsNfKZQjb5rFwfZ/EgwOiQWu0G7E1LjfsgWfWMcHT4DHS8RchasfcDQbFQtNs
2HS825K9SHWfFsP0faA9a6WNjBMn0vu0S9JIqM6egWCpy7GaSE51sym9mt4DJiDF
yAaiTYdA5UzW+VQ5SEiaEjkoU49ota16WVcJg9LojrO/WcqPVq0kdEIcKjeGOWhp
WVbCJmLhol3sd+OulFHorDQYUcCqg8slznG/pET4HJK4JlsmwhxHQpxhB9mOBDox
lFrk1FMlleCNaIoomKtrWMWSZHOGq73FaC2YgM5xnxW5U61aqXg4YEOHNUcSodZ7
29OXJmoYJZ580Ha18xHKaS8YMW/RWkfEK5wTmszT0XFYm3EUgXYO1c3mfBp05Kty
V534FA+BvFVmDTW0nccO9NSGwQzjL6Sq54yUW7GgL1ochxsOsOPLfYqnkwQcqctc
ZwCU6Fg2is1kJBswNK1/aUY5bOTr0iHbW1zZhnfjDXFx4lYl9qAFRnU98MOii+1G
ZLT7gsxfAAS8XvLpJMNJS+N0R40LWDl2NPKAYeYOmYeAe+xKzaOdXi9dksgRXxpk
n5Eygz37D5tCAKv3RFGteVrcYoqfAdAedTH9Nh/mjGm+SwE3U3J7wZpJC39LBhAS
CzqdJJ3qWyeM3sqmFo1oABFdQLMbHVHmCn1VS4O+V+59q/1yz2dxwDQJ5MO9zD++
9kFxu3dzlPNZwEZfrUgLb+kEsLnYZXlKZKnZawaTknGjjDSQpBFi22uYg+E7QY7F
7zIEMUiBXCe9fjdFOs4Fy+SPezzCJRlHFl6DnortdvurV04IHdYUd4mu5hKhBiXm
y6sT94r2HryPIushi4LwIggLPk4W+DpZeBnkEGOJpmINOLUMticMiHQfGPJ5sMBA
Xyf4eu58A8E/+6flk5jRAcjb/QNdsmLiPZnAlr26K7PES+g2N4p0eCIOJ9Mg2ofz
O+83qe0B9FiTFRL4MDMu5b8qIwNiQI4dCGP10uc9VhPsnjAEnwk3zb3gaqdkyrWX
wuRDsvH+OiOXU870TfcxK6VnINiSj7wD8Y0mrSGxKzVH9L1fzfMOXMYDAGwuB0uo
Z3iZ90t41UrfWI+XP6YGhVQlk1HdxsZ3T7/+xMLg7g1b2YskQ+tI4LztGOo8Mgoj
O01IGd2w8KUuUT1hq5CIiodJ8emBIod6bme+bhijzl8o7yJNznq01VBIZrMwhObn
sIjbiZF+0RDMzHdpquFa5OuexdTrrSdRYDFBtEZ1zNlNN5eGgmi4hVIc3tQDhs3Q
+d/4O4L4RBDEcPPMLp73O/JAfUA+621LUXqJvY5DmrL3RE6sA2taFlsRNygE9/CE
c0lnj1GxdoMXgRF17ibIKauufIZm48o1boYpQdXJzyuR8CDelN7nxSQEEwFE40e+
Bjb8BbZ9CcRPN2tXK+EdIvFLg7BUdzzlgLH+iy+nkC1XmQBO/3t0esw+OYp2W8Ey
bCu8htI4lEk3ASaaG3cCX39MbvC04F2gWO6S9gm7sXCgk78x43kfjL26xLB3Zu1L
n8Hq6NvbN6kgfy8mV9D5mGz9FFQzPWBOQO5j9SUfTyofL5MCPcOzhhhEngEZh6BS
3ud5s04bnDpHifsvboDYzGN7vKDTwtqDq9OpAVT+0/qTj3OkAGzKD+w+sZlZ8jdu
cFBgdijYmPBsksv9xARbC+AAmVsopxji7pn9GgY00JeGhuWyv/67lBvpWKX6q5Ln
nx3PfT/iNvPuXNZNiDdUxujrWrKWeGXg8VD7JKaQmx2RCxEs2n6WKbNVG8wkWUqQ
cAccBA1s+pLU98uH38EjFozI2dQku6he6MkVdSMsGUIIM2kseS982o9dk/qIlNZw
G1YnUI+H5+n7uWReHExSS7vodRtfY5rsm4eWnes0ELhlWufjpDu/ReYubrXbXaSC
JtKM+yTeCBJ0hG3SzyCUR3wDe613lyul3I3scJQmRJYrGdlAE6cb2J5mTJzNMQa1
m8oz0l+CHDGLN/wcZPw6D/M1BJG/VxDSjbBOkshqUgOxPuMv40+ZZCS43vLuw0Up
VAQ68+jVfMUmbphFMSkZABXsGtlEpUN26lwYTUexj7lQM9a0aCixY3AJVRPTqrly
XiVGuVYf7EI/07Cwn8dBrI2qF8LlV9Hb140x/xQzSJGMpYjID8k8aeMyUQ0a58xX
UHsszTv1ixyqTayOf8gkIK1WJUdHgvVq67j2KaorKNGi1HEFk9E6LwYOA8Vf0WFb
c01ITWCxk5R+jBDN1VaP75SyONNoOS81mpagA+vLS4sKQtUcVVQXy2ex0RYL+ynr
CYpWaua4em2QcT7AA9Dyvi0oJrXYhNK2kb9qyrgFYnPgF9FmnJSgB8U+nKVC9FVS
i0Xv6IVINq9a8klT7i8WMWpc0KpMg+4zso3NMShiAqPvO7DJze/t0jsx61dP2SaK
2mO7GGpF5hqPlCaZm3kz9ikQSASU3LQ7R15xL9+LR3IBUcaIT04bzK7d+nUCJjEx
Dtoxfxr1tJOQxyuSL4sHNsF1yW1fpzc7t/LPB4gV4PVQALzQ8irWo6uo6EPUF+45
eopizBIEbcYykczy5jjJrfxZHW7JsEvTzMQx8ylR5ilO0qxU2nKTwGw/Lc8xkM7K
Gsm7tjfcKc1tis9UouODhic7eT1MrcXWauFL8PF8pUZpquQb4AL3ItBTCwaMgw1b
1HM+bDpsbZrHdUP7YqSN9H/LCjJl18Pm9B+md4wsSQ9iK2iaZZVqb9ZTU+UDgjCj
6fkwaaAivVSM6XIC8pven0mLys5CbM7WvY7PEG8tGF81joovEURx1aLrfTMPFGPt
YmsEYOTujui97aYTFj+d7rkKkiIY/kb0TIoddvsXIvIPnHnR//Jhw0QoE7wMO1mf
gRT8tHR5K56F7K/tnf0hbOIc0KOcVKSFTxS6DdyvgNNfnHK0PfOVwKoVnrHePp+r
c9pA4d5qtGwmJi2GB0CZDJ7EF5ePJXxViLD3dVjH3IVltXvhz33NACBxHLdO66nF
fxzvv9jaTXBbu2ohHDX8zmgc3FfWbZZx+6qM18Yiu/wTu58VpM/s7kDm2SpiBQAU
6YReQi3ihQGieMrVUkfITLjzGoUqoc2BN7OjAwGxDL5eSpj/xrq63lcMz9OauWeY
VJLiYHnAn6DRxvLn0jVCDv6T+BvJ4qvASsWtt5m+6sPpQG0h4OTXl5s/RemsfRHy
FWUxKlqRTl0jIVjvDZOHKArQgVgCP/Y33+oCQrbL1XJUKYDXPcmNuJs500Syhw1A
+72pKSS8J6lbN2qff1O7DIw0Fc6m2uIayX69CixaUyWE2u6HWXDCWqQhjLIICZSa
Mi72qdwld9bzDTdpoSxprNkyUPseIO95FhAqmfIT9gLM1qbnzg66/PSFseTUTW6a
FAwPuRk8Wwjd7/s2LVWQniFhCsFu1Ylxpx8bokcDY/78IuMxpJ9HZzz7xyqKDH4c
RjLSfl5ROalDjFstF58Q4WZDIkOAPNRz+XffV4C7gwXy0B26CCkgT8ZH+qSY2kEn
cMorC3+VjC17ADkcAz5+5ToLSnIpOwGjw7hz41wfLtGX+7a6/avydVlLy+hKX39l
l9tgF3z8gwL1YYiqBAhYk9pPqfclDsypjUdjhsLmunY1xeYqvrbbQcR0HFa9e2tl
Rg+g2rkequNZZE65NHiq1gKeS/GdFQRMa4EMpouM4IrAY6y44aY412c+Rk21aPgr
GRdoBuOJl/EUdMAjJzmn3rdDefj5uKWBFj7CL+dPuFFDJo38x3lXxBttdxo1B2Nd
f+zmt4o6rk8ekFnKwliWS/Ni6+2dJZtF3MfvR1jy0HIrKbHiZoVWA+MbOT1IBht1
Y0WMqXIvSGRsDW+V5FviWGRf4uTC4C3DXpteX0YHCDKjUsYQRAX08dp6k+t3AsLd
9SH3CzjVDfFEw0zuKTYUItCC20Jlzmj4rzdDSyHW8aai8/HaVHgsQ3MpXL8QgPas
TvLKpCxfOPonCRU/od+LbJHKDCZJQEMYEbJkdhP4VwW4UpRVUYy1wtf3voF/BBXf
r82YIX6DdU9AYrDohfebI1+p56shFKswQbIpFn8tCb8o4pfeaED5U4eeJUdMinIm
UEzCAMq49PwpPgI2iBq5TbvhOo1oenCyxeoeCat1cSuD1KH+7ls1EwAY7Omk22Co
/HHKvX2C+lPehYMrzVgzlHHtOB1lq5QSTdCqPrupjaUbt8lYyy5Z0lovALJW2UU/
RreeuS4av/f/YT88UM8/5O0jOZkfBdCqV0jrPpAyjTDh7/MZ+f9R0LHJIJxt77Dh
pyoq7nNAxSZbANzkE5gnWdERAznONzRc8Pn2FPX7RPElA+LsLW8HieQnj41P7olj
dbOwG2q8w69VHi63YNEsUhXHt9s0tSBsQf+tdLl1EFM83GNpgHY8mlKi6XuH1v0J
LIPqh9/FfnTyXHHhcRD0Wo0b1vLGBXd4Lf/J6fNtmSjdyK3MHcJiwVn0xX9dDr4y
6mG0ockJMXNmWQizVivlMuK4c3fHAIvtxzNf3BcDd+hDje1v1Uw/SCA4tEe79kcM
1nsoljHm2syG2KqGBPr47pm3olxQIKgasgHiZSyH78EdqFfx3BAUS/0wVcFKybsu
tgIQ1+bWlAgeJgsf2AL5PlrJ/rPJiZJNdxoOx0vkGXMMeUsvihAvG+ASNlm5MBxz
H/dYsJctVgJlxXoTDL8kMswKinGMB4uI3faeRbDz0Pzhqz0lK4+EP2Hmm4pORn1n
MmsDx5A5Du7NmPNoUtSq6x66Hpi5YbuSCFfomvTNNPvE3icvDILbk295pWMj0UhD
Dz7WnfCE18zBihEntxJKwZnEw2zpGLTK7iPf1xe0KjVlnqt3okP7U7kdTu3tae0q
f2WeLDMIuXpIUWw6F+EKWAFqUdUqdT1NOqP3fuPm/zxcTdOVffhHUpWRYll4J2wi
7Y/B8+yVbV1JcrlX7/HHZ+rw2ReCrZBCOzc/ATB992uyyi7a1jeg1AGRhUJMvJDL
lGHyMsHMvwyY39YvUa+eCpAXTFPrYANVuFQ/0ZO79ez5g1rlG8o3H8IDiDJ7kjYb
6b+lNw4WUGbsgIlosBS8TDJX7w9LhwTogCkw715+3lC+fIrP6pP3+bFV9iRjNPhp
zakgaKWSgHuBr7+OBVUdyv5ZOktQJp/jIvwGShzUcWLi2QDveMq/EGG/+/XC58tt
D3RxiyyZd5CUvVLeMQ13IQoEicgel1tgwaJfEKi3f2/ys4gExL5XY9AhgiIQBnLP
R3JjCb2qRs1ALPmhMNNagSDhu0ffPFT323/vc7HljtPtw27wjIk2xEau9irocBtH
BLC54hA5coQE5jwnB5km6ezMQfvb9a4zvNq1dYKUne6x4Jvn45+3K7hqL9bOm0eT
CRBGAmoNXeaQqqTYgn9ij49ci+M+ibmKez8R++V/tV28JS8HlYMCc93JxzWMOava
rTLV64nuMGc2Hz8g1NBOhXhElhWGhmb7K8utzNPmwHoXO4zyxp0lJ5/KDNwYdw73
7fg80LHFXWNhqZFFEJ5t0Vcvv7GuvcS1JcJ5URVcvmb0RKSmj6yX+L+HB1II7ZzF
O99kahVOLHI08fkQe37X9TDYVMAHPHJcGRcUWU0XXwiNTCMwa4xETyNv622RGsOx
kEMv8v7h2kHYw4QJgamYB3w0O1jBr6tx/bGkLjl4vJovawSryhYVvoX9hAFpB2EX
XATgLLh4OBcswGJnQBtEZFYC64CD5ow/Zi9KpW/LwVFFbKHvNt2TrtKulfJAchoy
gsgCuRPbfR1Uja0phPSWPiZbcEMMU5p4sghYUaOw56zyqRnFpteDMhG87hygWlkq
VPit1L9/DH1kc5ZEnR0CrBiLFYCmsZmT6J6EufDricQrYR5rv7UgckZZgXp8mcyW
biaAGAhgMOfsE2CsiIoIBFWYd1QAtDX7nn/atSO0Cc0W5j87UngOynGPju8lu8K8
7jKsZYcijcvVvA3GOfqr4gL14o2uWpTyTUNUaTU6JM2MXsQH4gdGj9HpsDpO+s2f
Jj0hHe/v7dnAt7f8QbHpmaL2MnnHlDb10DbhzVVGNNz2ID54tv5hovknnedVkS3H
0Ae+h1CL/fjt0tTMQcHpuP8MKowdBHR4AYPa3yq5B/AegQOP/c1B+OMfmkdqpd6K
ulTjNk1PNRWr+p27J1AFF7wZDeIZeB3ZuI1AHhXMLMERkJluN0N+HDP0NLOSFa3D
WApOceJwAJv41IoKbuPq5IA5IvDp54j8A20DS5KrCuDQsM0LisFx723kKYu/6zz9
lSFNzWbFcgDUAWzUBaQbNRLDmlkB1l1+sNI7AWHJ1uTE50aX1vBEw2BcqMujXRgv
dJTwFNyXd0LVMpgBOHUIHonYGitvXcy/aiRM6xcco9gGNRmiShtMLYkf7bXW6ztU
uC4OXNq0Jbbm9yK5GkQPXzYCwIyUTCjw6MwkkC+mvuknfDfCMVf0xiYxUIWkHsgm
pwFT8AatNSMZ6dK+cnOSoTonZLUleMJx7PjR9Gwt0SkP6ZpCIS/1Ta4ZziLSzTUD
NZSuaBLIFlsDeEiL1+qSjaMdbq/r7BLUumTyRUboFvGwqmFG0WyAQ2Wvz/pLzlU+
YqEkyzkHVPyHk3B16f+/SwN1QZCOlFzH7bOZogHIF/Ydbbq+dWaCXTBkf97e1lOC
V2z/rBCawXGDy0963GhYClwFDs9/CU4ZFlEDSgVuFSWgpSzASdQ0e/duQ4fgfk/g
JFW+jvt/vn8toDs56/NxpwzAXj3gHcDA2Zfp6v8RLJF4rFkJS+PUCv7N84rK5xTO
AY7WxKe7XX/qzHxYb4CdwyWONPDuNzQRbPNawHx8YQJGY3iMBN3wVwd3jMr579f2
AndQhxZ/9VIn/V8ycDK+W8ripFkBFgGxXc48E0cEWF+f3i2/aS/iz61qj13HTUNV
gHAThsBCFrcbQ3vRIuI+6UAkJSeJaaSkAgGnY54NVdmr5TRWaIUd/tHtp8tUUCgI
x1ZIYcOpezH2QXNdXvkuPWoblWJOhBY0ANnl5TeMS3YMJ97Cj7G6teVsU1J4k2MH
kIBHlj42SNM9TxOGolPxMeQR5n8sTnTwNgt0/8tYCG0laWmk8auYBRdnpX2H+rMf
8TKrfRYmgnz1KuU7WkFPpKgmdtglrSX4u61tSy+OtVl6pi2JGwAVR8eGcMOUsXMn
/LmcYHeuDuwp689qUAqnwYWW528o9LQRYzg09H3DByzBkdFCYRko5rsWvxLfGCoV
SNzqbUwYYC8cAvxNTauDSqdMvi5UISY1BL/TcsQliMLtkitLEcE0tmMUYOwb8vVD
VskU+URuuaePKzBW44wun9v7TEu4tWMVdtWMUpXBB3LFe2uZClajZIifqV13tPlU
k2CpPL+uuOJx6TK/S84kurAwOlzl9CQtd3lk9ntdf6SYiJctAZgRoyvwxn7wiirM
nbsUFkMT/7KMTdo7NP2YWcAwMMCuoHDKkHl05oMe80zIZ4CM7BEddzsTBRGgytMP
JwAP7Oju7UhSn4TZT2hp/S0u6Y4sRjOT6XjP81rDWn6iLbFtQ/tvVBuWOeaTXejB
TzfM0b9M4hxjMsheNFzKZC2Mvi4XpQ0XGTBJKkeTHuAGB7HhKsz1qSu+3mnzZVD9
2FLlFQVyOnrtHFPcVIjpwCCvvgLBMvCtmQ1Yss59+OyYn9upZI6OuOXPMjkqo5rF
3TLwX4gJT02N4NU2mbfHCgxSyiEuqT3fcNT936JYG7BizVUr2tG1SMn3Af8RJaO/
9XhMjrg1H4i6hZvPMo4hAjNn85NPZaUUQ7wgQb+vN0lu4d9ZnfrDKHTuSwLR0+xS
mRpcmdLxhKSptX7uT8oW243dLPbByZqB0T0ikyYX8ORponY1O4f/Yd/r+KK3AaHa
xizQvz5u34ka46ifW0mhDg3d20mcI0/1VP3zyvy5qbrssIz6ym+e6fJi8+vkNkMX
qaw+X8L0Kf+qdPqLN3vKKivg19vRXx3OeoLckLm7Vpt8/qyTlVuDrUyxgfPp1AUN
AbvzSaHD0C8/1YH1/CN8c1/uHq17nVuEckr9oYybQQ8trqw8l3FrF95/+yFkEAeM
L/Z0gNF14twiU0iJccpSQiP/2phQ4yYaq+ox4lyp56vW3cd1j79soGJiYQ3g4EsA
Ok/ghBZPVYSQw6vOa4LrkVPTxKGt+USxbwxNVZ31TLhCre+XoUyiTyykRQccrXx8
4SFrcSgjT6EciMUcpoWeKOKNpUgQVT16ox5D/FbmUl3OoNRgWNNWgNnnWeTEnk/P
lOV8ypwYAwCH12uXvSTLCyCT3FsyV8Nvk2JCrelpzvpe1EBVqZ6OhAi7kCgQM02u
oOFQZmYoMhUyie5pAGZ/q8uhi9TG2R4X9uhju37RKw/QWdIa9ykcv+YKAM6LWuO5
JUpmAR1WZHLrzSev3TqImGl2UZvd0+TYq16WrEz9eopWw5/E3ejaKNuBbS/yzr48
TCQUQz5ULC7256uRi1lqSIDxAG1iVaRmNvh8+uHqCARubNFuXUQpBde1weT2Yi2W
PixBJQlZ5tzAqLAwOyK8AW8v5cy38hKkCKoCwFEY2xpzJh8D0KRxpaUSK/YqgkNs
cMrSt26BprzeojO9/wpruijkc3Ae7E1hKR/L1Pw68wiDIjZKz6uyX0vEz7vqDx6N
FEzsuhNA4slQGw0UgCDSmSGfS/0w0nMP5CxRVShvZhybZExHnZnBeRGVli2Rc0mf
ZGDpyRldfUFINtLcTCNyU1cA6RzYoQVosJipwu1+vlnk2Wv45k80Hw9czqxD3QbP
3CXR1xfFrMlrNySW17gXZsGM4CvJ12Zv+ZS1qOOz9cM8UTwx8TNFBqWS5hKBSozz
DKfd9aiDUmhvvl4POOAElCddtH7SO5wogTvjgC6Mo1xiAYX2gJgeJmd7ZgSYMQDG
e+MFOxy7GqjQxwdikAHSqPYv9/kQ9LZtlzsTGoyMQTMD1Z+NkLJVp2OKMAZVlNSw
H7k8yDjDOxTJUgl5vESjy9HGWrccyvO2tASVq2gTpFa+m/6xPJJ36o3TZwc25qKj
U2CHZk1AhhAErmY4ebA6jccKyH4gN8OjOe8wZP0/sXYeuVD9Dw4ZaA5+8FZ3s26Z
BJgUtX8GdNTZu4wvMuzBhG1JpBi0cIKQJiqfw8H1dGfMpRx2ZsCo7bUahA3pE3iF
QWyQNPdf3+0O4X5GL35QdbfuUxNDxj1mHbHeYn2rHgJ2ob1DxAu+VKbWp+pJ3L/Y
krZJux5U5ZVvmESOnFkWn36pzNoT9RPA4Yqu5NxpsuUcbIAVU210x0gPTtWvXFGZ
Z7FHl1bpLYo/MQYKTiJZBzp+J9h66MK4lwHjfV+j0qI0Ik644sAYAZ/kAK5f4tYO
NL/Z21kkCSIVO4V7T0Xo/xOMpxUbpUnYvqvAly8HACKaG9iWKdW2WstWdFhIqvL1
opxeAksOQNvI9PDYg0B+HGzGP84Fg+HCtV+x8hOveBkmu5adzvYZtU+tpQQWyj1Q
huyFxiyzoPMq9nDxxxWlkCD30WeAQabzfZ+PHl5L8TgJTfNP/2tcG2FCWGI/uIeE
G9fu2bJVKuq5HM89ckswoD7qit1RMEUR/AVqbg7PveKBxl7fmmPk/s1e7OxtsgF0
6o8vWMX06uhiBOtNmIbxvtdSmz3MMfBVrLkGcr5K+O+7TFRS3mt3F4xca++Oxwbc
1WtRwsvk1VEQ53dhCz7whXuBnyw8+jZZGNfCB2kDQEKtPxIYC2Rmf/2QctYPYz1i
gQ6Mdi2H1l95h8sEuVunUgiWnUKuFC+dhDujT3EcwOeCgHvrnYaQgtdMtpvgcWjD
+Rcr8mJDkG7TkHsPUFV+7CPdZfCCH10agOxChLIbdqNmu7Qr9RsuT/TAjIjyMUes
+f0ymalt8zTaSdE53HEL474959MnsEYUN9sgthMFXhCRFBDMA8LZWPjls0d7cOot
DP5KWuIVcRB0XA07PW9ZeMm+rZO7ua7+/PjNaSkp98Khlim7T3s+AWmvnFDryvLg
cXKTMBH6+I8sINkQa9WvEf2M77y0EBj3nIgL7sqRWjQzgx2hD5/rXXTGdjf1UvbR
zwxDNjCPK8PqlT29VQ1DKLDG6aludgxG84xtcYP2LfhRs3UOVUC/uRcqny9YrDXu
lenbFVU9zVRHYQSSUznQ9X59uKeYTvFV+BMAgVXuwyxAFWy6v+0f3d9iaWdr0dwj
jfVPZGUXBX7mQEh1O5v4RTXMGXmecZBJyhOcHnUkqGOCAxaEzZNHeJ0Ki9pCgIBb
Ajv2a5OnhKPNIN5/5VDF+2wcojxJjSlvbVSA2O1Ftr8BBgGHkvR4EzzNQOzRfGVS
uiNpB6m3jx4v70rk+ojE78jOr8q60qZl3+0coLr72EHDvnNiWIU8kBOWP5g2BIBy
NSCwo3zeif9eUrDsgOWdNNjVsuSKWkoRsPVn6LUYfcesMSxwsA94mzJnA9H0Hb3t
2yjFzeZ6UEDXrt33F2ntm1sH9YgyLb1kII5dVFBY5dUHpfEGGm5jfT3Pb9bhKa0D
yBin/DBV92avgLYtsCo97uGhC7kC8jgM5pvHFzTa3v/LK/vpFMqOwnK7ZRjxdoYT
rS70Js+GZ1fBOnsmcLm3dI8ODxlkc8qxu0K4XW4aMnTn/szYUWYDHI72R7+PoeaS
rvbMbgSo6nULXnRBXB7i5v5UN2jOqZfbrjU9BtCxEPWrcYq61Os1T4CGCgF4YQN9
c6Ui5rlSxSXjEG3KzIwJqeJTQhA+ddOp+qEdQgOBR+C1vv9/Z3elpp0QHl7tCuwy
EGQweJ73i7aBk30ElIYk/hQs7Y6iX7UcsSDTdHx2hiiFHzuwBitz3nDKS0+9NdOk
fX/5FLV7CP78fRY9W8zjXzyjgOrtLLKoqRBa8wkkO0bfhDhg88HNurWxSqscgpf8
3G0d+c5zwX7LwaU4GiDtoXSdUD6w2n8pgF7OiKnXsA+k5aSUZQ+s43QwUPm6tsM/
cvHZMxss4+zHvhO46yIt/6kGLovQdJ2VSuTOIsS+ZEE1a98cboIWAwWT83JgF6nT
RvKFAEzLh6evqlzGCj46iw3HusMPc0P0qZmCdg27m7RS1ZPjUBEvnVwWFgWwS9CG
qy2yDFZYWMwPpPow0d6PWbPgshp3orpZyKi+XeWcj+8bb/Gq+xk5c+NdaIGl65nS
rsG3n8ji/haB2jKV4DbxtadYwNpGBPvetgvLVrngNxpce54aY+CxNNQHeNUl0zH3
D4v7AcSBsk+eaEmWPuCgUAEm4pGyPa9q91t8Olo9qFzL4WKFe4AkYwF8jbjEy1Av
HI0g0si15EAtB7reefP7BOoc2hjo3gpj64TbF0xp66qq9Xb8X+Hxzv70Fx30Adnf
iVyq01xILewXQ4uDQ+XO37ujRvZouvXVsboUtYMenH4jVqj6CbGHMeN3JK1aIYtQ
OgHiCta1PW1t/pIMYyeYhi/7LeYfMDD6KeogtCT8+XMO4st2MCU9MSp44C0yrRbC
+7tcNHmAVtPdfJhrbq417it82YNh9N3W+M/XXpjGw7Jty+waSCr3QkX9WOTj1l5o
XV+7p8E62ihZgCFAktqICuida2pPcSMSGl6h+if2nTjgg3/K6qnAEle4xH19cARe
LZGT28NJq2t0rz8Z7FubOfzaXoV19UNgMSMMO1wHg5uV9HLGURZoIcV+O2p17oDX
WLebvQUQI9Xvf8DDcLL3EPE+Y9gSwmiZVgsn4CDHOEAjc+nwvaYFJQiHdn0Nt/Yk
fcVnfwE25pc1x5vKj/rRnW/Ru1WIT5LXTcScKPFTlfCCXGO0+nWbLNqkqMxjZz/z
Zqni6n/Atn0cbp5S4BwW5S70nCa2MqAO9rtg/rnGzb/jOqFgYsNDF+TTTsrpg2Dz
nmOzuLm3zQ3RBdckaHgaSa/ruhfMx1YfrPpKijTSpxg2O8u1mgqCHNjZK35Wp1Vi
HvwylzlYW8CoFFKNgwBFezKFsd6RIryMm1sm4a+tSxKdHus3eK+TIZx/8mn2ACou
+sTeV0/TNoxXpsYh/e82+0GuIzrbrdxqzRPly/WJ3PAhyE8bBPsKwj6SJqiUySsQ
QysGZvhhPGGSvCff5E9rMzN/ryimW0wopfSKp46xxX3cX4bnmyNjUEzrZhvFf3Ti
9JvkGXhfXCB9Mi2aXDUoayRg3Vdk64GeXYPSv5jTDVKRqCxMFGuCGRKmLBIPEVYz
oXJ0IddM5/6vOddXHtMpka7TcBPU46h8+Fnh2AKGFF92CoHiLcpKnm5Ij0I1Whkh
j5MDUUJHSyqYRvmxftogqAIorFEB+VCkjwbRzPWbkRZpeKzTLh8LEXRpEK3mwO8D
6BthRTI8V83YM0SY2F+R8Ks2B6ilWUl1psuP5zBc71vJHwJfEMgkZV5DCcp3+M76
GlqwIbjt9dyqYxA3xRwrV3Rqk2LesD1r30rNe6aNVXSWq8cRxDxFbYVYE5/l9OUx
NUl63Pf+xilSA86+0qPDQ4Fd1rV8Bw+z6NVRQBWjsUkwQboskTwUZQNYwG70HXwg
3AMhgRV+UjZiIxK3W4fGG1jWOod59uO5j3kg2QbPECoDZ+6Z6NOhVmrQXpqXR7qT
Q4YFFmIvPuMbk3Aj4h8RxZeUtF3UswH/k3M1xhsMUfiOph5MU7AhrDKxQNln4cDL
mYt4VWNNcRimDDWHnMAbxFryyiNF1h2O4B2Rc0SeQc2XJBUlmWFPofhGvgxPGUiZ
A3AjzRBn1lbIcKKym557F2two7zYvsHIXogcb2ovEbttz1CG96gX/4qTZ+DX/fYX
X9QryTvWkqYPUutCKlA6AdrPA3kNje9w32/b+QAFWCfZs0yJtJExXLNUjKgmsZ83
Tb2KIR+ggeGtLslHN3TRDKq+6khYmfNPcT4sLl2I6LgD1ATRxS5wQfruxvP8RPIj
bdlBmglCHM4cc0046URuSOBlkLOTaoyMNJRXFWAgvzXzjKKLCXR6wbTdedBG293H
3h4bxr2gru+UEMjswYMuEq8HzKPQyEzvYui0HDQp+K85IYwvb/MBbyJipe2UMBGh
FMKPSkovCEC82dNnXAHByDL6q83a5nq4iFz/5OaDUh8/iGv95bGATnn7OxBk2S0M
XkOTOrrFj0dyXpiJ9ImOWZa64garO1x1Jvg9nrt1zOfDijI+SyxCmyBtPwNdvtAP
L2fie16v60CyZGkMNEj6JiZiAEUzvaF3XgHMJ8iLW2SefU9MSQOUBtgHORUwH+hO
9ICnfM1VP9hMoEXnc4wxovVBrdmPAoMntshYki5SWaOF1YT/PfgZRWh8spesQHQp
82ScIiUqShwupAMZ7KEli581zknGBXEHJk+auImgM256mLP4pC7IPkDiyR4f6sq4
6wh1PBUDQ5UC7t3j1LVS1vC1njW0cR3cpMWCxVBTUUbQzrzcI36/6d9mULtSxGyr
x2qYqqINTBNTE2uU2gY8q0hvIKUxyw6dmrDIcSjvaRPprqtgY8X6RWmnBzEzFi48
J4sgh+8jTYy0xy5JqB+ddJRlbusSA+ewur1MzlBGmfpV0oBSLxYxZ6TRXvBooICO
20kgz+ZVibIYERiXRNPgmeMKptzTtEHCP9uWRdM47dpao0D2y5zAghDLL0RHyhdy
B+HVR3lqPGO0IgBjGBdOBTmnUnLaEsGKxSpdpOLEiYRLcVO/exxjWmPtFjFGwrrz
fykO2WbMrtSC9nVCLuBrQH7LU9hsSJPR86ycZlmHmX6/pftEHFwnarHsw1lVRWsN
3xXAfiSg5FDg/k5uHtkr8FoY7VuON1Fa/vd4mnECCEmQygldGeeyku08WJL2UVtT
FsdgB7eHQw89jdWIwkUxC05F+WSwI56IeVqhP9jN7Vi1iyvAfAg73jsMX4m4Kz6D
se6ZRJzYx7CdkEsPlFQkiChTHW++ShPZ6lzhsw91460r07A+Y9SX09UW9vrfLOYW
WFAgMgmt7+rUsaU/O+iygqguhuH6NNS4RUKIANA4fdrEdhPC7VNVYWUGn3AJ4OZa
33zN8rp36E8gKFFBD/dLieLMMwVHl6ZW4CmxkdK3JhnpB9Whhp6mgm3RmOovpY2D
DEYNenpz8votpRQF5pRK/A3fyvx5K71YYkgCEiQH6Zk3vuAdQZC39pe9pnmohLD1
YPoE+5G9HI6BiqyGHcDRgiuOYs1PiW6w2XUDtPtVehP9oFdyvG+faCVvnJkWb4x/
bCS+5md+yZGevUONNwfkZQdndcl8d8ivmunshTjCyaSm9zOo4lkdzz4rUNcAr7bH
SAj/5jDPA4HWb7GFNiSro3bGKxdTn0WVrVa2GbU8l1rIs8a//+/+S3JMHL9IUPFL
GueQ/EngFQhbzC200hSEqEfg7zFJsCwspI8bJnJUGsLRfy36l5WR3Ex8Gq6x8wPo
`protect END_PROTECTED
