`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMtdszlCWPJRl/zNcwZX5CalcUKkgQ6PCvTSpm03WdpkyA8wWcuxVFPxY4FqoRQm
O3VsX2JyR5u8u0fjMjup0SUaudHViwMPz+VA7V0Ps9Ispog7VeVkJ9ebUCQfPz1F
1kkIGn+WXSZCk7U8H0qOaTegFimmACw4GSBEaznDj61MU+wZXzuHtr1Qe2a5ildC
NX2pMrSv7NAEc2rbjI25c/MHAPH3rarvSFEFoFI7BNUmq48XTqrh9Pv6/85osghS
Pk+mLSkzpSSfqMCI+dEBJaag1MZxFW+MqzZBAzSQjWTZJBxNWn6r2Yx65EQlGgns
elXrai1oN2q3uaWgyMpDAT5TVEu7HFMhYxugoP22N4EBglxW6IJhmI9jFDZmYRJQ
CrwxMMJgTZ93uG3tQq8vKtoCx3LORmQBMwADx2MQGbzQip5DmTByl1PgfaWk8sdC
7quYBnFzNTecAljO5zEHqxKJuqmQZQW8pubzn/a32dJQPhBLw0BFrjaE5KPI+ewi
gJLe6nyRqdDltiARV4O31N4zY9zjj2XHs1iLRRZftfn25wLW5Q3wIKWVubEGq/SE
VOVUan8Z74XkxdY2yZqYmuTn4Bqnh5v20hIQPQk6fJJp1SUGvv5gjnA5WYzVC/sV
TH3jzu6M30mbCKuMThV022lTpcGn25CmjrhP/9Uh90cwkBgcG4ExXoLyWlduPSMp
lrbgSe08XrVVp6hyO12VqQZaBok9N4bh/WPvJ9s4aIT+xqWKl4uV5Foi2OjzG6Yb
SSIhSWW7SlPojcIe/X9xm9ki6EOcPpKc13LmEvtq8RvSumlt37cOJzO+bK878czS
iTpnYGgZGsEOmdczX/QLVf6/7y895tlyUESFhVg9BCB+TW3VQSGvbKEtvB+cO9T3
mqk7iCIHrjK6/6aLqP3ED1ENCAMgzqA/jFAjxTpvcrQ8pCS9zRWFmH3gghxNYaC6
LiCFq145vqaePibN44Khb5pp3wOH5IBY2Y9yDqALI45VJtFMIQLj3Cz7gEZyFsgn
XHOeesdmUvI1SGRfY+E7wZ9swMjIrNTQUqAWxzym83jVWznLDxWRF0GdC6eenpFF
VNJZlyUYYmx/KjImeDUULWbZt0mowm0qiP3J2RB6sYJVLIypSEwi1/zQj4p7wxpG
tHZk/eeh6A1fcdf8wzl23lBpqW2GoBolXnA/J05SjzekYCtkoFg1Xc/EWuIhd0Xe
W9cyra8aQWG81RWukM+stbeuXQz6e08ZaolUGPh5TxerhCppYf2JHKszqFccr6jX
xGQ4rGTPhugihPmDvNPfceQggGfjxkUf3bFRVdfm/TFp7JGW2gK7HJuRo8dpWmdc
HC7MSmZruAy9IrK3aNK3w+Om3qgRyWyta/wfGjhDsNRWd/3/1DDB26sScSso6+Nl
RdzrTyAB9KjZDsV8WUZjUHZMjbArj2NBf16ToxhTVocRuBMIKIF/jvP8lX89JYKg
A/dfzf2FVZA5QnvjwHENtcy9dWFkicPV3thLf/mxkzw8KifYgZeqMaH9SQGLNf7h
hnvM3LEnGUt2Z320TYX1ClzDrUh8aHFm+KmZCj7LxiQeWcJ67t7nyUf0n2oeUWuz
04uOzfealJsCbuSgiBsLISvfFCF01mvH5QuxB+F7XeoUZBpy/ivohhs/PEzyL7pw
AsM9IR4ik88dmFXHj4Tyfpmit9Fu0hzIwm6uvg4fFm/9y4DlyKtBsNoGVCX6Uh8k
nS1fRYD/f7j9d7Y9Vva4qpcZKzl5appmnlvyVt1EuRcOUruGP+jqKcgEKc6Ouyhg
cfI+LnU83Q1CfH78jnylIaFh17j+iL3t3d3UhkwLx/bGITF3Kbhew7eg5G8x9Vdh
/+HCB2H+7U1NkUvlqsqvYMDCHcg+mjHcDGaAyDxmUlLTHGwbT0OIDjKXw/oxDWXA
iliziVAmWq7fixdhG3m3nQHb13SlRJIyzT63hDnikFduxl7yk6qNdoydTrmnX5Ui
ARbz4SD1T+L6KtNW4wQCd8ftthK1tuz/mRlrfXEd/W2EePZXW/KWEC4svpGPq1MZ
4atm71zH2X+YMGUyBdH0Mtv5x3v8up3Yi1+GsR5zKuBnQoG4cX3Cb/EIywTd0gON
vBoHC9zIwprmzkhOWhCqf84Iy3rQE1A41+jXq45+t8SS9ivAA3C3P2kL+6/XkDoE
ZPjYDrWZbaojOIANcdiDkfKsDDOofeCOzuMa8Nrn8wmrGFEKRt7AqA5hQN8tXkOe
d38AFMr7b/caVvABTSUYVpAl8HRLD7v2QyrKasksznqkJ3HufsxDJZT+ZyP5ZMTy
9mi+O5zDTadkNHCR9Hrr6MLAox26uTaYbZdP3OYSEJBshBKx4Vh8II/AC9WgtxD9
1MntRkRjnpCylYN3hqKPtozEN5e2YVP6j5Ht6U9rGJTd6Z/8BcepBTRhMMqeM+KP
qouH3JIKznmxJcpaWI/aJrBw+MxAm7KqWwXXKVMoi10vlzf0ikyGFrU7PbB5EJCG
I1vWZQW02e0YVzE3c5x/pPBkh0jK0+lNdtl6ukUkmo1c3z5RXvyPOmfoIh5aeWVW
sRFD2cSNfjM3fRXPLxr+yCeIN973mP/bI1WIfGygDalHehBFZ3XojE1rjUdbWxNY
dhMnxHCjfCqmfB8DjJCFTvSs4UFOaVfnHiVlyg9xhGICb2hd48jBENM3eLoxZIYc
YGtPJp++FoGLtIGe1HJ9SQJHXlgsYhW5F0ETUiwYDq9INtogz8TlgNRN5AZpZBLe
9C0Ry70QB0gmomndh7YTLVQd4fC1iepeBnUHHhhNATm3zPkrVFIKTbW5XU5m+PYr
3Y4DXk8Lz1v4oWOAAzfDG5Nhi9M0NVwS9wsWOl+8KKFmwMaQEae5D/RQVGqm8ihD
7Aj5KR/+NOHvwCf6iBUN8FIL5/JVKo8Gz6sGySn0eXC8ZHInOknJ+QdxoPbFVoSp
lWu196vuHacX9zC36Ez/o8l5J1TqfrFCWOY8QAqlFulh+cwAyCWRsOh5iIf/THIk
FC/wtuYOMAKs+yNlewDnVbWNVLXYNTHpH/2xCAQ4neDscKVPy5RR38kRPcMNdTxQ
kETiYWCKM8S4ki8/nf0K/lXq+WVZBfz9XVWa47rii49jyARL/l3eoD09kyjbZpjW
JpabLprbydkMzbgmohahtYQDJ6PxktE0XjVOkbJNsXtwjBWmFkXMcvMk9EEKgNpk
8ZbWiDjgTJKjnH460LUjiIhV7gbE5F1XE5QiUbhzARY6IdPgQ+977HhyH8UgaGlj
TPthHQS3+KgdaM6/Ejx4gJXSVZ2mclMijV7iwt6S3No/4ERJHwGbOCh3lxrTOLv7
j6vD2u0Dfxrl7jguxIcaV0n5fAww+eYYo6X7nAqIlt1q5pXvDP89b3OibuX5XtxT
vIXEro+8Yajp3HchJEIuGc1HjkXfNooFe84FctyypjxYyh3Drwac9OSYdGRTyCIf
+gZWhtjDLl0zoNhJpDG37ed2Xskm9w/uDq6xICNEC3cCm2D/nIknhqsDvqfcx2+9
B564VCy1iivRtsu/PCydLFoMA96NTVYuNOEGz1tmeIhzLzkPxlFvlPDYaSEGn1CP
97SXmYPIt3vsx6Ef3FfK9GiF84dAT4IgX5JPez2KdESt3eqBhed//8W2ec8y5pqY
3aUQwOaiTW7aTu0YJYlkI4Xr07xROUrEMy8r+g03/M/c1wdcrKzCQPcU35bx+lzr
b5Ki5ixvWUslUxFNPhO6dVr7klj7MlwrKpnLFiCzMvTaamW8y5p21uFoQta6rm0h
dDu5gIPHoiQda0mEPF78I8CDId6iZqIk22Qw4fLUF5Hj6sxcRDsIBRWtteyQ8opt
CUvjL1YMOwkEmVJrlou0zhasiHYn7VNowxnyNgZ+jFgcpacaIfyh3JjoVWVZ/LwD
t4ouFdS3JNgMjM5oDtr4IJPm48EK9QocDIAQ3ZLrdagkGtSL+XO6ZLMlGtMAbdcT
7U3F+2AXyRKJUa+fpbDpewVqPWoHAfIQu5E1rVxGGYVfn7FYPXrsUnvmbL0+T+Z0
UTSV/JreZ3Q0HKJ7Q3kt8FFHt/JU9m3IkvkB7s5HMIoPs/I9oeqZSVd9wDkdF5/X
Ffjh0+fbXZm3fExgqSdoZ38Xr5XbitlrlG2sS0DgWW0JbM8mIUZklnG9Y4n3tRL0
pKMTIH2uRj5HhR4Tv50tTGFRRlkxOWYrVRErn0srLcdUkBFmCbMmxeeUiFeEEwhO
+9c0JCh/1z2VEl1tG5fq1OWFE2ttqgSPp0m0tBJosHbju6QGCC0r/hZ4b8vWMMHT
FHKx6id46ROUX5ZZ2/b5i8FR7JVIWXUzVIW/+vvF4Ia/5rDLGAzcQwyfbozWh19q
11WOSsrrXhkaAtjjOsl8Xm/2e2rLcPzcKyjozLIOEswVdalLIKs20hh/90avsztx
IwkXJTP/73CfGaUTRnr9p+53aAFeMuebtid3i6T+752TsjxOvE1Mj1v4yiIz9a+A
JEEMpNNPBEw2nU1uZZ0IwF9niu78/hSYeSVumoLC29XfrFKyRlqrkwvJxBGkKmz3
mdOy9tyqU2eWDV2I8lsnSLV8PYQhVsZMTS1Tra1yxLGN1UN4z9Dm0KJAEMn2faPp
A9iiW8YgUV9Ajmec+s0cFDUaMojzJhnFSK/icSLb51PgrfST9WiFFA1u59ledUWm
bi9jSVSvo2AIZU06p1Ol6dguzRZHlAhyXA16jGNgz5ayjHMLfboeu+OGZz8G8oT6
ufYleaz31XRjaHEasFifkUwb5YLKdubmh3dZflUvGdgZvyl5/cGfz/wMtiu1Elj0
crIFzSnL3LBdDkvgmdddo63eO9mNv2LbrX1gIZnRUpifDzWJooKPbGssA3yvCd50
nJvYpfmy3ZIH4ktL0/3uidrQCcdXc2ZtoQYijqw3Fsp6nLcoK4aGgRiMmBrl45fC
cRdC1RPyRj2uKK1fh+hp+EfpQ918WZmKN9sUWlwtUZw0uIouAsHkOiV36g1ENGjY
Ye66y9rdbUXSUdqpWiA8QjS7cwHqe6IOONy6zapl3lKftuIZjNKUEiYHfJ0Fr0G1
GTbb8WlSn4IugokUg27iy+VqaFHkcFP+oLIRpfYP6TIxiz/E4lhU0QPkzrU7e2fn
57WxRVePLywAQoJ6wLa/dF9BQLCkUOO9GrvdAkyX0TJY0am54fU/y7IEsou2zPyy
Z2cHI4PCoY38/xpShqpRHjddIBjIfg+K16NqiMsPCXDIv1dHim4csEoV6B2eiqM1
kbDs/SCdSE6VpaOQmhnjuiQfDRae/K42HtEp5h6GYMD/ZX8F/eOjwWECY9FVPBVL
AjAI0rDJdWRfoN9KfK92TV3VyhdAVmWDYveGwobJE/Tx/fnoug0qS2t/7hWRQbI9
Cx9FAG3SnaCYL3BrryGyByXeWv6elq9yv56pRW91JJN/dSTTeiK9ZuAeiYOJInzf
XImit9Ir0EtcavByGoVePQeDiIWE36tQHUuccNSK29MoqriKSEWKtiZkvNrtbzzg
39rwmrFQFBpb/eitMzfkFur9lFnjYYJV3FTQqnnnbtTmvc7B2YPrBS5iuQsm8thd
ne2SC64OYP8q/vwTTH/CogTi2+WVwSjQBpsXjFymKgvmiaVB2mGgFXMAnQHdnzLX
AadvfT+TMd1ZqXi6V3SoG/1irCCQ56RZR51e+ZPBOZ2K20W1nYZMxpRDbLJFJ97g
0cAb7S8wENAt4OB9oBxP50CP5k5W0BlyxUsgQ2nVAcRk1aeiLW6d5bCFrIDlPfyg
OWOTIIKB6Eats7UlpeuxV9MOyPIYClbZ8Eyde1yoPJthaNHGucWsQqSPtc18gCYH
fdQ4yZFAXuG7ae47Qa0TeL2HUN2tguLbwybOlQ1Pomw3Id/6KIjJ2DhnsOYgdqID
AMTn8cOy20nvJO84A4udlhtwamnQfoG4g3rt5aLPJ8+XsKMGdlTEkADOEcH3PbEH
FH1c56rZYJE0NuCoCJfOzbGA2Nc2wr2PN1Ho1nvpP0TgGoz9KGLd51sa+cZoE+ji
sJ1EHo1i2WsCUEBzBkG2yOtZ2B/7uzepk7QpRgNIdiPEE0myqpl876PlM6y6psdd
otBQbIpBQCzc3x1poI2vS/286lZX5eBKX5IPxtiRhC6oaRvjwAwjRmCg1LtMPzJx
g16diPURMvakZjsOI0jfvRhURmxpLui/6lK5WzJNbbxqABN2LDh3Oc2jBZNlEqvM
w8F3Q4WbvRrVhqEnRtIOekJTEx1PtJaQ+l4XIsPSQJkCB3A9NayUGL5RQba5a+nj
jauQcWcoyTWwKhL1p5tqjOyhmMMmS6HmkmJ0pCtEOsTvYNscR8PM2snyKNKDIt0B
JCWeooI3ouRTTr2nTrVEDK+80ik595aTrD757/cz6B/HJ018sS74baVQ/7auxlvK
aAlBnO9ILMUOIQBSaYKvAE/xICVt/4lSFZTWRbZeATbbmaM8pqesH+Q6CvR+iabE
8N59evNwS2GcKJSgYxs7Xp5kXyuRYRWhxiu4MIwTh+S6F65XnzH6MlH+wSymnaKN
DZ9Boaf80ZTKTTLTzZUzt05rIATheQaI92QevkGXhMOY9xJy/zYdkQkdK3vh2c4f
WqWDSgdO1wNAqaMa6oVALbXEIUcn1a8eWOYSoKaouWjF65OIEACQm3wtI4/XX73a
y9ItUTRQNh6xg8BPWTevO1abibx5lok4S0iOHDpspEy+YqOOUFvHvn2yPoBmh69T
7bwPNkUimGwk9GBfccIL36Uwsn/m1EjPzDK/RsbziLwzednI+vxo3cbggdMy7KrV
LGoAtY9tknmtjcjoDYH69CH8JCCUsWn/5Zo4qqMjqP4xJD1ha4+zR3vvalJ+EjoS
FXdXQocJ2rDQkiQrHRaa2TF7FINvb6iAHts8yQJPD0Cwr2qfu+xAW1R6a+z1AsKN
GcijzDV6qHHbK+OBQBevaQbBONUWDNaym29Z7muTKq2k3vvUhu2KTNxV5E1E7zlt
Kvw0TpBWBF5xDlC4fZfdpAL912siKWzr2QEoCgomQ2dq9Dt6aRw6H5UGvlIJvo/g
W8bH0z1SnL7yTypmIOHtKy3l/NOC/TsZ4mNc15yHdUaCMn27ntlQs66wQE/9dqlE
KAs0Wp/xONVBi44qRItQkR0vuoq+BLpm6wcGwzlpZziobmukaZLSc8w3/GKfnfXs
4DtErT81y61lbV2xRBjiNVKylD4DtrR25ihz43g4HU5kokSzhBnFIgJt7h59ItKe
s3PFgmrD2pfvDlGmT+Izydw0+EqqfKoQTq8p7YsNBGR/jXFE3uU5OokjH/HWddGR
5Y0ZY2Yp2tDmz0kXaaRqnLq2kxNvDaKRDzldxLmSDlehKAtUVQW4niQ5GLP7YjCz
0V2nXc933CST139l76znNmJyXTo3DOr/rsrrLoUTLMW1ssT4yGVVPOmdShZAEZBI
9AKEn3kpfGgA6E6LiEfOO14eMhX4iHd7INJflGNGUvVFVHsd2MIOg1OsSKnmtHnj
QYhEwSC3gussSR42Xn6Ysk6SUHHl2z9HNnOKfgtlgxQ6pGrSJFfay5zK75nP82i9
wzv78KPA046kZWzqSWRgikpXE2lyAb/eNeSGdpJIbAhBo2UkzWMde3qfa6Bk2ecj
wRfzEick92grT6fRRZ3XxDESrpjqxwPWgYoJQxsQ4NDHh7Bvx/+Tkjn8tTvuBitA
3QAaNpfaqyvn0NLH4D4V1l06GwZ2rxcXVtbJTgETlDkepY7LpGO+UqRht9C/7F7l
RpvPNz8G4P4wHElh8SLp8SVc9t2uOoaEgBbUAcP49qSxg7GbGLnPJV2z+P11XmjD
XtedD+AA/Hj2OwgAtvUlmTcXGEQoYF3UodiTweg+BGRhvJ+rhAdQcshlwsC7soQW
13jBHcP/tzCwf6K4TjoyGGAsh5oeTGxOXhLnHvs88YIHG/8WjdtTMifvs6etNI5J
l2OTgw66InOB2d2m9t4LYVTZs2IxSHcfV9Q3cRVuXoHgxaTHTfL4CH8+kNdgogaA
0Qwp1nYq9f4pXBwn7HgK+f/1U1FGygTWfnH8S3CR6gDXi3W1pnOalsmwOIKgCbmU
/3xDNOIJY10gtE4OkoRW293i2HoG9zDh96p+DTlHIEg2K0sPP27JAkt4S3qx1Whp
sWZQUTZvIHOmFMjoc8ljbbyhVRoovBMawTdmulMrWzevMent4qvCKWxI7APqaZZ1
PHm5WYa6sQU02PDVBSktXEF/IzcsAbLiAXqPjm0RF8aZUAukwANXBVMyILAuFer0
VnFAqWuWhetL7teTNoib3/BwccChIEutXQL1NLHvkknd5BLWmNJOjaD9UHHKAaJ+
DXAqzxehLW5njy3AEIetcoR2XtkcEk+sYwxE2o+6MOKfpRt2X8e9z8+U4Fec3JxV
Xbsh0URVEcfjj12bpZC/G/OgxAvNRs+vaGtVQ1b841mRDJjFcdAhlCVXQUKk1I2O
kVmDtgnQszoQX+zbG2st/AFCUeA8wRf9A0y9NzqjnfiYKBwuvI1Cs1UJZc/vXPc1
pAYoPtWaNU2KMICU4eo/8FAvTULc/5aMf/+soxvv+BNwLf2phM8uYZGh8o0PddG0
HEW/oP7LjhyrurGeBAxg2EU/6WYwUzyQauKeOhiLW7fcx7114kdvhkSBhnii0RIk
OGHDchhONRaNRobZyNTKuL7TgmSO328Gx0/2uNQEREp0beuilnpEMVg85Nxgo+mP
q0EyfzcXnuRh34KdkXC1FpD7JC5tZuVHK3VqFnGyJrPffol/IUiKhPU+iviOzkJk
jjrcUfTlIxst04gUxFadmpB5Cn/HGOSl0EMTbHMoIzWP6JyLruFL//VbaSTODoUO
2PEoccVXh9sKmr3owGs5EgQQtFzyDt0UcOtnsw8K/une537sLUojgeZJMPtBiJPH
LIHfBUkDxc5mT437c/RbdEoAU2fXy+zCHkuIt8OmZcndDHh+3bg/FY1tR5aS4O1j
BcGzKynIKebWPJYAyQb316tMJHOo9eB3NaAHnAkOB5SyoMlGrQrheaQKp/BwxqD0
nqTeMgKFJmqnx3ucM6ipSGKVDExxCUD3yN12tzgKegY4AyoijThL1pS6O7xawIaZ
Eb68PQQ3IUg9bjWXcPsz9olP6nkOENrxosPsv/4noRFVJogeYErWyDGPVz67fR7/
dGrgvmmh8TM3v41UP6G4AV8L4Q4+7Flr9diVR3+6NEfeKbTUiI06+7Xk+dWI4hVM
JugdCpo9/5L9RYfNPn+h6LiC6oWRPtPUKscvJxgd+EeYQu2XfEdmlZVsOqUA9m7e
kAEeZ8sCmoApGVcAJuptgp1vdWdc158c948N4jWqGLTP8xxNuUeDIm2yRyH7bumn
YPsKq4tFvinCo503ItssTLvWQ4c5ziTQ3+12oVCqSyoH9/SuJtvCrU4DQAjB40dR
bVgB8m4S2BHZ9js4ejE1eCBRBXMqMhlYLzU7+HBO7t1du+CNIKN2kab7IIoFbE7O
mXFjNG8oiPe9E/RGwdVGc5qxBqYfkm6HEEHg20JQe78+ufrJlni/WQvVSF83BrO5
0zDpdR582/RawOuj49QaUZJV9sMgxiPCW97ohMLd/MCLZL5dFZwg9jadEtytK4gu
HqMvATTHlOKZrbCva9hBXGbX8OEq/HOY7OKhexSZs7nv7pFOuCMaHtq36kFGsuPm
7GKysW9eq+RjenWWDtRaPyIhsfC6etWDbnW0dEbUg8/fjQOuX/hFu+JXN0gWsYqZ
YJc1wIukqVISAWEvKCJ4Qm8uujstQGmO5+1UzEpw4k3TawwaYrKPmjU7HkLAfM4a
8pRClHpmaVJrHaytqA0bgA3WsMANVJMy+65r+M8XZdHp9JKh2TJW7JvWMra3RS4x
23ZibrLCxn10IzVcSryqJc4uOMjPitnwYb5UZM0tG2suOED+CWokLNqXMJEyiNL3
b3mBb2TNEibYeTsFlWKaIVRCNZkLXiPC9ZQtBED0ZXEitCvm6VD+cQvPNBW9YYQq
hmh/FkiDlKMhhjrCCbjh0iITTWfPNJjEEshF4NPxat24k0zDd1VUtvLDxj4zNxLS
k/Ww8Ut4DW4ie5Zcr22ym5ssOU4EkouReqa6SEffoAtWmINwql6lulVfteMAx7He
kSJ7WIQs5VHkXVRXnMJvASgATcVZumcbFmW5luvuNPp3LEE9E41WC4KyvISeOs3R
Hcw12v4xArYrSfQ5EFanslREsQTIw1HHpEvPjc15GgW3iHnRVf3GNfAi30mv5eyk
sG6AbZ/1pOgfTEDVQoBrjStaud0rEDUOCIrkMWi+Jf5k+0UWtM2NtD7Hm8Lq+9/+
iSnntjRnSjfc69eDZT9SVW06R0CHGFCMQdm4iefIepzpAbS6DO00l3B9AoSs+tU4
epoBPAPPnwQGZnKFeXmorOqLkSOCs4lQsKmS4+GK5x88mTpcRiVavh5hLig6698J
7Seq86y1k4qA6AMxQ2ZDCnqtgTjjZ7jubVwmpArgm0S5cd+ZkT1gf07+afwGfF3T
5cBHVuAMXr4RLaKYYVHgiZQhSN7Ac4YBSyvXRs3RiGUQ6AxK1rmk74pkieaM3J4k
yodAVLS4OOOFXqJRFvbUM83bO/28fng7rSsn4ZYHzQIF/0YQCUh8Qk6MewUGsRdE
CPDjzyCCK6Ou8SBrPi1JuGR8UW7GUVNn1sJWnvb2ORknsjzJijb5OwtRePw/Tk0x
P1+b9WGJVi5+dqj7K1Ad9ncCc41//5AeDuESifRMitzPgB11CXiBNAnz4P6LhVFD
nVvM0cwVsyODF6L2+158vy3BYaJLo1JYn/WR1mLxhOnnEJw7vEHZtPpvYDfva7IF
//96apOY+Oiwz3fX7+WPXAhhEcvz1OCAxWnFIurzc7TH9S318mwMHqb1yEJBB1PZ
2HljkSlvhgdnjBI9p4DqG5mPUrctDITRB8f1aABWBFuIpHxVq96u4wvSndARbPNY
WAYGPYc1esqoUeCl9GGs4/U0I1Ynn0P3+2s+Py1bEHXkEiks9c0wEIgk9D4TQ2PV
pbuo6d1TYQxth0gtrXVtez0/QbPWblbFIBwfIODXCGCvFrwp7kvB2MvjO/PTcLth
2e4tuV4XUv5JSMf/hQjg/3hcQ7kKfujND/kdANh6kfILP7+B5Gqg8nWiK2xmnS96
pkV+rgCLvW855oK4PiWO+IqkbwF22b2hOzRRi2h6lp6UGR9vWF7uRljbeCgOPPMA
C5UZmm3Y9GOqeZy1L+abt45VaMhWKgRYiIT1308kc9Z5dGJRJcO4M9WHaux4W+ER
ls370CmAPUWgRe+SEqohjhlnjOk24LPgPMPImoX2UQUBri92xkIb6kbt3gzC0M+L
vqHUUd5SPdrlvfKveptl3FsOIMITxNqpoC9lxCkh/u+0RIZGpFmVM1Qnrr3aneFw
o+a1QQGtepJsJn2Ao6s4KVy33tDMcNUockoSzb+rhC8KsXXsw4oaDz2Xh9z+CExm
D0wgMLJ5YCNPtadZgQh6b2jwW8hQNCSScDwGXr/VZl5jsv8RM1aWXBdKAVvzamGi
2a4cBIwk9uTXZaedgsNdKIP4BZCnaXARikKTOAqvZZkZDbAVXHbS1yQ59MsMdNFJ
fHlXjIIF/oQ4NDKo7i5TzXwje7mUfHEYVlA54cv91XLl4k9lgmpsEKrHxfWhUhDc
kstMxaO9uNXmlCblzxYvv90K52sOYJDOVMkjNZan89rKoDNB9veywGmn+z9Mjalf
ILgoteR8tas8z73wSz1kpFDTEAbznUq2ipsJekUNoYcrKdblSOH1KknbJQ5SPtmF
qOUgx8PNcoKn1QpoJvfWQmN93kncYTzvpq/frr7WiVgJxWv8RzazebQWxJHhdzIj
LINnIC+8IZCzdGkpDxycez8b1dvhfZVdSLVZIOyysTxcT2T/OrNGk/HYRKmmPmfN
5/jfdBdl2Dk6LGjgjtZTPo7LTwaIjAguMc9an8rCkWrv9Q2lW6IaLtTMLFhpKRE4
hcN9khcn2Wlt0KjeCPmWuvkdasfKg8MPkeY5nIa3TGl4ztb8HV5R1DNUn02jMpWh
2Cv5a+BLnK/ZHiUSycynqt/0/hVXtRsd0C3U7u7UAmtyDm4LniFGROuQujefJnY6
Zm8uiKR73mP4udmeldxru0DNavMIohFnJZdhXnyBoNPM6eW1xCu17K7o8pxQjYPl
XE50H1xVvvmqdQxCsBZvPY0A1h6tUDBic7DDqUphTY9rnH6omlYklEwnFggDOFxF
Vqdhda2ukrpNT9VffUUToEx3gpR0oJocRDp5Joh+NKgpBamRZZTLphhrilNon82Z
eT71kVAon8hokuTZx239f/K6ggNCXPI2bTdCIcwJarKt6gesFRDaZtE27COxZKbf
U4QchiMOZjG2SHP1mr4m0ssxtvL5aUEOilndmvhSD3J/MYUVL8uCVoB8J884BxhN
jzZeHEdmREk4IE+Ebhf1k86BK3FIuXuBsaV7aZifsH2p/nb0F15Q9OY5JnpC0chZ
b6f2598hoF521rsH1yUveJTuBP2c9n0f4FZA8f23aqRpXixSHutjbuXFVhabaFCj
dJqFZJPqXMksY3ExM8aQ/S2lxhvQxEcbI57P9Kd/QJA9/CzCnOyiqIpyzEPRPKFk
AuLRfqiKDJaUGzxh9t55zLNIpsUFEid29/HA2tYmD3YsQdoDCnxxbbHZZ7IQbiVH
xJxQn1SpdbHnt8pkNxl7TUOgsG4ZBGWnYVVO+RpYITPR++X0iwArHXNzJXmVqViZ
Fie90VPTm1ogQm858EsxCKiDZ+OSSlh4cMorEIb9TW8TTvTx4Q1sk/Bx6IKaHimi
n30zqT358sFWWvPiBUVmqJT/qARGZGCVBEc5X7VDKvCrLrcKkx2NQ1ACr8R6Typ1
J02C0PZPVaYVrOI8jJ2UMhO//ieWBb3DGVIRFhLD0rf9tuEpg8JLlwQq0LxMkY5k
g34dv7Rd1N8Mg9tDMVHSo3AnOEDmKdK6xyIag3ww61/QiMoKZOsJizf9Dh9+hFod
nGVFPYImanrv4EZ4/bpDC2xC2Q6JEvahS6fTc9VwqZw5IQiTPKRrmnEOWuXwV9mF
mG+yJ7oax8cFMyxFIhvtTRWfoHwEN8bdYxHXa/EepfH+xOhyzhnnlyABGv9P9vCm
erkIG/YpnxEMecYISSFyDKHDtK+0UDfO+aRcR8Zz0HcBzSi85tHkRuH5qkr24UUj
jR6cZJYdRwNbI35Tw1UmtQwqYLt++dq71U0Klj9AC/PacJKI4ssfmP6k6eSj8+Lh
61nYPeZ1ryFOG7w/eVMImzsqfB/qgiclS5c5GSP6m49PFkScsRiAHdsjtgpq5gkL
uTAvyWwXFs6nB6A+i53s2UWk92Zrgvtzo5fl1xUcLUBioZMOycMI20YFjwawg3Co
lRJom+55MI7GU03rm2mftToymlKtqLykYtaVFtEcBwgiHWj4f1Cg68W+yBRUQScw
vhz8TwPmRLTnDKjXLPKyE1qubZlG75S39KJtLIU4C0E1bQJdQ7Y1MsSe5R7EJXXS
vnJ3UihNN/Tum9is82IsT5jIEZsJNX1E5j8c7jhwv6En5SqBdlIZIx+qvO9gHbUM
TtvdKx2WfrCqdVBeFkIJZ+LvdVfOAdKgv3zThXKvpCdwBzJ4ihmiZ3iKA71MmH8n
1vctsfvddJLfyU9JhAQW0muBZZX2DOCO0g2MLeLiRU8+nyaKWXDRPhoVorrmLvMM
WKC6rLWnBtmhpA4E8QxX5Osv9uvdzpozHnCM5f6WeqYSbXkyIxi7Fj9VfWicvxNL
zhZJQKzJv0KmF0SUKfmWA9QaIweUEO8fJ+bvCPGismsgFZI8o6gVCW82CZeF9NFb
3f/Q96/GW0n85BSM5g4hdMzcpkgaF6vyCrSxiJA1ahAmMxWMnDb2vYFhWnfBv13o
Ou86l7vZ2XDV3ILofCaVEd8NgJvI6f90Tqs+AJPJe67CKuV/y7UOMZb2bErIucNn
MnqsWH8dylq6V0XJbWmqZlDaug6jWJ5LybwIhu4kvjrREkfck+UawWyFngx3FNtF
UWrYmwQRb/oNUYgw7AmvC9Hn9jbUlHIdhlsKAzmxVbHJdTgaejiUNOfMGh1/bGY/
WrrKUZht/+rI78OnGNoII8R8HL49QD+sj9eE4kwXDbQiwb2+8hvM6vxuLpypDeoW
WyJRiReb7JFlSjWLtqJ2ZhhjmnQvZ/gawCERwmsrToXkyLpI9XxRf4o0EoLMFsAF
1foBp1F/KakZA1+tskQJjx8s0DwW9gDynxtAn7S5JDcsfa5nvto3dLijbbJHUN+C
eWq9PJcxr3d5hai+iEVQ89Wi+RYGANYDQrq+6t5g8cWtOeAEpT6w1AM0QAcbQGfR
MTRfHfF5QRbhicExbB7CBYWegiYGpEyyUAqp5BrnU2Lmyzw2obcl6zZa1o6vT1EQ
HmVGjexxP1Umj5gfFsAAIGBzjY9Q8WrH5FilZBImV7VtYPchik1rCacW5pD4qsjF
C76thdmIQO1kod2LuzFJ4KCQzU8vzyL7y89SEKrXFcXQt5gGo6JM5W86O29mlxQb
03+/3iPbKGMXGXExvjCSTrpTGckZEAitG7ElEwk1rJnLJxFJelAAebvnHXDT4vti
CNCWccSBaSHz+H2e038Z8zfIYsLbvN8KfkoQYUXb6uNh/uFNTUAER6x5DcBzUZQj
UV7fdhlxnW+YR9S15N5/9yfWBI8S04fQgromBxkYQjYE2lsUMa0GHRC/BKFFPvm9
t66e3pQp+ZFspwFrmk8vTC1hS+BdLjnXd7JqRjhk34TNgQPYNnPDQkr3XJ1x7jC+
czp4ktma8t1NDLWE8xdU8BIgkXoWgrtEjc8uyN87Fa8okvtWAudR5S6DFJFP35xC
qi0vu9R2IkJYTBbAphuiC6kgjoSrCM3zFzjNV+iOLH59GIlieUNJulYfGzGe9Ey0
1w6DcJBUyteZN82d20305NPzvHVNhok60UN43bVnfZ0iSTFGtMhky9DiqHnDiZK9
Z5OWdaMe84sNU+S5IGmGmFlOIbUQXY8RXdfWDDkabLqzXKgWTCPRuL/2c+5h6BL0
FKnxZc/uvP19HQK24V6C1MmbwG5IipHlpOEh5lfuYRiPncptVpd9m7HfnBC08Yf0
zLQz7gzS9V3Lw7Nzcmwu/nqpKprK6vXHSsIjl0AhImbQ54sFbksAvaTO4mXYADuj
HRMdEGYfdptPrb8ePOPPOqzwKAa3Vp6pDevb4xEj4Kh0gG0ZZ6w+OwL1FUhghLyX
RGjb2HTXLxqXLQRM4/GAd7NzZ1TrBwFT9G6A2aTe2GYGqMUMf+sOz0bcLO4VmqxJ
VhZdhMpBndeUInHjzgSmYY3VbjUX87Xwzue9qADLyBDCi+DQvzt590kdErLKz54n
/NwySU2NH1cx0Zt1ayVi8eHKLvjvQods60cnANl9cXIjSxqTx+8hRqCru32FLZBw
KIWcbwPPdn0rkDTSFgOaOyrhC+bGb58ATQHSU9Hw2W9k2xvR+jIdR4vUu73TGxiw
Fij/93IfmWxahPBt16xkEK5KZIOvGJ2CNldS5roR86e1CIPUUZDw37CRErFSTtC+
9JH5EDOfbO/FheBRmwoxW8weJWCfiSKiL19mHap3baxjsu9DXLV9I7gRqnkkDipk
gzOdHgkJr8mDqpxqwInjZb+i9SiVMpFuBVtM29ij39Km7kRarcuSIjYmc9CPKPtx
i/lMwmGkyh53qu1bPaXaA99FL9bTl3PFX1Q6zl/28Hp9lqyJmV8FPm/Ps2ywaoc4
XxOCwb17SV/a0mSjRLF/VbOyOzh+XhP0bqGNCPcptcAnkhPesEbQdKb8Eeih3Ozu
qy6+g1s643CZwtMkZ2xMulZrRnAilOd4Iuzw15Da44l3CS/GOdjjFirQ3hWzt+pK
7+RFPPkcO5Wnxx8QCDb41VlqSfhYlUAXDng3ZHVPa08/Y/K2tFtLth7G/U7nuxOg
y/9Mas7NNAG1Sj8ZnHhJxp3I6bPbUtTfQKSYdnD3hUuEEHhevr9inbDKtfVdWvMM
5aHWKy9JNMQ97uZMFFCMzDtR4HPKOmtf/eUAmGvbeach7xYqvKygoV2dunql0rAR
jahkNc/7PTd66x2JYm6dPXLw9BMXkTt6Wm31shCRDXsVyjoYENtaOakjgVbDUJsn
AavjX7jp0av5noOI7gbwK0vcJzW6QuxeNX88Jl83DpIrvTVuxmWqplV6y5OpmaLK
vMArCDOGr7Ckl1EOqJdfkpvvhhUdwbXK0q/ZlezBGkeVx9ofY+TBsLR5uOlILBi/
DBmrLz2e89Hl1XpBkt+yAjT7xH4mJXBX7TsCjanCV5d+4jZS9d07nmsNh3Bmvj1C
Y9vrwMY2Cb9QHQ36OqTU77IElnFY41iM0C3OjKRSgaaAuEChThwatHxIe6N5R6Yr
NlexoUiEmJefZ3sVzKJtzfBZHnkStRLXVobTKsVfph1Aa5E1n4zQ1KAC2x5Oae6E
HWoX3Sx0eQc0+RNyYgXR6EPzH9zn+f9jP2NdOduFMCkjMoJKOC15H9zMPa7ktDZe
ju1yag1N9n+FYGE0w5Sn5U7gKrBkCh7oGh/PfF0naHXfAlmbZmsnt8e5l7aLQOej
gnd0kjg0Kv/G7eQLdpsTTWPb1+GyMF1TtxHbh5x8JEI4mNhjVwk9aLkJpJCTgSMz
I7x1j6D0G7955Gm5/XnInZwzc2WOX8oHSynH7TDSt636qkGkrQDOh7u6GX/SAJuk
FlNIILlBG2Oj2v+euW8MiUoOdpNqhmrtAo9s9jOBcyYfO7EpOCmc2hKxkYo3bbZ9
EPlvo8eoirQkfGnyqBF99zVLJz7B/PbLGScezBt2q2O14Mx+b8y6HPzNI2Q66h49
WTSKUH15ZUHxxoo2Vi7M0ckn7gB12sNh8SXMexCtME7+6qkaia67ukw6d1zuCSux
5nlx9Q60hxFVnTU7vfDOWSxsvO1AHZYSZBF63+47I1FQOwC07euf9k7lJWRxS88V
KHMWeWYJ7dsiFmag7K7PMuZh6QqBF1rFvcd7C6GJdsDSGQYH1Ei526LQjPMpoLE5
N3bmOZi/thmjzSAeYKBp8sw/NIZ5yvM+91GdLPW6Yqjs67/NvFUtwoVUhsaftwua
9vf5O2cOE4W1DIB3M9dXDqCOIsFXJSwMXOD/nQ1y7jhWxzQ59t0UQgOmP1maNCwc
W6cDQKJgVvpW6BG7rjNRflcyGjwM9Z4wcbXUadqon4oytUE493HRp8ucLb/2FKh0
S0Fir+R9IiGrsOXbpnBuFIHBWoaL694rxhnxiwk7aBAz/pHNHzvKfJ7fugY26Q5Y
4oWqpxiHXZCkgeEEAQMbMIsa1rp5laIO3LlAQA656VxpTI430bAU/D1vs5EUjmVR
lwVhfDWGi+vnf/muVTH11So3Nev3EHosUzBrTmp4762cHShjvYtr+8tmEZ9XXLo2
bClSwjeqGwzAgMeCsJiuX8bSlx8tLk0PwnetC4RwVEDlAbTCdY5rmhb1ShL6u/6g
aZ6tr3iRMxeNUSbKqH5bRSyQL7vDn3AZ8TSoeFlcRW9q0DvAl0v5rL+S9GORWBik
tfFixN29tj2A+NElFSlQHbGfKjKTSvAzfG8VK9BXxEpnuT1dS7CQaM+fp/e3PfZh
nZAUYRfo5L2sN0/v9wNhd/7XuiOtx+vbDh5XgcdCDey9ycBf2VegVpsh73VXpo9Y
VToBSZSI6kMiYDcTYtYEoaj/uVcW+kl2dOvVS6lPqiQm5dT0j2l9CFgrneRoIW5+
/vv4WImDBeu46M7LLMMZUxbzMIvjEHwpOQyerc5qy/DCz780odEs4kAuuPpo80dk
o1kH5EGuEe9z3DC1sopmwr1tmk0nYtuwkTG+ozFCWpGnqXQ08rjL52i2X/YVxPP7
kpPz57+fuy90boTt1scrkOAFfm9Jf1NvBu3bJsYFQZ5VRhQtHPdpuRwV/pib6EY7
maf2g/ediNEuHJrEjEShR/5lrbWRO3HfgY+/QXBFQWWoMrkgj9/+jq+ZHWBazKHT
xqTh0k+hyBX3aD6G7Ynlp+PjILblmf0mnGm12jLfu3YAZNwGLkrZAzG1g9knz1WZ
cbIl6hV2u/bQBCOv23erRWl06cFj8omU5tyJ9eP4FFY8IDVx2Wj91N7TFxY2qnEG
VQD39l+aV/K2MXrv5xjpKKiY9lYkvZ4ERpYHpYX2NiuNveCJx/Eoim+H9ZaTd0IO
FKy1LI869JQ65qwVwe9rUg5xxJaUVjPyjKsC4knYYFnzsteRuJl4WHmii3e5BUzo
AyobmXoIwFP74x5BuGqC2opQP8jldTAd9Udd57QvtZlVTmsBQ/GUa5Vmm3T/jYg3
3+KkD5YwV4PASpAzWpNm+bcU8/L2I09xfkolpl3RhcVB5fZw9IHWJuNGcQ0cyhAV
Wju187us0Ii/rc6YF6qGr6nweW1LdjPJH/7Op+CoDnoufIIAAXlht+8ZAz7GHPwj
FbRnsIOPNdEgQ8xfrl5j6L3+NfmOLT1B3j6YTpnTvA66nJoxS16MjLHe5240LaYu
F3EzA/dMD+u1pca0902YHNlzdHj4RdKBea2zJjdtH+V4JqIqKFJEEJA0ADMTeiwT
GpiyeWkQ7NInSgCh40/CNGxAa3Mid4BOcOlWqdkeGJa60wYQMi/bhp/jy2xL8MkZ
BvAiDuJ5oPgYskVJHRv+Q9KGPlCILXNQODsLsM8sqwcZDfrQm/czQL91s6EHPyqs
cx+kzE/AwCmZO+Ez0szHb/c+DBhQVwp6dIiTQh04SOoAVxdqcfPUBRyZ+Y775alb
8WHYUC5jLBlp8JxM4fjkI8TWu3NpIfMOb8ySNGMQCAQ4fEtwSOdrQOHbmqRBJB4S
RVkgs/8vkHpypejwctNUd3Iv/k7aApfSw3Knb77VNVdfJa9IrlYFI2OLtkfhYIPK
4DiQ188Qn1hBDY57Px5f3Pn9xY176ttyPxEGyXUmuPDYo5zjFf61w2l03eDB+54N
8rp+UsysEAMusopAK69OG+yT2a3AkMiiuWHRGpdJJQD/V7dlDyuXA0c701vvOx3d
bZS//KtaoTxuRlF07/8yuKp1bylXeJVawk3rEaYlehRw9E0W9hGEJIqz47Bem0Iy
bgY2ySAmocr32BkmdCFiQUbMAcf8thVmXPszQGBZQza6dvFz1oRV/Iz8HWO3RlaG
mqgZb9itTTaP2mYSX5YKx4m0bcZuy1lDCDyDquefAefPSWyxeZ8htzb/7RUlFkNH
YNjcNrO5FGgLeXP0Ob8Xb1azavq7zmBRNV7oZd6nzBxBisB+baYnhRK1/vnPbhx4
dGBkZmnSUDbAm2BsKtf8uXvwrMxsOxW5/xgBgIs7VJr4bZaI7HEsTzlNvYDX/sRU
eB34hJa5QUIKRh4w6w2DzNIriHxxclXShw8NlHm4t5dFVRDVFc6eP4BcCW/57jFT
ssvWsfoaDbVsIIt92cTozpb/GfOc5+bYv/BRpUcEccwB5WnumXN7cJUu3cvU92wn
cYI3J4yrKM7AWeLHKplkcbsNHK2RN3zGBL6eOiZk4Aze6PmVWknJ68FcIsQR4+Kh
fQEWYQgN/m1vuC1vseIUqJxEtS417JYWiYgFPj7MZGs7jzhniyTBVTjfEHhzBN9N
LupMK0f3wcakCB2cZ/zfflB36JwudJ9DCN1dzcKUsfsah0G7K5l/aE+kDWtNwsNc
0LRNT4dDUDXaG34HJpcv9JBUYUXuCLtIxRnKz0lxQTy4i7U3ZcO7HNAPT4mTTJca
8FYZbYQvAYJv60FBMaNWvdQU68s7FhXqtTj9sEiJwTUAfhDmuigzu7pqkLycTlzb
DMPfx0pvnb8j4UxMSpTSniS/Y7K1r22YIl5vxsrxWWdOmqxqyicExWyE8bdH49UV
u8BmI84LqDvs0zHdnMQsYGYb5mIWrqPVqUkt+lpm+AhxU4oywo6VQSxZkrYjiBPP
qUPre/0DuFLlJmtBxjOyOvNqQ50gG/MnoeeI8d+S3OOmJUYgL15DqYWGCW4XGHSD
D7pWStL0SezkPPMlPx5s23BrpZxNXRYx4nTsTxCP7T84c0qzNkXOPEh3+oZ9WRgn
gvMf+OEDJeBLgjzmrR3GA8dx+zViKzaLZ+/OoygwXAGHkgedc3TAyeEcupDKoDIh
Ze4D/aAohKezFyzJuR2cMTMyp4/Bz1JtL42PDhIj3CAYYaLHQSBbj0lvrcbuqEYV
M/EmVAxIF0+8JgWPYa1Ad5ipsxvBvVyroYhTjdJ2/HBvGJjj7XQfJnfPrHYyWdda
fBz5t3hBkDi44veuWkw9w502GnWDau9t5Zn0UUZHozr08Q05jZhIxJBTFOxQWVL5
Q0BhIwCLwWkTKkLnQbNb6XypfOWSWt4rt3HdfkkXfx6RfhOTFRrrKv9WzjSvbk09
jBRu38pl5prZGycmcrFkn+q50/i07h3F2gy35INxQwzot/iJFyqJN5tEHl0Cwtxv
gKbeIWPeFeZ9q/ddb89fq0T0jvwtcVPY2tTToPiHMtXlJ8TQBwRnDIQ+BSKJhSWU
EUvLuGR8JfPvY+sJayXi1VtmC9SRUZ2kReiM6t5We/v5dw8OVhmriEHKzYNsLFmV
enyJdDhpvXC4bI7xioCPcA5gSMXrabURg5iru7uCacEaWocFhzphZru2tsCLQK2v
26dOaJLtSVumaR5lRgckVJvo82A0PeQztgSL0uflM5ZVsS85uBHBp4LWUzteaRf7
AvVzBMbgCG34ziPEvLfrpVmZMN6ghp2+afixjXh5hEtxg9Ey2qaUK1AvLTxtDMYb
eNgc5xRssm54kgvu4CI89VPqzbhZy89XKyEGIMFc6LpE8wvFWNJaZobOn5ebtB68
0vsyRSeTavnKRTxaoInHZ2I1dCiWbbQRunhjaenY5bNJrg9epQgtHdSupZWD7Mvf
dzBHi9s6xa4UoeVQjb9ddY7XDrLoxreOX8QMFZIuUVIDmsbRGsBHbv99Vrcr8T2Q
Rj8x8Wny7e8RZQhdA/G7osPUyQ2XG/wL/VnNAU0XzryuX2CV/KtSrY279TdjxDWo
V+Gt17zpD1OVqhTPR0OmUmqc32AImZARv2jdJPjJ438agxrmKnilQLHS5cgon+nu
UDQCbf6sf3dj45NbvfeS6AiQ2ymB7qd8zrAWefKxx8g5Eu50zk9P7rppURlB/wFK
IIbtwDpxswB6miEbg0rQWYC+xhPQ68sxHHmMzwCPEDpq+zjxr5MXQKVJOXGkvlVg
ojRGD11/v1KLGYO5nSAnlyTYM3IbO0KOHKSKftwrRK7YE82sG0wCB1bfH6U/Zgea
oQugegbJG4dJ+n6RvPhl1lprAy8JjQr7+FBicSPpu9t/Wu5eYWzRKoV96MP1oGW/
8CUD6Nc9EFI53IiOvoly4Evevv1uL0L7ElxoG6AMWUHraVeXMdxl8nkyR3/WgBpY
ZQKXtgV4slQ8oLquMm/KWDO5tZ6mKJOP2FLCxCt6n8IfaWXTMvKEvanzb2ANiej6
EoHQ5StbROdSkEhREnQg/VEWyPUhII6B+cquXUf7Aczz23dsLuj9T3lRCLRvfbxn
xk4+C57RCqF7ubOT/JeQ2o+QdGQHVcs6KYyhNr/pEeizTSQycRsQZ68EQMNq4/Rt
iiqnG7YVuNhTpcawL8eiAZ5vR1CaNzc3NIKNzdKV1ZGqI/OnX4W52v38J87mtPW7
Dp2kcDIrr7hthR//i/q013R8fC7hXGKPZ+X1hUFx3M+ahixofzIKHvg3669OrMji
/2eO6ltlXetDniyWyyYGxkYdph1+laBrbWwY6bqTDxduMKzwRqxDl5arfI6YG5s0
C6105epRS6Dhn9oUSPBMwo3wiImpDCxPwx6e/9mlBg9wjWqhxwX/wdVVKFA/vY+O
JphMsTeLk9P2OV4x9HhxopppaXmIjoFsAJYDAZJmITeVJZ/5esYpdo0kq97GHrIL
Ii1PwZ8JBqKUEs1u50YxvKhEMCO9YMQTuc6nu3CIpQCdVh5DMWTHaHjYDGzZb/a9
lPKw/o3cVVx33aqkjKrDifyi99gHNuz/MkhIE8RqCea3IETSqjHJM+xtpahdlR6v
OcX8MW14T+3a4lT1g9320glVEOxhw6SlHOHUL0Ax9eHvy4nEWoSUfWP28Gy5hFA1
XRbL88Ouw1exLPWimFSnA5zJq41BQBdmTdrYcgiY5Gmr0NmVSpupYF3GUQbEWqN3
ASuiYf+0EukMw5U5C16Bv39h3SlZy16TxoftcYNC7+JaC36KcTTqiAP0cbHzvOZC
pVwzF6TmyTHzDh97I1pRmKDdY7yQj8bcfHy1XYTFrlKqEPR22USee5HskBipKQfW
zhyxXnKYlLvJWsGzWJ9kiAEvlxdDR80teDvuKmNFoTGMXKIqD7TchlVUhwElIYfV
l1MdggQdgfzFh5axKGf6n8FLoZsUChuXT9y8aOsB7tdVI+0KyBHKIfzZGVt9hppy
zJBlAZdw4kzjvsK7IA4c2yu8E3xCc2TQI/1OEi8/6ZN3mNszPrtqf/PXcHruVa4m
BhJd5R0J8r9ZWuUxex9/5QtVaR4+/OoEgnevHAgefs7s394kseG90SdUVeycXjGm
9TCy+yBVHXbaAQjlNTUdTm5nnN6f6yphwUirEffCMymxUbe0bOlhUQ+qGKZjOu5t
Sx6Vq85UlmNKUS8A44r0p6m+SCMG5uWK5taCx9Mw1ZbeBwP09SVJmrc4SzgNEytA
kMYDomksQ1Z0oRcoxkvwlrGrUHfMqXUXw2JJlYAp5yvRv++ZwCTu00f+xjA8Phzl
wmTijOGM7iXG5bK5oyw70sMC5ksiq/yhkxjJ/dGz8Ls6sJEpmJbCq4spH08wppTM
qnknH3i6gIWPLD0bf8mt0uttCEwHZyZ8bOeTATGI0GGdBEMexGUvKlOiurY0/aQ6
pWttHxpzRBBeQQYXiPj/46UzrQbh6odR8KWWhxGickCioHPxGw51JEr34sRm7goQ
OTkQjCAPGq+zSPxWigine0SVngpXyaFd3ZqIueCBf5EKGg7TM7YCwjWVREfySzJ+
W4oFeGAYmnQyxhAQlCfhImgYwG5/QAyKfreVgXicmzUVkVirs2UsUS+6O1UK0QC7
kfK3jWv3PIpJ6S+Xwt20pqOvOVmQxProsj+rV1dV9l8fSFAmZ24agfBeY8hKfckb
z+18HwF4oc2zWaUePPrpvGIE0ZZYsXqoaex0rsxnMkXFIB+2uCP/eqZ4lhoENbSV
M1jWyZl99y7dshvSt/1SNq26D7qLkSIRALMrgfBTqgxi8g09IESKbiob1hq7B0r2
pxsdO780RMfZZMmlEb9Bq3m3nhfGn//I+xl4JiefuYU5IS6jTx2PF7M0BYHOOaqB
GHTukMDMsfSuUZzi+r7WRvD4U1rDSEC9/Y/qGx/C6tM3MpUHr6kMD5zgwWgIfr0R
KazZz3JF/ZzQMl4MvLclv/lrHI+n35pEMekzxNFpW5OTOiqRE4PhsyLBsRgJvrGi
mONy/2b6RkbzjyPmGeQEnIZZT7L7fUeD/qAP4iuXS9fG0VOxlQaO2I+HiPYAPJB/
2qGdBsH/RcgmnZ3958Yn2p7mI+ElmBJBkNBLlbfWMJRjerFHJzY67rwaegGp9e6N
VNKUTYxQOmNXsXFagHw3U+Da6lQtJy+X9GUBTKnFCafOrlU01uXlyTfiC5jYZmf7
ffL5j0Zfb+RqIVHv3aUqiHyPuUETo6yROUpKfhtfDLToFl5effmBYoB0XuWzKwfo
MbO+0KrFbiaMgWIu5py7w0oVdSMCQgoGsKGJDeL5zl2jdKqLundAuzCaAMLLlrch
xWbaV+7IFplgBY9OJnJEcuMI/ISybe9MOW/x9jpG3m8xMaYrkhYnK2CYQlQg4Cnn
H0XV8P4gTaZ9HtzQzd4dSu0629T03ywivDSwuJ44PAkSgJLa1pKOvZx49ik+c9k2
RHwIJjXAl68JN0LUHgzIkDDtsuuD7wKBdE6gpYfOjOssJ2tSgYb187G7nhOjMCBF
eNcjE3itqLu5MdJs7WE5rEg+vKHMoKn2Y8FRxKpP95C7D+mG4b9HGpVWRvIRIUId
LL3ZVIg8B+EQY6uzbguw/QxD5xBF9p66NqpOT6slGaLl7usGsyk8CNE14Tk4c/Nz
hCla5M5B+FhnFJSdngIfyViI2tiSdJRmaPfm8dzLR5uKrG9LgdlxBGeEUBc6cjOO
/lxW8Uy3pT/PrIEYXYrSo8+hMRab0xO944wSMclYJ+zgSCeYEJZFijJ1XpT+JfzK
qAi3Q8hfkPQq/AuoSvebTl1tuO6rCCgaxVT7RtIEYmcUDYpnPCnNbZuDW1/6FOS7
6EJ6N0EwAxX4tCBz4NkREpZbC+nMuFyM8fKwQRLVnQnALWmF+jxd8G83MekRYdtI
vcvHvWi8UnO95ingu6K8Oz4i0c08ZWxk2fkh3HUHMWLWbKDAG2+yIHKZQesrUmM7
4kJcYCFTnOtM+vvbyk5d0mqGDS/eT+SxGjhMb8HM7od5bK2ztvjkSE8X/Hd3PTOr
0i+4ZaGlh/58r+YSHX4qJOqunzITV44bvnFHGn4Un2B41dIDKDErUTdaFalro/7A
WPKtiIq/9q+gBRxJmstv28ZYXyiNL9f3GgCnVGEf2dCBByC3rA+wx3FjC1cu6D8G
TQEnPGe5t5mM0VU8Cqst6cUhyVfNR+3ltm/5q2vpcuuHjHdqek8zDsphzvzyhyu0
/MqzUobTHNXv9vGlftIkR1QqnXbpLTWaEfgjBeq2wsl7A22mBzUQJyqQ3Gw/3ro4
6XtjbGd5DlQUZsh3obrVC7C1q/7i1e9/Lc21uK5IPy5zlf6PZvAq/7CQG5b/3heK
+hrUHfbnBK5uWtYdShwpVWnpnKNLDv7Qw3JtaW8pvVSOi+N0+JUkVvntTscYWy3E
8J+cFPfAzmHfalGoM2jZuyGt3vWjEiMMAVPwtN4xVIDRdG9izpg5pGlNuj1AvHYc
70ZKnnyruIsAjJtYyFJyZ2KjIFQAaVQUUoBjYEcTSxfC6dXeYQOgo1sH9V3yFqXR
Pocwux42KeDnS1ti81MJYC5qd9RYJ+O+HzZSAyL7OYxZ9c6+QMMgEkxMu3WLqddl
sRCuo7gRG6Ik4OTsxm0gCsSToHw2t20XfFB1ImSh6EzB2fQ1l7AsQmpyDhNG1Csz
NT4Fs2fyGXHhrV5BXoUUlLWjCEBSJPTrm790mSj/ImlIrLB760mRAcoPzTytC0sC
OCBvN1PDtxZmZpye5iSXyqOOoNAiPxnlD4i53M3AwW8lnCCfmTmtMlavLV5KjEkp
0HmFn/TmemH0PevaX4jkYTiUeQPhXmZcNu5YFcwO2Rfb/U8PfOCLpd2H0J8ZKGOL
eTux2cYAUQml1nKNYeZUVkCdyjSovr1zSD+dgxofJxmkGzxn6ckZJWWQo8OfQS9p
vAK1g/lLmQChUf3kDdACKHn/1Ga53et6jK6Tu4cfAgELXA05vXqI8V/qzQAWvI9R
2Ffa6iKqvPffq39MN1Tl3vDs9QAuftI0155f3EoxeLN2NAWI6IB7T2YFuR0JULgz
I12zsy1Odjv1Fked6KawosFN+w2qPOzt3amYDqSFT0PLJzTlxlT34fp65GgmHlTq
S3QhaD4cYAmuACjN+jV0xkDNTOvqWDLASHvHMOCgUaDx9dZD7rovnodl5nBnC7pC
38P3SLCGktbKi5xIQcP7JFZKen3gbQ1xzuAF4Qb8Qt9WuS6UTxuUbTvGN5urwvJ2
YvK3kDbsdh8SygPJI9lZqx/xnsMgCQIQ5DZraGEti3kwB3ZJsxeN2eijZ4mIP/Y0
74bNnk43BqHxXiEhK645AVNt6wKjeSAXPel3ErErtLTuiusFLJH7lWPu0+IaxSP8
wFJJX/3x5H8QNubDgbP3n3BySM2LleUlcvxBlVrotrdJGynlyufaxFSJUMwgDmnu
p9eRp3LZUzwsC1+mvR8kWIl1tnMLjl9+pQN/5l3HSk37GDZhWf0mNJy6LvE5KLjG
Sm6H7kHFJzcVLLExpPEJvf2E0t9uAYuF8SKBJDYVHVX0+gKk8jg2Zpt1hXDcZSJ/
lJOVy2XWsXEFCpm7f3RCiX9I+f4CCbhdkap3OA45Nv7bA2+ZXgAWGxny76spSGWU
5BG4MRhG45SU5SqDOlAAT9O9OwsiHcGJgbq8ktToudRdfaZeG1ysvLCfXEze4e5n
FvsPwnwQQDoDPLR5M9WCKxgQ4ifnjGWAb+yZrbQ3jG5jSx1++jJiUupBOowobVn+
9R9NkhNUdy25QBZIsFZ4jXRsh2k8pNqsNAKmwZEljslQ9wfNgJgZLbcLv5qJ3Uey
6rNGV/FDmL143Q4HB7TBMi+c16zZFwJEGxT6k+Gb+laL59n5gfGpsDrZ0kzuVSv/
4JfONEYB4hf+qrEjuCzDp3ECAXPPckJu3uR/kiObpeZRT11Xcmo6iu1IrE1aZ6UO
SGQBDsG//MHL6zZCmLLTrWbeT9kiYbjkVDsbwEA0kfoSSDwtdIF9byud/Fk6UeT2
vTWUWVmZcafEfzp5owTxEPJn6NlQr2KdcxdeDHkXKK//5kQkaEEafOFDa9pos5BI
xkqsERsBepZ74q9bNj7CIBAYlIf2rg0q5RPN8pRfOoTpK+H5wQUfhiZgurjXekzU
T5xVqh7Zj+DaYT5MvIaQaaUk+7ITb5kqA0DqynQa6xommvnfP1KFSaeM/s/D7KBh
zxfRIzQ+QgbOuDmLaBK0zaCUCH6krXi44i2vlmJ232kMz/QgJ3oJQg3F091zkCvT
KLz/BOe3inO9rFPbQaAeLE0JLBel+B6fkZs4s+Qx/FVWAT4JaVvjuL3JGdyNVQqu
poXHcOeB2Xhp3jQm/3M/EYLj0WlBo3AY0Soofl+yeFHRsHKQ0Ke1iRQaU8ooAlB6
jkOXLiAzSvMGp0oo4YFRykFf0RlxWfRhjZWahcAydEDklRzEAUzy8iU/WqX6gMjx
06WgBPBWIOuGl/YvTu4fT7VydFMVJ8FPX/moG4OjY7q8RvihWhS7p9pZwgslQ7r/
LA9NrN4GC11VEjeRrqbBzxmmbCDywJRzRf2bVYpXT+TOPisZGQzyWQJdx4GiCWZe
JjQjSOIWMvlAL2Dg7dqRiS1hTKTIZeSmkM7sKsNcYfPfHG5S4PdNbS5aU1PhwiGL
hoIoHFiAR5fnd4KRJFp+mEXkMd/vDR7WvefXE0Ob9MaPjZ/UawfUX/V9GArVGFOB
7702j212iX4dMkLXy4anQKOv/AoyE4hV0j2j/V9PJSfGONOXOXgC1E7cyzN4I0QW
Rs3wnM7M0QU0evG1IpVUBD1lvSb/hHwqSWlPZbAeFfp5VGu6gj4mpr8J0sQeKTZA
YoxVhgfXtq05R4uGUys0AlST5oqzDDcQknf4Nnzp3SBy91IQlgI/YPNtcyk3W9s+
QGMKARWN7Nb+4d4EDhV308QypIG+B8QN+bIDDenV2jDW3ybuQXU76k505iTSpM0s
oCMmmRpmnJr2SWxzneKzkzmN4OMrgQ1JV+5WDaCLRAAURvQB5T+8XnJKlYD1g9os
T2DWvIOWbkS9iHmWAEaqP0N8ZM+/gxRfu3RNlymNr+vuati7gJ4XUjKKjeTjmw2b
9ZWXKE9+NDJnpyHuB0OAorUZ/Pf7xmHgpwDqYAOQ2v++FgDflF1jmi2Hvj12DUtV
ETiyAfg7Hv3NT9J3Zg353iSwVDVJtRxEzXTcTwHsHpH6p0Ov6h4lrKOBiKJfWZj4
F44Y0okWziJGwxMWF86rRwM8E2YDTNlTS2ABtIgu9XBxsLehMgcwqLgaHSIisyWw
HqlbVDWu8mlBCOWYzkqXO7nenTnf2Qg6gBhOZ8PEQpJHviJrGa3SPOc5htOQlxog
elMMV3qbY6DcUfI+F8eugBCsazmytXLAG5j15bsd+dg/K2Mj9V1AzEzh5rkSgLrn
fEvYj1zyp+s2MZnT4hrqhReXm+kkaz1ETR7P8kBr7oNO2lqDP1l3xVaFSgyO5jBs
F2RFOBKcJ9wQXjEqFT9q76/LeRYt8gWQzm4oLmjaWM7t7kk3RrrYjkNEbA5RRAZL
6sh5PtOF22Sinqs3+MqUsvng3rkY3JQtUDbTa/hQqBEBWkGuOKmiA5H4E4abSs6N
5b6oWM9h0FjtxnPqMSyi16QGK28GZTKyurnmNkxavFHHF7E/RwvAzxrBN1kjSFto
aDGm/+d6YLTKfR467LxLOmbIjNL0l1m6ikotIFw+agGG3AWbhRxCTmKIWO1HhGos
2PZ/JTt4RwSIjFKz7D5HkzCA0LqI1MsIiLi335NdL0zyRjBvW57JWVqn/khoqfW+
pqyX4ZP+iSIHq01yIlnusIGEfkbLAFkJJJt7dixAGLdjmltST1jz1a2Pml3/+ewJ
3cAWNFVRH/mnWZ/9Cazuy1ZRm0213qWcoxv0KUYW90+gMy6imZawPWx/lacSOhDE
87iNUQgfLxAm4lMfu88mAWdrK8JAumF8oPRLHCPY2u7dMxI4FIFpT6cdR+rBRLPP
QIM2ezG8x1I6lavAMID8BnAg6Ol4PYYn50UuDB9+B952sGzdphGgPkLyeRm4023K
zQwMrVQuNcPTQ/KhQaw/q9pKscTidUhU4whRVkf+qBRVeFK5QgkajKgrtGk1QxSH
SvlRM5MYDajaxUX4VnQdvyrC7oOcuj23d8f/irzWQNFqpIdjp7tWT8uJFe6klUSa
7fVZb+ATV1D7wHjXWmnICFXGFwAHvx5Vjq8cRT8YpZVTcZ6vsZPx/dLA+UWad3Vw
MIE0kj9oeMcYRllp1zwGrH/DRKvotA+Al0WWOaoRu3xcly0q6T1Cgq2MFCTj4Py0
kFAYkuSbgEE6IABv7HkFDp6lbOeWod7vLA+a9ESjTm2atsPQRr5hJiuufc92zzgo
azg9yhdcD0ViqYkp1ITBGJK8KAFE8GFahPqRFq256P26kmZIdk9v8RNfvS0RLMeG
oyHxwEWG3iN56NeLLK7AYkTVJxia1qULp4KoDqOou7Zvdn5JYswi+rCe2lb4bh1L
gzrtc5jO+anNnf6CgrYkmdxrg/1xbhP20Vm3oGcbqxAXX3KTg0ApYdsL0qwnBcEc
xDCkSoOpR36QnaEt9238sfLxhrHztMISsJgrZdk9LEFJDgBQTh2KHsGWSE47E0Bt
RInrWPW34WO0DKTRSKSvHvZHS6tzuQyrPd9Z2724Mxq8GmPvEkWqrnmQbO+btLcI
p8WVfDwGtFnF/mPdS835dnNwNLAdf1Eq5qBlbYUdh84sAsHfFMt2Xr7Bu6DxYrug
YsAHKj+/ga4ArETAUSEcxVT2JfC2XPmK/q9QUFI3+VIEzu6tCG4aywoQAu1u1EZw
WK+0CrU+c0OY/YQ5yYxAoL1bdUUBdjC2bFlxjCceeF/SmlFfNPnp/BhUyehHBtMH
Yq/XgjnkhYUiDBXt+1VeydlRJzbQc4IjNu+MJQuuel+53rD8A6O+dL26BFyThZTU
TSRkmcPWTcF6WKQeSI+uPGAakXWSC+ByiFlxDI2GdOaC/V6dlwIbrZ2dpsQL9zq3
euFMEwaDjfbRRbqbEoGHJKgllxzztYjThRKPE3kdquNm88+bAz3UlluyPDumdtvO
ymMqiD1gJiWxVFa7DsUoUcT5aTZG7HwxkrQnoXxxlevS+r4SMIXLx5e3Iixj03F/
m/9001XOgTJdNLH2ynDUiwagtOl6+Sq84+IMoWfVFZYzwckwYiSNh9X/5EBYLwkR
EcKMB4kTH5tPgqf+gYKmx+OsdGEQlonzNTsq0iLubD4mMZxCt3+HJqSnSkworNq5
IAyQJ/aZABo3C1xhaxTw9B6kja+iR/fa41Du6LPzM7YVoNigeI2k1H39MJCpKO4+
x6x0ez8wleb3twKrWcMmyQfyCREPCZgUn/qwkmFGky0nY4SiwhwZ5lGY3JmgF0Rh
t1RRhASzqsTwDm4k1MyrfZHKOStvUnBDEnPan0O9Km+bYgVGAzDUZ5aZ0YwBLeHw
nAGCKRRlWn2LFfZwPsl5xWGAu/9L0vX7O6mfHCPo+k5c0LwbEPem2CTxo09/Wg8f
kloXBiuoE1IRRkgZJzacU5QZtYMJVw8bhfS5E1E0cjNyL0YYXoNHPfjDJ4DbgjI7
YR2FkXOLg3idSEN+hkPDqAFXGX5zFN1CJ6S5lOYC3dx0noMZv7rt2xsBKYiN+TCQ
W3wMkwtl4JqyZVvdQEHh52VgQ4xC3JsRRiY1UAycVGxvRj5VQVCAQbTuDyWeZSWl
ZxW29HrX0UPsw9wH6SlALkpPQcw4pA5lsx391bcSEJwT5yzwAAuG2grQpFYsh9JX
/EKUXbh6BS/2DEMQsMFBF1s3WUTpCXNjxHJZUO5osykOvyzPkOd7pLlNAsMvuG9n
1FcM6/JDQX7fo2RBN7U7uQxGu/KUTcMoRWagaUJBQvPoHFAThqhTcUpWUHCsmHG+
KgN4/04Zh6DPf235/kUsYyiultGO7tR7mx8GByt2MhHHFYm42E4S6hme93GJq46O
yhAKstgnmScBuL3+NbkAoeqNErOeVe/Qpj+hMTJZiqg9DrXAJTqHDn2pb1+kpTQf
8GtWF8ODlEhSWJ4W+v99TbTyaQaI1YHr6zFzzqmsgDmKCJ1ps35mCGAqOPGw9biE
nZNNs1kOQNA6F4ChlJ76I/MqbBsCbCQp2eWfSGe5V/RivY0FeaNJUvIy0+93IvS1
IqCqjEi7NNZh6lT5/kf210SnmTauClboPTPMV+klRN8gOy7GWHH8NOXWXGcaDeIu
E8zoXORkETHpi/MT29M/qIpJA3aDHiv5WTo0xkWbtf4QiuVNgN+sRTBJaDiUn5gD
Pj7ku0C16sgKyg1KowDCDKxr50J0Lk+JdgP1WlFgD0PdrU2exA+5c74yTrEIAjYR
J3D3725AHDAcE5aAb9FCFnxCItrHh5pNKmwlL8LVvLih/gZwXqcJ0UreCYFaaEe4
4WwlY8moEcTLZL/LFGF83DtnsCA+07ipN5XFjCmGA+I/u3SNC1TbpLDagcYlFB5g
RN8Hlh+eByHyxAs/Y7G9LMNuezQKLwu6yQdp9ixLNBpvSYOPU957lbm1K0dqsODg
ouD7l6QFSukBCNy70UtkrsJQKUON24wBtLcEO/2Wh6jVDJhnmnhvZ9XkPqPbEcWM
iiym/pLj+1gxWpdeF4ngtWCDNcmBwdZAQ8TD3Kiq62ymdYiTnN32dd6Tawiyafrr
vZHAYg8JEj1dhkD8gIEaJXPhxAgXZzZrFhYktaqvnk1pxGulYzCeGik5pC1K77QX
x3xDhtE9HUeLOPBFyrdYOZf14tPDzDMtzFjqlC8YPznT1TmKbi3tKUWpVgqm3AO+
a/XT3rYxH/fEqMleYszKx4FFXaIjxI8+skh7ctmghk83aJm+Lg89Nax/rXQS1eGz
2oGoMsYvdQHF+S9VnHPQsJbsubd0TPUEfTWDNq0Pqo6uxtY3giLLav7XTcGqk/AC
bb5fTgNVmKJa0yvhwWd3W9eh7uDifSpC/kgFs3oJ4wouWgkLQ1/f+SJASu62P1/9
KFicGthY1TidOwqRIasZ/5H4eSV/kdivFVexiUolGFqZ5lsJpNz1zbqDY3wdx3FN
di8nhQ7RjRICVlTN33lh4V7OxjAKUnOo1sP3C6fSd9ak3a+ldIe2f3WJn0qmDN04
0gVPYjDylhItovzCehOOuT9e6UwckUWvQE7c3xwfkUHCsYEOtkTLpZngwemWfezx
U4EppJsU9SFKzdCGYV9EXv14vnaSZx2XL6Gh94Zi/zxzauUNi7l8LH8YMINfqrNd
n7jtrr17000wzkUEWIY/C7/9Pd6YP70por/x9hj+oFWBbnDLps7CWpn/n9eVUmWH
lxw/d4lMOa7B46+TKCjzHzKURJWDd+oSn8/7TjT+fCN7zZzSOuvvONWJbQ500mlT
nOUqkzMsmziMAKrAWHi9qq5sMIZVpZ/CQVDXJM+RHAbG1gRgQ7mzcQ9nBs+7Pqz7
cwKWwwD5fXKRQW970KzfWiHTH4z+sytFQHRwAxi7Npj2wHRejT8hbVynDugmAe9N
YgkQIjRyasM+/cAQoRXhAHVDppBJbCd57L9vMfJ/sqFo0fs6/zoSiZuqgpftX7gG
0+IbNosBONvluViHME/ckBY5VjRHnYDBnHRJboh9fmKaSCikpgS6+qsKDIBpU6ha
Hzu1CSMMMSHO4LnQV1qX+kO3hyL3SAfnZ3eH9/WU2/JmdgSiaGfdUNsxT2tNcUHM
eCkmC3Qp2sRaP7ezeC348L7kVID/oFp1Q6xxtw1wKTZpbNYdSR3mg8pG1hQiwKnR
rkeNX9zuHcxzo6gbSz1N6uls8Yf3aIBnxXRCkxeQIgkFG/RsJ1SJw6H73pBH/iPS
gJLKlfbw5kxQYc9XKMoZWWtd1q4pMm13ShIe0cs+vPR9Y5Wu42bNWR1yHpGjS8lT
kDOv2wKCGpifNPQ4g92RsH87bSfVrLBTGlK/sbcvZvg9dcTwcAttcKut+iZB2OMF
lYxyo48rrqXGJFhRpq2QvNutwFKrcU2a3c5V+SUdr039kGkzdn7u3KgKPvwxMf90
yB0drwvShbiAHcVe+4o2YwUpC3wS5yL/4yXe+PRvIqF/ItVTVNZX9gX8tfxXyHfw
EFIsTHs5R7Zwo1rRwhaNXr+HhHZNMmWA/37TvJQ6V4vT7dnge7BQajPI78/mjGYH
Wu5wrasCEDz436b9UVIpPvbT+RfZRTNLUP/sZb9Gs5t+TqbCbLJUDF4vZIMigViw
4YETM+emmTTA0oblZ1fgqDu1v6m1NV+GkiEDnf0c0cuojq/Qo4e1aaXm0IEIulwh
xLiXasOLbNJOwiaD6SHqta6TSoNbRhgkBeQIcNV6ms6s15JBuP9+Mll/8swnkBVL
ZFIy2WRtFftU63li6Y50IeRKzV7exK+JF4YasSmbiicoRRKu67WjRE09iFpCR5nE
vuhpELkuowSuX81TgdyVZ1mY/9HSgI3Q9byVHhwhJ/SbsB7c5XreSQN5Qz3ijDOm
NyUXMMFgtEwH2o4Jv69mF1ygUL02RNxtTx7xj8Hn42+p9CnRUJCY+Sv3aOMaL0Sd
P8o6Ra8HQBzZrwLME78uZn4DhPiKtwGwjugZau7xhJR2Y9w9E5/37kB/+aOwSJIk
+Gzs/KyRQx3ajXd6Ube29aFFsG5YjeY9FxIK2sKuXrAFWS3kQ6ExWjvtB7TARO2N
0M3KtZstJJOBYVlC+PvMS6N1dGI5N85AG3lMhkYzLf1kR68aC1/3W/WaKWd57jUX
le+kx8+XH8ysDoMEkJh5hEPvv8R/RrnQzdmSSVkcv0JD0gdtecUc/J2b4wuZNJOe
AaGrhUdtSsH6YBtgkhDTmgQKJp1qII1x2iFy9/n2UIeRPmh9oUM9lJupFpjxkvre
y4bOta8qnofGhXqe5d3iDohCd/chLgsGMStqjA32ZkGKlf2E2xYd1vr5GWhCwasN
eljjymLzrpa38ab4raKpEdfAB24TbL8znIT1um/kGz8bo5owPymbi0/1s2OgQ9hu
AI7kHywDB8M70WQEHJJ7H9ryEx/3zh0kBw3zbQA8ApNKiwAy3QxCWzfvybtFrbHF
kGszHRe4VW1I/rWcb85Fk/gWRxGmV5pmr9AN9Y5rvsLmK34UDOu0ImhBN4ajANXT
qJNYMgi9JUWtBQMCH2wrCn9e6tTsLwjR+A9uxRhK2+xFo0Os5rxGPsyn8dNNQNX+
PLXEWW6ALWr33fJTXsRBHX1LUWCT330HNMeBmKotMi465YjUMr0DYUZR5kvI026j
F+NcWZOXUiY8C370Cex4sO0vQtAOQh3z13UWdG+0bWX9sxwtISNzkCb22QWtSuMW
kUlwk50X0A7PBcYyUnfZTrbRJZF0d3agH6OOnTAHSMEvaZ+a5ExxcerWdQSpqOXx
wUPLV47tQq/aD7Kx2ris/YboxpkvqfxOYxGExlFVskJJAs2JUHmI15rHncZLCtEt
V5nIncqidijdXR5U2DP3KVsMcQi3L4S7YFXhR/xQs6/BSdj9ayUdkKrvI9OsDMu8
PF8+h20Dfb29f8EX1HxsCnKSDYNjTZV6dUlyM94AXUgmg3MYZUIWjryE1hg2vgVD
r/HTwzrV2shZYJA6mvzcalBZYg3AdGzSGlU/oqDrYEYSU6zH1+HQ2IAcGn56/W8/
CNgPBFtqqMd7FFFphQqawKL0PLM69wPGoT5BoeDvxXZ3rwSC5/Dbdw4XXmzf6uFI
9qDzxbgHM4sW9r1qOfuPm7izM7GyFmQf87Hj6CXBa7uTTKFCstOF9x7METv4w17Y
27GAn6M2lfRFUAzApuW+/fJKRF4VbWfZdig1Ts3UcKVL1Mw6uuu/UV6C/TJ7YQmc
fX17EJpEVA7CxFEorlGVsFpdE3kY3nys+EUX971lJPGY6YCiwylokrwjg0dMrr2S
ofkHlAlrD2IuD1YH2mKBdYPDWpgMT2rikROVzHPclzBRzOPH3k9AwVY2rEQM1RwC
v0bwZ0Q6/2lYreXDWTjayUjESimMi7X1m2vQSfqKT3ONStbxD8o1EkLfTWYVFLDQ
gwcq/5DfSZl4OJMMjJULtrx6omtnvSwArr9e8aB49EKBPvsMaU0fpDUBkos4vDGB
Xkull5ZdPXx3QYcFm2ys5UkULdUDYHRDkXKstA7Q6/btedpIev7EtEOyIGywE+WU
GTA8SkWd2Au6kQf10eZlQ+cDVcXGe+nc7Q9s4LGT+ry72z5XuPWhO4qCi7GeOYVE
/0VQizYXKzy4ULeL0hEFnUE06oHZAqCfoDUayBT2ZdJwtWmXTIREE0kmUkuFJBr3
GxWZNmv4hyHGsagZ/0Ctsip1nTMVMfL3dnpfj/hcPBfvwiauWxKlOa+5H+E5mNFZ
mL4T28ECGs+bKk3248gDxqygSQzCdQJoAPML0F8gCw8JsvfKaZyRR0UOP6irnj6J
LUKe0oe898fYFrEAP5tYkLQ1r6p8T9jeWrfNHNA4fnstazj1Sqpg9pKfJrWYxa3G
IGz59b7xcxK/NAtKxOIp5vzfpBGoFtXfYOXepYq4rA54Ah34Adn7p5RAVjD0cuaB
Cts6q3cCDbEkSoLVmQA+cjCEmgQQU6F8lA2EAAC9n3cz/80JaZjBUrdpwwgG/NoJ
ousmF0IzdwMvne0NEhDXjX7NABQeDQXOYA1ubK/yO54zTi7USh1gESXGZqX/eFTy
uaEr9fUvcyXpTMQBttdyB3MttnW4NmbPEoDIg2UY4DPkvut2GLRc3QmCYWDzPyWU
vbXez9Lzi7qDWcfyYWcYfgawp1OWhVyDbOxzveyCbLnBGwsGoG1sNiK4IN/Hzqm7
yPECczbO06o7iY6ui9TvzBsFVr6jpv8mhRPi9jFYS41u8yimJX6ibqt7bC5sekfU
1LO+hhXLG3iGGfgFdOoX73k8l0JrFl/rv2L3UJ0wlGbYb21v6pD8+Liy484dh9BN
C8ORKR1rGJWDgS7zLnfJSfJm4kjc2yTeKrliYxl9iwcHIdppewrEkp8rKFiVi68i
4Oc/ho+V24GfImyBKTx1r0AaQ20E5bL75IkxLQ8uxGiVYPgVUSH3UH94+4TTb99D
vhxibsLqmrW9rkIq0LpeE3t8IwzxecHZ2gNb0+t0T2WMHfYgPwQnmfnpVwKmqfJB
h2aLRhAkj3tX5aieHH1zmgG+YJamp8bY+o5mFC5uZQkv1l5OOqmCKZGsz7MJuGgW
1ZrWHIv6ltQ03dGMGbMOyOO5c2xCg1UA8jVsqcfGr+TLhGNhtCo/V+yBN6jZ8fwf
V28IJWjUjzzph+Koan8vTBVSxMcTdxnkBoiZIFKRQuAukSztcadtuSzULuwr4750
kiyak2vKXy3r3VuyTXumf5gCt+euTc2kgJWvmLAB9BMLAm8c4+4yj7q/9zPLPKGh
zu+t2JCRJ4I1yCwh34bLCiYm0V9ALtkwrCRl0dcwlcZr+H9eNYVIqDxQTmaU8uQz
tgS+TRvvXDdZbW3Z2dmxswhJiugK1NgAP3AWcxDqafSNAIt+/1/YDEblcpkC8ipe
B7BfsK+kXct84YdJRGzNlH2xekl2By20ZwjDeRgY13LdVzFTxb5Uz1MXfMjNFNqw
5GyVnWbL7HSJJVZFwlUy3a/TNTY3UqYUZXgzEMZiuKhEFM/Y2tVBrwoU6pKooPUz
cFznucxRafPKDlLlecVdGGfAuiqK/81lCu1FQPOUvy86UTEMp5e8y79/2eLJ3qW2
NHPeiaNAU8V3M8rBDQQhENgZi2iwLiKWnqTWGn+x2Kuekwdd1vWSlVodae4Qdn1E
5TYR++lIqsqlP6BVWi8kRvYwWXpMshO2jDeIsVDfmFq/sx9+UJlNL85u5pMT8Uc4
9t2LVsc6DD6hIPJO/Q32KyFwYiFmCWOK+9pVxwZm/lh1nHKTeWGzWKp7iQf4FhC2
HgvKT8qG25h/0iGTJXb4j+Pod/kVwh8hemBdtVRvMIk4IK913/iF4o1ZmpC7IT9w
qZfDrD6uuvAfacSE91kaFGWzgT4TOOu1j8jFd4I9t9/vbsXEGV/pwWgH/22tZ5pw
KjqLpAM/8zmPHEKmEpJTZ+W7nKvmL6eprrZ1v4Secvj5h2dGf+E8mgplsdyBT0xp
jYVeTrSkYK21xTRE7JXEKmySApHV4YknMYtt25HuVvau8FSnusAEt6rq60U8GRsf
LXhpbjdgN0cWU5nz69+kVul5L2/olLtVGvUWq0czSj3T/Dt+Ly71MfABGuXpjnkM
wdeoYG29tmVZ1YMbJgLQn/0nNFLxHOmH0aU30X/Z31NSwgPej7DHNuYvJjdc2kkq
YqYSz0n99nA3Nhj8fEbOxk8jeLE5YnVLdJzcjL2ieRXur96yVf5UdhYbbJt9XE65
nbhPiHCV977fdsUICSLoK6F8KkSYhtmPPi/WDmB++9DilBzLwH0WTFoD/TlUvdob
/Hb5W43LsZyvAB//tLOXXUvvTOHu4gXeM/LmX1Scxf8zGV/+ap7HE8v0SBKkRqoI
xoBd2aIkfH+006YhmgLjwFiRmIyyFyvIDxHI+5c3nlw7vE15a6KWTLqPB91PJ4RM
8mSXDhPx1oP/rUWa7KJni4cm1yrk5Xjb3b997O1dpCZu51VpkgeqcDCHvqdTWx1k
Zir/OGdKsKv75FrzPTlQ+oMB5RgYlSoCG/MTbMPdniN/pjbsiJGmh7zJNnv/4Vsi
S1ceKEK71713NbQZvBBn59YJdvkp9Ktdfg/4T1xfBHrI/wL7ohbBdNU8eiJTenfY
SZKTcNfoEn+yQ8tAvFMOSC6QnN8O4prPR7ZtVcjCsA2W2Y68slpdngWWP3ga33Hf
Vfi/C6asYQOwyd5IY/DAPGQvg7wFuleVq7Kh/xMrjAYd0gp/4yH3q0PQyxYcjCEj
AKYLAtz4LJTPBHKNfgn8Yo3COAt5+gzv34MpNVxqUoMw2sVXuF9G1blw/N/JEtwB
RcXKdfF0VB2edfxyc9LORv9M2lkhhzokXvlHopvXO9yJCRuCySk3h+Ob1wPVN7cn
mGl5jq1FxJvn9b5uADvDWmYuMERTwJjoeD1P4iB11j+kXD8VMTrkjsHbCvWCAoeK
jzTW48C0xn6ZVvIyKaT/Ft6c9/gODAS7mvl0gDcqlMWUJ8gZDRU7bpq8f1T4LZpu
qPD3+ZhnoKiX22/gO5B2ONDEC8lW5S7yvHUbLY2cVHpfhWHOZ0S1eZkYEg+Cq8d0
KNF/pWzgMQt90vkaBnZr0scW+l+7AtPxY0yE0WRNls0IhmKaG+2ljvDtLqAor/WM
JOUaG4bRy/uVOD0kBFwRCRrDoQcS2dfivk9OVqwVGfLhQ8xBpTGT/hdBIEN6e8CV
T43X0vdQpVgdGkUl69fU4B7fb9lO5ClNLhMrKDsn3Te46dMrv8wAU7R57cuAPmUh
OyreAewuvRyjLywpdjFXOX+GXz/K1IGmZaHzzSMPBKQgGhkxAhTn5Sryiav6Vhl8
SZr07YZW2b1jgfI78Cd6KlOdh2UPMAQUhpVJBcRmwpfjZ/Vl5pRLxIvWY3m8HhId
ypR7680RkLhoucDoJK6Y5VIC/dOTqvukW+c5lz+UFJhm+SSK8jY+zpbhCCUKPqcr
5ByNbOtzReyqrdI5DjehUCJk8gBehRuHaVKZ2FotatRCKCWrmh9JqJuKsLC2+zFy
IO4WT8Kl9Bxo+fCmOVrM2QH9r+Lowy8+EZjC58q/C4twIHtk/JIlpbd5IssrG0tt
Jxx7pPTUpUNiqloHaBAbA+5jdEHtdrOBQ0xaq6mfIME/o5aow/+zB0W7snmAMYFz
PMP4uMY64KwTs73DXmQ7FAXcULti7YPzeUav6HjqQXVHIADdOxi1+Cpv12pr6kju
JeCDRlkFSsUf2UtiZOUN4YchxYKH3w5o7YjdmvXQn4M/4+d05u0Pylv7o05m0wdG
a2zPOOiKFKP04jugzy5dSuqNteD0RYczvb+K3UfqtwEAryKV8ldb9YgfNVaHZeXh
/INmom4TtSwlnLRA2zuFmyH2DYuN5s/a48iYm+z89Fq+zjW0JYv6+4S+hUADUdHS
aqaP9Coz8YNWt2ON8EeUhb9Wpe4io8GPA6MMQw1KY2kShhXk6B1V/gurRtbxfr5m
UQ38huOK0HtYX4eGbohEAl8m77AhrtOMn6F2AvdkYkDHb9TTT6YIS48lLu+Of9iD
cJd1PMYQ7qq8uxscF+hgi3vyhIjso9osiufeV0CqkRTMY0PKF/S4p8v8KT0fxXND
P6lCOEzdcK3tWpUdyZ0vZEQU3x8nxddxxumAVltwQqh5d872isxcpyOsG18H3hlX
3pR3z9YIfPHnJGjkH8MeeLQ+wwM0SpwP7thJFKyVIRN3H7uqngnQDaCzavEPYsvv
smtxxqnnhoCgeR7jZhZ4cRacxQ+VC+AUWmqgHX9UT2r23gspcDLx7SDEKrPH8pKN
a7UC2/dvfMjSGUbhLIYDveHAyvzluvNybRef2yZc+bQnlu7M7n8aj/P4uR5KUlyw
u90Fp8YMHzyKi+C5Jn0mihdo1ucpnHBfVi5lEApI0toQJUGmAv9T/5tRvp0P1mph
gFN3OtVQBnWOj0186omxzNRL5zX+9CBflKrDFfKWVZeb+aMbvyQ1ecVvWzwrJR7T
/8L1DrguWoT/rSPvo4at4SFX8++ovB0nwngzbfpdUKerT42YcduR4j+0nGlUeKa4
LLlDYousaBhkjSiXsPYUdqMg2hbuFIoNC7HSwR9PcHLL7gPtEDJpdFUQg+ryqpKM
JT7AV4RNWmtB47OOkwJFCuQeWzTdZale7T1MFBAUbAvNeTHNlABFSHeoPL8GTkRr
DkrbA0M/EgrHG5kyPl9tW0kcxxTwISUA7ZoALi2isxm2cOm1EoLcJ5gqQtPMYZ5/
QnXWv7Y2cn9xaAmzGIDtg5+rkySmCIrzKtjvTKYBcvUdNeFpnUxneuzDI7Ojlx+b
lzeKJFt/0WRIdttgHyMPXseiBm/vT9V8gPaRxERLFImS8/RR73tCpBZuqI2gDBEO
ZxyLKLG+I1lf2FotwEqjDLsgoUPzbs6wSDTQLdCMnYrEfjWnPc0KKXUdljhMllYg
TOAXuSSjU05NkzrLdD6MEcceUwWF+tiKOlD2IWVzER86qWvSTrcHpApL68WeUa/o
D6Is2E7wbe2U/grEo3/4hQoe63aT6qxhrLQ937SriUgQdLQV5gOneyemguIO+LId
Ti+pH6ML026uRXkbrVKVCBr87mGI8ca5eQsEtpZmT23Df/jCkQqEIrCao8qTcAD6
CP+O9X0Jb26cCEmiUlAI55AcyZWGZGSwpKrTaZpX3lEEcFYFUt+UQZTav0mmXQc6
HYqWgVYEdHl20Qo22dZPs83LDkrH4mrprAHcc+msd34yU6pZuncrGFUpRS+2Q3BJ
MQ4iSKh+MrBvAiop6eXkVsM3L7aMM8bBqTHixShlmwKljggaRbBwzs1fWOhT4KyK
a22txIAkQWd+SNZX4tKOpGD3D1SLcxawb9fbWI09khuliqHIUI0Y4EoJgG4tTubK
0vKrYKb4JVEnbldn7J9BMNUZOR6+o9SNwByrJo3b32SqzBZxYFdhoXUh+wRKvgjo
3JODdIbDORRkkIXQHdo1I0JcdmMQkGutBTwLwTCVF7mFdtxCuHfLbV9FUby2o9oj
isKgnMsHVdDkQjgcrmNa/B6kbklAZoNbC8ro80Vyzkp/9Zf8tQ5idoo2HueQk7wj
9A3RORcsueKPWQ9WS93jYJlYMDHmLz2oc86DQaPczbhHUkIboylxQLiBqJaCTESG
52lO8r/2VDgnoXQO/LrDae+gqiPNZvF1J6qszRX1zTJnJjLP8wg+kyrDahMdKKac
xoR/xs5g5lsTUkGoVJU5FdT9rHtGAQapfha80UxNBPwCFOygExknOFlJiLRJTDbb
79PdiQ6WFmYKrljn9mBh/kV4uWxX8Y2h/L7g6uFoMhNLCBcE2Qr7gJk52oboSo+6
IipBlJ9Rp7G6qkHjollWDOiYiNmBCuIhHkxL+P3RBg4yrm4J7aoARbpZIaEfI76R
BXt6UgJqZ6SYAC3tqbU45WMTDzqGi7DRHHu+iAc0tzhaaxi0c8wbwGFVMGNTJIn4
wvehQR7WE0ldkVKcKk88inSADh44EXhCgqd3HtGNknZaXLRY2WEzMvQcr/OICVe5
YfdYs0fZcczrDgOEj9PiQo9vB6cZ0KPyrXa7vNc4y2UQLHAW1ZWk+g9tFjb+O3W9
higxoi2aOfjBSko56HuFctQHes8w/55h6sJfUhUea7tBFbvypRjMTs2vaqLB0Z5p
+FgRZ5vgLx1CVI3CXJIM8JMMzuTq58wz7MDZ42d9cDCDDv0eJ5y6m7426V8mzrHf
oJ48s+BP3dYSW1mqXQMiVvZlzOQv4RnLgP9RLsq7Yjnc7WTg1PDcsX4xpiFBMsDq
lLCIFLFEmQ+zfBkpvVRLFzmluWxfa3ckFG3guP+LBsOVMN3GTrKe5uQL45vjwFEW
3LfKzyKwMkYB4Ci6Vv3psR9xM6/yyvjSelg0uHlkOEupmpDCYWf4giMETt5iRZfD
GmY7usSFrTcqVOafsoBHvJXjSKt8ORjZDWzPMzIrc82Qh/Teo9OnKkyQ2dVAx2d/
wO2YHrmziWR3r925JoHOoSVHbgjPCQme3D3KrGYryUSuUlguIPj7rAT8+6muVjbb
i51iuQTNIBm8AGGgwB9cs/pimOYfpC0f3q3VzdrgxYdWQJTRcPZeA0iefNi1D7/D
v/JqQ3KdJN2Mb9m5I52bG3Trk5PlsGr2RRuWNvfAI9vVrDbaEjrxhjfzMQvh35p2
D6wN/JNuPyr6VoiX8WFR21jGwygUSwHmXrnUs9jNQfJD1a1Yg9YizYuZv2WyYZrD
RMdH6E2MhLWrYtHK4/v9NM+UwHD3IdHGUxZaBESAQlziFCMs1Mpx3yVjxijCWlpi
7w2w9NNcma0pUQJrS38G2p+js4v3Uy/dM3xq5Pczc8FR7uqRnLmuv7D2HyTkfeNc
4uvirv8LiO1w83O9MLCLNU/CEcBpNRlaJH3HBpf7n2PhOKJEkTpeoXKfoekNZmqo
cIKJB3Eujdvhqcz+Neg5Cn7/7cZdKxshnrtA+MjuNDQ1vBKoHipQhowXZBRofcov
3IDzkAU3picdRx67x7uLO4r4RqeMgMilBtwzZC4cbULGDNjmer6h75nyBSpqlBj3
dPUIncTgiWP+V9X6fwgJreZBKgcPRRext3QQMj7CEvv83ZVbdlT59j33doWzOVvu
H+TQyUxU4paIT4Kw17WYAxRvqvsqnShzNUII9NnJZAWNY9o7oC8S5N9EjssMAOPF
HsnwLB2pQVBXAB6I+hIXHVJIM7/uSF1oDTrV3NKV94kTa+U1IogQGvTjYoDYKiaf
YZbXHv+o114zIyxJwpH+M/zl7f5WNfn0s5xSTSEqTCt23Db+R58cbt5zXzpqDVNt
J/1T9zu3JyrEMAiiJU+LDuqGCsEjBfo7EjqSSrRp5Hgo+9QlrCyU6pdCUCYABVEM
G+G2lmTq5ZYHNyf9TmzQEQJwSWFiLTPvNE5WUOQx06IXuwjqvYlf7CS48TLuO6W6
cKW+con8Oo8zQqR3zB/8qAnM9mS/qpzvN7MsHR74TUT4GicjFGPDU9XYAJwsP6iz
zoWFXqXcFcBWjKyeZTnIpuj+3ZEBYcb9EbhUrtFbm8KB25rDFu5iOEeFaMUnzjig
+fSWjze7Q9AIijmDb5k+H05s0WqnBJoikS10VJsSzaoXtVnCHCv5Sup5MMS431m0
y8ssfQEY8Cmw/jql+S9+OX6yPOTlc6ZO5HWDgbCE24cTEM3pNylXlNtoZraJgokH
RF0aHJFFL2GqZup1v+6a8uAR5+BT2SveURAM16r/IgGO+xT9c8q32QywPF1fYjkc
lL/Tk8gBmuSWUE2sCzTfZHcGY9QKNHjLaIc7znJ3mZnMTkl1tQGhrCyjqO+91J+D
PsEIMkBTPmOw7Rvw5MS8nujbw0c8GnNbPLVXKKgwkUpcxE1WSRh1M0SGnMstx3b8
3QwFRpqmr9ilJQXwFyw//BE72TFN6VMs+7XJf/YlDO/tNXIlv9bt0XkVg3M1Vl9G
0d75oYSa/YtnM6TPoDe8NupfC9Nbdtvti+ZFR3Ok3MAPG95ZqjDK7+BOK5hD9tAr
gKsl5zF35s1JhNfLl2od+EtsB5VV0j3OhMF2gwgM+4PP/FZWKqpIj7LXistY05Xr
Kd31apCJq/YCmrtoiq7fYeC7vjQiNbRsXA4nEJObriZsOVFeakECQlECv2YvFnmR
Lgw/qWyPL6TrznOW2CWH3BJpLzH8iINsEPEctk6zJaGkY9MkrQHJOi+2O+a1VKCa
ta0i0PrVdMNBxJcgPdDkb9p3KAccqCat7MEy+mmTGB7zyFPqt8aW1k03TzEEFGOp
DN/WuSdnSMGTenfeF3v3gG6kGhhe5VnrM8TrMvpOOaz8SEdS22rJLoap7PE/zN2m
xaaZUz3Tad1czsSVizjffwsc0JKi+rS1CQXQI7nTGpzHVBbC//168hR6z2UaFLe8
Bg34k2T4+UyAtUqSEWN1nNXSOdQDadVZ/MwQO2eDTBgDn1wZxTV911BovEcFbKIR
L2MOZEd/eRZFv8Ym8t7W7BIaXyJgWm+ERKX4W853qKkDFd6D/1XpJub0WVCflJvr
i35HxzFLIdt4OF6T3nxjFXLKKFcEdh7Knc9vPaI+x46JhRIaFkou+n4TvVb2znIF
CP/c3/iOgFGyUpQOfgTTqHR0ujp4m/DuhwmfUugVa1OasyuNWfDmp+YCEC4H0m2d
F+APrPj/5OPAgSnN5PL+NBkhdZ1Fs6+XoRrXC+yczoTF5BGDzUZDXzz6my9fvl3u
b4wEf2S60JxdhffryNT3JKE6WiSvmK/01r+ylwTcvu6kFCbRu2X7TMQs3prOZvZ/
4czL6F7GjAenLPL6WrpROczQmRx26QZxzV6djcyBVLTj+gHGVFBUYd1+kqa5AYkR
9mS5yiJL4UDLz42YyjlTrTHfzBvQBLdtnNzAsVBFa+TYYn3pONg1PzUj301apErd
eMq6pFfhymjz48gJxHIrV+lrIxD0mP6c+9xq+ERy3i5mlHGin7bwY9jdiPjnTlwF
dJBIk0aJeKmXYjNLQDCDKRsAiht97+Fr9aD6Sm8ejVX315ljzpFMtlC3000x8UIZ
4hJ7aYmgRiUvffuBL7zpOUb9gY1+Dqs20o7Dz6rb3I4LfNOm7OBHeViCp1y45ye1
OBuXIagtFydls/eIk9qVzGxVhYKhBRJGPQnOwYzw5c/9Kenbtw9rtOMzRebDtwF4
UTnD0NnfgFUG2C6ue2jW5lR7/hEWAqH217+EdRZ919Oq+Xorz8X9PRVMmGg/Qhv9
BECzEi6QGlB8vjMSXf9JT+HBYaYNUZboW5VbOpEPqJbMiJgc+NOooPPnZxmbRCoQ
dPW4NzOIBjsW6ShdGXbc9zHSOXqHc95XS6HjTOHzIfkaGqFXi9W5SBPNjev8g7KT
eo0puuRTZlACpDWYMh0b3rcTuAy207E4M02bflizhQU5y1OU9lQauLD9Dw80ZkQg
kAxJMPs9qaeLDXnMGyo8hHpAK+sQOLSKRLMeMppfzt4uou2Ac9IekQFqUCRGgFe+
DMY5KVgF9CqYM2MWO1HMuvxY4RFKG6c+7hmIPAM4IGSsly0ejbMt/7Dnqo7tWADt
0ZtlOwNNCPWLhMFHsVzkh2y1t6azAFgCTUvsA4y83PycCVUfRPN34Garh0Q8Z1Ek
8qgKLGQTUsy/I+TFxtgRHwd6TPo3cZfcQEFDOKAIaIOth219iH0oDFLflYq1U3ez
LgCdB8RQ6I7oArr1FQ54CbodrjMSozYwKPMfVnUQsPSomVBZy4rx/2djhbG7ZjsL
vysp809WTJQPndaL59ws0MZAzBaLf2t4iKKnojKsGCE6AHNDD2yacKFGKt7ejDqf
HqriNnbAoOK5voMmEsoSjJPIuB9+nvJuc+RahHoF8QTGblBO4yimgn9d8PXNBGMm
SazqWH+2nhYW2b2dY6RAfrQxZS4Y4a0IQL3YDQMrZtAmuRUALBLWxqnodmo4Mzyk
NdkzL7JVgcPvKMwjPHJy9sdQX5IQsywbk1KLAsmvw/VwI5CZYKx4o6i4CoBcAKFY
5bLHmVDo9v7KVRECO5Phr9napsCBXhz94DlvbKWPKLYdkx9PR/zOypOTUMsqloWs
43m2gu9YDG5ahEQPN/a08VYd4N21Q1f5RIqfEIjz7inW2mNa2Fe4kqgP9oZMsCFu
svrkuX8iQqxpJl2NCKqHe52sxU8Ko82M2OOdfEIWmhN+bBMusNQqfzgtceiQQHYj
DJqUXlHf1cgQL8y74FFrV3NSWNf3IsOEZbq9SGXI4sAXR19mq8/KHfGKu4QgHt1Y
1wQuk/z/5Hkvdj/gQ6zIjVUKqRuQIZjasi0HxG+JjvHT4xWu4j/mVnlLCRQKccUc
YpKXToQnpTgptcz7qjzemJzBlSXFbHOX41lrWJNyD9NmtkRzHJuQE2HBMG9d2ovH
dktA8qjnw7iS/ZBYx597OBOuqkyID0B9u4myMFfOCW0itdnun1SHt5QSxiCLV+Gl
cGlMaA0h5fL3147sTsN9FakOuQaFRb7G+K2OYomJ2Hih/iv35j2ss4bHAozic4F9
yQ8jkvYI+kALi3ttP4iq9CdUpwPItyT/CBJSAmQqWhs+jB8Gl9ECEf7Gj8z99YR3
zO7oPaK6qW7d+ZM660/eQdxIP8g4kh+lPLe2/0optw+jGNgXOMAcJjirl8oXmBbz
1OGB5xu1PkI7HT9dzfO3Ambj+L3Ysvu5bUM49AUmi2Uu+atHcSQWViwyCKMkobM5
9QLhVzGKjGhgF8/dQvSZuG2/lcfPchhxaXP8GzD5tjwTUy8qQRBLUgg+PTmbb//o
3MTCGZ/2mNwHi9gO2IavCwzlub00iZVSbZDsy78eWsdD+ZhpEPoi8ahYR95VbjnQ
Gcj8iGpL2CIFdx4dsB/HjFM7CqrElyCW7uOhJRYpcK2UK9BG4F74ktSHSasNmKbQ
Or/mfYFUDkFLV5eIiil0tbi0LuhItA3VCXMTqizIzP735JvhZoyWJvw27uYQ0vB7
o8Ibq1YM5ICTiWF+eAfqYy3x+tfUWBweXYG5/J/W2uigvQhgKbvX4lTtFVrQM1UM
5cxtQmXoPtJ3qfkyNzTM02EWePUKfFMS1N2uTOpTxjL/J2d0nS6VZbM40Zw8B34g
+hAc2zDeUGz7FHkq84fqRDxWwCh69oRJ6IyCH/X6FfUUHKQ+Cba8j8RFWhESh3NH
hx0g25UDNCu/t232a6A8P50LKeHv785K2pE1rHuwcASXuaPNSIJLK9T1GlEjKZxy
LY0QYKiDpQ2RApCplvMFeNs3f1zE/dmoaTU7MZiyJnnMzd8MH5Tvam02ocs0mf0o
9gwBBVN7+A1C0v4Jh+lOZCyi8b6wRLrrLIhco5zZQhlQ+OskT8Ld7ImCZ7Maj1gX
oN0ScGe+3QEWrTJGYMEbngp0I1G8m7SuJULwAgxe0zYV25wWGHkKeVYGI/yeC9Et
+JArc6QQYhmVcIkxacmkRSYAsAp8BgdfqP1+Sgo/EJyVoG8krSrnbMTKrr6/yr5s
RmRd7W3wflMpg7fE0EE9/QdI6DsQ83bBVtUrRiFQINSitPkUtEDaEV++us+hKYvI
nK8LU5WXdUOraJ+0Y9Luv0VaWUHpocoKpQ4Psj/cCQDV9SM7c6nnsA/drEDBg8oL
KXIZjovmaoG9HesEumMGjIwLTY18cjgxNzoby+YAY0+b7pTBLpl1i9upkOINJ0Wo
cp+5tCmZKY2sGP75bHV2e4TRBYH28nqFgxIyHR740brw8EGsD34w0HLmm679lGv5
0inQJWNc90uXndwsLMuWKRnkNfPiPddJJo2pI8eB/0OGNxQ+yM2ueemNTtW9ZuPG
T4Y5g28a7+TPjbWTqvJHi5TuH9OfT68/8b9fX0e/GYG0ztI1DojXh2Orx1pOOi3b
dUTMpxCARoIRYBCsaU0bVysxvhCFTCp4NLpAlM0/fiMVlpKyDvQSf7XtY7gPxvyu
jp3AqErNA3yNFq8mctFSPvtnZLRUbJTzUqRzlxJWb3dKowBCrpVEaBLFD3d5jb0q
g98+KQc5Bip/mG0Ca45LDmSsn8vuMIx4hGk+v0YuzNb1O3oyF5ZnvTuaIZ1vWeyv
9v+RaH+yPJsQHA/L5A2/fClOX9HZzvdMjZn7ELu+0bMCgs8cwrO+ngBGbNk/rpZT
CtR4xbwyTpos9yBl9aqTGaw3WeID2659iXC96mV1RjwY/YESOuQMENXpMdYma0Rj
mj334n63qbZhIqWuW4s2kZ+wTJXt5lhQv4GjBYWXsv1U1DKGO15nx8u/rpu53up9
ZF9afvMvftv3QR8GBQarfoeXIG15myrxPDpPlhMkWU2Ah1/Vk/YVmbY/yuDYYmZS
FRcZyX8XPN5+Gk6lmGQLmhH3zOnWP3rqDZ4Jds1E9TFtPBhBG1zXxJTphGkxB7x/
wTD5vJk9Ha7EXND+NkdSVVniFxry8/4/L5klp8/m8QS5nKEB6ZEsO4wEOjecLs7w
18BwrJYjWEqHlOBhYNO0Aj5rUQFXh1h+9fzqZ7cuEDU84MjzVXLfdgEMmEiF15o0
JLQm+08muTu8Pdt2AX+NizWdylH3QKPooT8WwkkBXx2wutYfmsKWKv4HmQpezCQJ
MPs6d9lx+u6n+31nbB2t9CatN6Dpxhf1eRixTfuL6ddhUQqUZmDkxfZjfK51UVSL
za4BdBfO54+nl3oFR1VFQGlluAGmdJX3cABBXROHLP47EAKziEvCVPcG1l4skjEW
CiT8BLQhmt9RafVHyBrV/S7mH4lE7YZgDUThAn/fSvehkS1Vw8PrXJJlWrnTSJAf
OAdxcie+Mf0x8iX5lWxV/K8QBMiB9fdUmPklLXvI/SWEi/h6wEp43YDPdLCBW1mX
Fde49JH4qyzVDe5OS5M/yhrPFD6aF7yZDGx4tBOrfP3MvMAYSiXyZMY5OrMx8A2z
5MghLXJSl8aoneKyKQq91ZTeEdCxGxLIS8tC9bKYL0CsI5GJK+9skJ2oVLrycBoI
v9GLJ9EL8TL+et1ewL5WTAysd4ACQ/d5nGz2+iSNw8TziEsmOrKKU0WSMy9xNCbt
C8UXWpEzFX+nXGEbpQmtqooLGidN/2j7DdKmNYDpMw5R6gYVhmpYENx9e/DJtwCJ
BYKPQGCnXXGj5PsqOwWpd/Vark5EUkXiN/HpSdYv8kirdThZ2QUh0grwkD1jW2XN
5FJWfkOsDPGVG3XtyICDaZbWw2z6RMTJYAUCEkW7tT6D7l2G1+E4Q6bEab1QB0al
yJjLGxKXgmH2GC0WNXP+oyKqlwznZfby6rWAN7w94eV81x4+BkGwBCiWeOTjXZzp
6RaoG6r+K8vZnJl5D3nUZ7jpE7q0zOKglrr3pahkDDChH7zFjYX0mtTX2WV38RDj
4t9UIm3XF4WMhYsl97EuYyOFcn3OyqkUK1d+sbcwZIWoJFYlyxl9PWSGOqNnhn26
35hmOx9up2TWbzZHrzupwyD6T7tO5bcR5Vk5awYTsPI1ynYPLArHY1Dfdh1uWX7b
diSGJp9VS9Ysd/oP3Iu8kxWCa6mr0FNId6VhkDp0/waPzjHQabv2Xfb8/IA+5CQL
79D2/yJ+AlLfAHXZxmjmHm3qVNcdIoAFyxoK4bUa4UsaShivQr6wDyxppOD2xEY3
YpOM5zq+JuaNIztmGTIDmkfPbdApVfe2OGXjJrBIfifSugIuHacXTzI6vKsiMvPG
ujKHuRrGZWlJbodZl3qTtRKrLRcjgipGyA+y+A83SI3TQ9lzIetTFXxONPVvDE6V
ZxiqhHh6bsMy/bVRB9wDsk7p85Wvg2nuAhmTWVrjVDrAci5B6dJq+AOchaQqa3+A
N7TH6+GmiDTSAX9sgTND2UPdFE6UYP01Ufn+7BY8N+4BzjXGDEVfWyusNFsPe9nw
k7AL2YDfHWsUNYlvydni0PlA4u2Tnpz0dFTcCBKtlhM1A7u4MwCWF7DRkd7P1t7X
XEtV2deFnNbTS48KYaCXzoWd86NNAQwfAzHvKnjDA0JwpJmzfDYiw78WywBHaUOI
p99CTqUSwlaIilr8LSNJgZf/80t4Goli7EWU5UBFaxYFX15WleEYfWDRgKQukP9O
oY6P5Oa8XcYeCOTy0p8sssQca4GMQPW5sJc9i77LisyFVcq/sDgj9xtoortPQ2QY
CEAcymH4i+1qlNJby2yKtn5K5ctKZX7F6TPtAlws7/h+swz4M+kVNTmeKdqrQx43
V6ptRVf+e1ejwwsOa5aCBHNdIEN1msWt0iX0EkWONTMHQUqnsPsB1YsGUNCO9c+y
5F0ttvTQCIjpfFM1L6XjoyCJ7E1JhlpYnmhVwGt+93rh9NWMLv2VmUdpQwfOyNMr
jTCnAmOrHKx228EMu1IStd7DPb3h+hZBybzYU/i7YLR3LhugG8o7tl6tJKq1dFpy
6HG3eTO04CBnJPfa352ts0Jyl4rT/EXR5LJF72UbIq7PnIBonadP4pzi/LS9k5C+
tv0DZr0Beh4LR6p9DL+QTvb+OHJiB/5oGz+fuRKDCM+fb07YtZlZjd/FGiMN3/GB
hBF/Vb5arNNIuYrEaB65kMP9CBLoDgaDlaqxyfUq0o8FxSNvOuXfWJxvjvOjyZKo
wR57fX1NQ21McsnF2EPid2+dRF2pZWspg9M6n0u01nFe7q3BqBkvj+XmAt4xbo/H
v9l1Z0di3LOoYydibh2XVlUEroqXeGSWv+F1u8YFYxsFt+SFfUIiPG6v6VI9Qocn
tHGzKtGpmoz1kkv9Pm9o7RI1h8fR0xCcQ+JNcePcMyfNsqmZLeYwvSBPMuospZZU
vwTzCtvX5eRwp6IFPkJg3jX/xu+fFiM2kPeaX/Ns2fYvpiznNUxZoTS6uAlXDBeD
YHw8uEudKlbFPTXaW+NRLCYD7nFr9Lnho+MTcI0vihNZ9DxTPR98zqkqP8cFTs5w
J87j5rfZtLIheU+V62YkDWjOzt6c4hqePdXo+77/2SqkM8JQKGx0zPAFeKWJFhss
v/LbDPH/uuDAhmYbqQLkc1dN2kCNwr1UH2TVM94POdHpnStBMEOj2xpFNdOrDnfw
ICepi4/0f2jWdAZn/CrcU1nlT+xW0ZSsk8onxrbCrGThbd9DmJguEpKzQRT+m7w4
FmTA0Wv9qxi3LsHB4gYnSmLL9MjUbMEUgrhhenI7hzixpejx5IfFDh8uHPTssDpX
FbHeRASq8W0LWSxBA1RFdj4MCttfFvzp8XGiKJyHcfgRqXKfn9IPBeUDBv4lECPb
vs5nrSd+dCXmnfmUxeGO1Zmot6eOlqzjS+1pgoIfiX/7rbmuseDCd6FjJ1XmNl2D
B8okuUNqOxCSOu5VDnp0fS7q6KZ0Y+BgTFH7Vo7cenRh2vFxJMi1Fdk8anHEHal7
FpxusOYvBPHkYzBhOl9RZ5CTYMGMSGGVZRTZ/2GYd5hyj1oV1QDCZcbIWH9EkHcq
HHQ318nXHAj7794eC+MCFbkbTK1OMP8rP7ExFesbbCgI+1wT7dbOCodXD5yWLwvt
ivk0u3EuGyr1KVsau5WAsI9AykFIsVJjm9o9VC88DATHNLtjUDoyrcLkhveArMk2
F3pcyQl3zO3LqbhhPYTQ4yMkBetKy3LI12QCtiGlNSBMs0gjLyicFZ4x+fXqnhxM
fJVFeGwqAavtiovdLdOT4SL0/zepMhlcyIz7R3Lr9zNlyy+iJv6rBPVp5i3rKk+z
rB++0GhEQivx5bkGY8vSk+HR+TKig84YgD9Jk5TAya4xpkaT7xQkyDpFsT24Bikw
zdi2wMLpWoG2XG9dpatas6vy9JEWNC/HGJEo2Iu9ZZnGHdQyplG6eyTf5RjSaywu
G2VFEMcp73dlIoBJnN2QYY7V8w1lB75ZiTaMP3GQrD8gyLonNrf1of+rI8O+SvRb
kIRmpTD6GSnJAUe9/GTo3b7koBzaCPzmoxsG1rUlv+R4VMiByQnsul02KN237ptp
360tLyVzBwS2o9qy0FnzWJMffS1zvgQ8p2MkejZMwNtUVKpsmHPgkAsKL9CUxEr9
uxP4sVJrDkUePrKRRaBpkz7V3moQfYbHZpzr3CxBP4omTZ4bZpcJBjHljN6y2Ouk
XcSGrrZwuwvpzVswOyhItlm/MFruqFnfjWElbA++Jf1jU0vsMPM4/CCcFuCi358k
MIUhB1gZijXl/wRqzCNKry+nLg7XB7XeWqlkoUe3dYUnxS/ry8N9FUiX04eADAde
idD+J6/9MKGXjN0Kyy07rVht6sfhqpqApc3VBJcZ3INVf6jNfNVP6Mh78d4HTH59
9g5dL/a5F1gzKokjxVMyBhBNarJNTpgHyqGz13hLL7XRTZ57+jazddr61FPNWmB6
fTCI1ErWQgkmiExXyc/+nx/TpxN6MumHc1UCLzW0AnGrqMN+ioIk/6tLxOzqq8gg
sZ3Oaafkazy9w56e/AhLuVXFI3lFf0Dq7rBGyHx+UDHNsQ/Y94XIs6kHAIzc2qNH
Zxl3vgn26JJ0Tu+96dBRPbvNE2m9S0ndCobdfnsZ7xdBBIxCocbQDIGJLEi0aVz7
lMtr5fTEYGyJrC/8rRZ2UItzucrX4jMKtEFa4tNs3YjUYFGKpz979GRZ7OGsbIy+
wtoDymK6XKL7bGDLCstTTy4WpXi3LKc0aVcHbt5Ey3PqsL2SnD90hl16Z+P9vMSS
pBs3oUV+xklIEq5/34QgmSO74b6CTd89624hudcTU9GP6Tu/C7LMyuH/M0h7dUMk
rAmvyRnnL7lvU4+QQEfD+Je4sMmQg5jrEYsvZdvVkU1Qt86oo++WB+hBlCegr/WZ
D6pAzIR6cL1RDYP7E+70FoQPY34zHwhVX+sbTQ+TfUiSJ2u4xLfGZugUtaTld8rc
zLAPSq8B8KdQtOgJ1JlZHIMxPk6DYZTUksmApu/qJ5NvNADy0EJ+XZqAOc2bO43k
NcpCi04c/wmer5Ek7DesjCazX9OpCEU1EFF7+z2vNnoAZzISOI9BuB/aXcYeldX6
6Hl6L7ULxmG/7GBQIx1xHYAeQoUI1qP4Ei+OCbh0Gi00uFdcYDyi4ONrtJsCPR+c
ptCMxZea/KLxFapJUIwCkZldGHdOTM3MZU+wTBJi9KluGuZwtnS8EDMD3SMBcr10
CzPMbDgilTByinvrf8YSRtlJ9hQkncaFjxqVZScDGkl5F/NFeiWjWPZdfWFuHR+o
nYuoj5NUfrl5NQfqLnJo+sXkWewfk04bVtxeALB6dNjEWDnb6AJF8PhleBYNKXqK
hWV6N5ZCAKnHTVjRgD/DnXmuRFpdj3d0BjTNC2zSssv3GWzkcKIuob4BOQB4+1PH
CI3rqJWmc4KQ6MhFuBPxNEyf1XY5j+QLkHeOODyUytslWhcBkISXZak+oRLz1dfA
wJuxFo+QwyODmCiwyH9RIRtM7lRxEaVbV6vPuNq0kPsOlV9tSzj8SC3bkabXI9QQ
GbDeu9OmIwC1xC2wKa76BmIGG9JUzlhQNmOV24msy79F3vOWTDKXSNpP/A/1srNH
3zP6FrEK8ZF2/eg2fp2RauG5Pe6/UhqOALLHxrTNC8LaiwEi/hMZrOZWxghK+1+p
1Tq+WKcpqihccJ7j/OF0tlmcxX7jmg7tPzqGbSFeaOD2Gylxil1UJTlsoPbfqU7x
f5RR8gY43oxltDFshpu/mY8cQYcwFptz4OXQRCMUzatj2+7z+Ec16wYn2vFq9vPX
BzZWuCr+PuYusAdKV8WBKDJr4ffwOAbD+N1E6jrL0ZmZNfSZt1fGcigLJ97FeL+t
0uFTmIpTPWJCYkUiwLzG3/cnEZt0f1DloAL0wvn9zIKgqRjx0PGX7BGUpRGEr3JH
iPB0LNnDDOcer9Dlteo0SuOjDCoovEWYgZwXXCXR6iWyLMm+JpaFZycqdhLo4/F+
mhfcBC0zurtj4+mt0xMxHeYwB+UdNiZea6vabicgxQjqdgyDL9CgWncvKBfdba3r
ddC0ZbBdYFatKYpTjQer6N2SbJNr4zOlz23F9LMJW7Gccj2XZuu2KcUxGK4UrtdO
o3uqlfkAdijoty9pZkZxL5IFC4teDqguLNB4mDrtEXMoWF24PrvU9vbCqb9k7Kwe
xgLvxCAAlIT3NOXLAVMMDBKcDKDiXheqt1+PfeFEJBD7qEzrQUo/ajuPq+dU33p8
n9BpKp5oUSjIpRxVr2I57SMy54y8rdSNWQYF0QzUNjxnexHXvKxF8vr3cAqzcl1o
WBkBxhswrz3WSWHwu0+T5gV6AqbgZX8rtsO+DIk6fZYknzPTn0A2E1Bbh/dTC1Fq
I/CXaQnJ2z+Dj9nEzHaB1wVWJKvLMVws6b+YW3pvpS99A32CoR16EE3nRGmEmDSe
5qNjcvlJL1h64AXIUmnFeL0Nw90CvJs2jR+qwFcOHM6dm+lJ823y9YdYsiPnees/
+1rE7csnImMvOJZltuvRc9AOARpbMcubrZL/hOeB4gU/L/OqL6IKCwkZ+jpi2oIc
z69hdiIxmeSlKtsJZgZz67kCOMMu5yzYWNaJFFErL0gT+U0KdUcL+8ar7B4bZWFn
9b4RtyL+QjkD/8hQC3ALc6WzlRE4GxxeBQXlZQkeTR3iyY33Nnnn8Nu+Yqgd+qjc
O41q5qTXcBKdw6i+vkASsM7eIH2LCS1Gk4Geb4rX9lv4Kj84d4ZK9c/eidoDi8uz
ZcEFk9Pldq6W44NkuM1zJBkqq6VfD56Wa6tZRbg2MwLP/XyPi/c3BWQ6IPGp0Hiz
rd0HNy5Xb7QAuKGA4njt/CirWQ9wwB9YNI6fJWEY6A/9R7AXF5OoclVktoITcbDu
ja+R6tYZFPIbhEzW8hjzwoYSjGz+NBFux0ZRPA7in6d32X+/tO8iCawm2Y5AJKhh
SzpKAMwBojcSk0q3ph8ZbjxMrO30p62BAROg6He1fk5vL1420kkmGa8lPB2iHDY2
mumIwhjxypFrfqt+7twM4Qax7Sr2i6SI8g4X/8RkpS6TGbRMZIZAfq9eqMmrS88p
7ic8LyvYZlCfo/0yv21G2eYQN40D/76oAKouxOID1EiZalbd5ifugjT0tY6SeHPh
D/9bTNnP+eiW5Brwj5ototOd7190gpY7gQg0ZQnjJpKgqplixhUjgXeIWbpQz52Y
y8ufehnf+JkPckaRqgkaLwl33brQZSW893peNdZiX+bOZEFazSoLT3ir+LDmZG28
UdvDeSJOktMa90CJ5PwruFjlk/1MTq8LsrWzCGCOTzqR3KqD71iPmQ1w1CEdBS3K
z3ejfByVML5IFskc4EMHAUNFlgsri/oDTgIaICs0IGiyJYQJsmcB3CWKbUgLwMep
orwNkymihz+J7z4ppVStV09WGUZEXbtMLVswCyXnZkg/ofK2upwU1gfiXZd5yS0C
ou1zm+fSbL39LBoAF94Jsmp8Fi1r4ND/vu1X/t1lG4XoQ4TBBY+TTEAE9L+kEfGl
vb8awxEnJHN0CfHNZsxME07EqVLq+jDGWJKCY57kRoncCobfvQJaR4bpAZMWMqtR
9zAd5YJBO5qieyCCkxTQqz21wKOwkQliCVpS9797PNR1F6zKlKiWEyB2S/iX2yXq
9S5XMz3jEMJywb8jhyJknWgLl4xK7/heX16c3YYG19qXrTRKHhE/bfdCxjkfCrNN
opbOaVwJv1+K/UaBfJwsWjCzmgGnTRDfSDtomO5YyY5JtHDDm834lHhNj+98VLUo
bqBn7h16G4Jmf/cY8/69ceRM9bVOWpWk+VUBuNfnIzI1Ar/QLL1F5cEUqM+KHyAG
px3NCLwOxe+iX9nFfPWN+64WqGDe1B8xeBgpMy/hpSkBjX1wCiD/U5f+2j4orqs2
4YvBm6FZ9IO5t0jPSJNGhnC8jcB9S8UAO8moP7dgzeTOH/ZhCblKtVp0VeacI1TT
YF1iWKswgQczFCIYrtyLbN2HWk6C8C1W8ZrTGaiVgb/SvH6fA+1cHNljAOHw4zMF
JUq9I/Pgab8lH1cnNPrBN6+vKhqAwbWXj9f6WpfWWMF9mZT/1OdKk8gJg+6pGwFA
c/tk3+3ay/pC21DMEw2+s5o7RIVUR4uVImtcbfN3ErVUAAEq4eUjWJsG0du0cZ9e
QyWxN7kSdfFiIrvlnwpIkK9y6rjqHHe3InT+fCMuqZPpcyHj2runE4TuNU2aWYX0
1s2KEzhkKo7nxcXr0WSFSm3/zVluMjII6HMPSS04l4RXK5e1O104UnZoyJA3y5mO
rKnDxV5MhRVlsE6I7nAlIpedHzi0BGQJtIBNk+FLmSFHJZGoTPLsDOW3OUli2QdK
fWw4DCYKc87U2bI2BKn+gSu0DG6pZiERue5p8Uy71Qdc7cSkxsHjhWflCOoZURRL
jDtkVmmsaJOcpxXIkSXGJ8MJ/R4L1xSpYJATTReZWj89IdgBIUTodWWDn3bHHefn
3tFUDFn1dk57W6o1zEiz0d64uK2bcDoFl7V33KX1j31UKpoX6Q49LP+hMLLUg+uP
EISjlzRr4cOiHjvxlCdbsu8eImJc4M562UQCZ4JCjIrdWnLgs9ILJqzeRG1TNuKS
av88ROoblvl5Xv8US4idjrd715TcmpN4oDGIbU6xifdxn6rw1xPBDTKLxq8695ZK
d2c/7PYPeoKSTKQZRNZgtR+Nj/5KjsIv3lvVeOgnygrq0VKKo+Q1gCPtAxnjyAqW
rLVVJX0gsnzM40JDiCukwMI91W2AVTR94VjfakSgNwKt7g3ISM8Hjam7yLgVk55Q
0XNkWZBib8TLYfdEINkZW0gh9e5bS8kGCvp4V5yVUY6GJK4UVgwixvUVQziyX3YL
+JpPnCYeONJ/Q0wS8WigK5jsETr7ZWsW/AHaNG7XK4m97D1XKOwdtM+vUzMTylnA
+s1XcNGSUoO1fCl+FL2VtNcT1T0+BjwSEyPeBaHx8M/9W65+XFTZq+gGkakSuiQ2
FDP1k43zjHdy6cbarEvoGmA/eJT7ef5GMoxJlEdAIQ/z3m8sNbiZpTZvrhkfonG4
oO04Mm0Vx2vP3mRQ/sa7imGqRD/1dc0x8bYL9vy+XJBuk8jCkker8ccK0eu5nPY9
WPjGXKzpwU2xA8G2Cntkos89JSbnlrm0MphCnN3ICD0WPf1ZaxB2jP1JhwM5Qs/V
9tf7hf/mqD07KzdabeoDynXADgXIIQqyiGmDy/a8cvQRlyWMZmFMedWb+XKEHivI
9EK7WFdl9r4k92hTByhZ/ltg73AkaLr9XT/2uppcRNG5qMFv5oUbc+Lk8hGzlmEV
pSHixbYdIRV1m/Y16rpAKkkbPu2rHddlWN0z8u94e/XSJoXk/CkQKqiA9AlJIPXD
djaXWenVC9R5X699kGQb6AKSzi8+7BKRGNt0AHU+83iO25cXOG+WSoVE8d7w5D/h
gwsP/579YO+up8VFoKLFEQvk50zS7Za3FDM0IeIauRu/YkSUIWlTqFjFCFGiCHAd
jTLHLIA2SItZGfGxPj++0qGiwQ2DlL3kBO2O90vavpwrbxTbCYkqoGZ1uBdzbfRM
m2Y2MBoZSFFbxN61t6+e3ReddFBgrQ6WpNFgZkRyJEeEOxYePShkEe3nec53kA7n
PHCnzEuC5aWgNZoHsmKbWsi8Co+gTL+IsasgG4J7xj+nN/fAr+lBM9BnIUNOl0Wq
Bnd3aIHrbqrVlP50cqgFgD1B/BVB4fZ89mMb7hjracGmoj3AFi5ut/91j2broPVj
BDppq2ofyA3M4lAEyI097zAc7V47J5YRUahEkZ8CUELPxHh51tsln/ExyULi3/b1
Rb0IA5Tl9A8Yu+/w5kAVsPzlZd8hbVdUBFafAqp1ZTs70rmI5VRsjU6L+CADTNud
63Anb4Y2VQjzVmRnRyq3ann2G2AUSJ5Y6jdsScmxtbYH/mOjzkYZtS3/VTmaJ07b
aiykF3+dIi7A7IJV/cEF8im5/AvsJGvjsaayrLr9lb8uEdzNYcWwQtlLju4EMARU
yxHW86q6l4e21V+NqtFMolU9ADo8VyhSz1a2e2VLosGxLiPtmeDeEBMDSTBBCkEH
mMa1EEpLprGgZ7XtyskKjxnAoFWK4MS82GsRQXa5gZf1+sfZTCAi5Jqmb6bfr9F2
fFq/Zf4cdORoqQNg1VAjRsaQXXcidrFDj6rkkGiFHfgwU/kax4qlXf/AO97STUyU
GM+djNmOIzgsDSZMcL8ubUyvU2r6DZzXNLRU59Pd5Ng+FTLjETGpavxyMF0FLSv6
eKKXRnhxrlzlMT9bBqiQUZ5kKFZt4piPWpkTygTozoxVUAmW/BPYU79RwyzEKDDR
J8dkPvFiULcujHO4Asn8f5SUy3RvphPuZRmmo/V/gI7O5vKFeHHg/vH1nVKya1mE
ep/kYdtQ1/1lcpNCaF2rQ3UOEZvavRmFBJm1CiH0c5YKArhhRqpK0Gm/UyejNjrA
DKzWaODHsWUPG2YbjVfa2g310XBRVmVoDO8kBMh0RLwpBdjTJIo5byEiN+LrB62G
JepA1yeMRz4mtUAalMeq5ckbVb0J2XrnEmbZTENM9lLVdvo2XgqoyTNoGrySFyrf
nUfhzK/q7i66YSRTR+Sj+eIkfxyBq0wBlRFdNYJkNp7pEj98zDG73I2Zv6QjUOT9
QZGSfBPGRKzUIj6YKuD3iKGFMq4GnpsCrpS+oteglxTVtUWwHI7zA0bD1yr6vLl6
F3WEluy3r4jm2+fQYjFjJxokrMNK9cNdjlDPsXa1G5TbagizMqQAWLSArqdJ3kN5
57Cfa2ziOsT2Ksg+yKgjRHJz/lRGzE1YrF7L5xGVurifulj+L1IKxVEQmkvl0Jjn
ebTwW4yf3xyyU8sM7KqAO0mdhDMeyDAU1xaABrkzfWDknXsvZwThAeN72LzhYTvs
AxL8hp8QyB5P5C7L9nEGD3UdeoYl9c2cVkmpb0dkE0WxicGOfIEoqrsdGh7GXWRU
kjai2+QaMPpaMQeqqNvWuyUMHlfnooaJFaRu0zjbC3g5OGjs3xDV4IDFPlUmkSIH
ulx9LkcIOvLuRjiGTDomEVbq5HAeJTr8OsNDIhYNZvRB95dTqBPLKDsaUg+5k3nC
dk61lqUeAXvNI9b927TgtYh/tqJhFjdqnQohhw/wpwTHcQf6MCEa9+i2/D0pSR74
/tccIL6+Xyca5ugWq5/5ikoUSuj+vVVJ1yXnDjN1IPzunR5lreidOGE6pzOxcZ6T
pXK0yi9qZFfiR8jNN+YSMTW82y4cwdPmlbFOfjjyAI/MoIV9uDSnxumAUOW8uvDV
WMsUduXmvi04ATkmlA9D1JTxRO04alY03ytKjPx/bEWzwcjhkQ5mO525oXcdwHwa
bUmh4N/L4x4PY3H6Z31lgVufip4J2v+ggRFZrLnHE7t3Cehf2/FYjQWBBm4oaZ5K
Cfu8gN1cifxky+C5E+6NQps5a6DExk4cvTZaMgHQtiRpFRx9H49CWbYXavFO4imb
TtJlCAtLOCGeBo4qjhIBijXPZurEs9xrf+FRvLuv3jnF0OnUZ7JOOWgQSAsRYjxX
6xLyHS9+6GlfJ9f2AckjJO65spIZjpl/t6OZN2uYWB5Dg70pKF0DsEt8CvpnqRsp
gPn20bmlF/QX09NlbhFdyZZRxDyFBD0zRDCRI2SQFqVlmllWgqUGBLRVsBeVxSKh
OkOMgx/7d1+RpbIqfDBXceQQ2zp+G6iFYeIlYTb79K+4h/jUdYCh12yGM1mWGyec
E/dUbsu32i6lAuvfbNc6JoUagk76wPv794AI9w4B5bNzAH9s29a6dQlfLbEqKlC6
8ZszElSEJ8Pjp9EJRmzuU81479Mt3hc4ysRvdLXFK566rRsOm9Vud85tric9MDN+
iwxsHveCpRYsPibhQSj3jdASg2NB6JftF0WEqUN3CKxIxryTCRlUi2+JlPzElXzw
Wyw+gW7ytyEu7Z5Eg1Pmrd17pjbIIIDAQEyKOSUU9NHmPSLvBGfY+7tjd/xysD/X
xHzKBMh4DRuTYW+jUMO9dtfCEFXAmhs7xmuLaKWCInDY97YdovrB2s+sb7Y5Gkei
ddmXyLnRMX1Mcc6gZQEs6hiMDnGwQt0mMeJ7p9hnZ2LvRekGrUk9bq35WcxQJ4MT
VhnrQ9Knf6W77lQ9u1OOP9ZQFRnqX8h104O9yZ/7EcKbGf1PsumYNvEooSnZzhhM
qGQUPYUHRMwxhQxqOZI7YkP3VNYBY5h592XeroO03+U3torsGGynQ4GzGEb0RMNg
rvyhSL6EWIKyBlsvWZNaOSuqY3aXiwRUnWqpaqrhE6abHI01xDVyAw7eXqwdEM1R
BZQpcBYF8ggfncZs36Xji2XKXoMBoiaUJ0WWceXNJXzvCjEqE50p6041b1c5Ywz4
JaQCUx2G2HVNms0cSDcrp7qondAk83Ts6sjq7HK0KzU9MZjrsOBHUn/54V2eBIwQ
U0HDrqzwSzEgSkELq4FBymIVhnG2pXisrn5y5gp3GrwdPfwQr5U6hae+ZbsREdB9
Sj0HUMboBmw4lU8/6wXDJVue8vckgV1bCwmyRsjoP0gM4UznwB9cv1BF21N6TbRQ
yry63ZwU9oB73d7xeDvX7aaDsXsiArOkZ7fkJbXOLYsO1PXuKa4oCPxnOQaFvzgy
EFcW1Eo9XqBdtNQDzQLfKylzqPAuHgck1GDjGzI2IOwdrJfxMWS/1nEkBIUb7AdZ
/SN4X/u7m+F5ZQQ0kU9X427l8i/DYIV0u19vMk7V/l/J9id4cL58+dzQfJ/E23oO
wm2BsWNS8JFAzv3nbG4N5s93IF4KCSzp1GSkniPJmNSRBr3uoak3VSjgn2QIsYyn
vKl2foQIuFXzk5RNgGKXR2W1BNYPl6q4cQIrE0P6cLGnhIEvbv7ntSTR4t7iqdtC
RNWqtDTi+Z1rlmc9WCfkvFfM2Pvtefm/bzyMDBmDfoZGikZuAkfXCo6hVS/s6Xqc
ThCzwDzr47cUnI72lS0oSw+tiSAwAFw1QMo5rV/Fy53toY+iulTUf+cSK0g1xA/4
303Q+ezyIsa5e4Xvjxp7lq3iZrvz+rx1NOv3bHKOmtpMqqSAOWAM855vJ6PGc3mw
q5kWaRnxORddcpcTAXsI3WGLudloW5oO2qGAbSmwiCVXxGHWw+8IVzpuvtz/4Jz5
QZ32a7C3Op24jBG6JaOUA0coygDrRLhrS42MYO3AXgxXx2WElofhAELXAjbeviki
eU4wNyewhx+s7X8H3gAbcXa0wDAA76qajO8QwZ70yRL3HLKGL6j+I7LavRvDoDQx
nknhrsdHBWelHrCrFvqTo+8bCUIcjwOMwWV5sIYb+X63SWyU0PhmfbeAhD9Bkcos
f4gC+oY5L3v6+Gz8ZJSStG04xIcgiqUm51e9ATRxqKtVSZUcZIapOvboo64ShCi3
S3/I/ConppAhN0vqWXEIGVIb13OpZcxZIbGy2cv0HZPC8bgK79IpNWiaqLe6uV+L
9ltSz/1NVaA3kTsaqzuQ8oKGrGGE/pa932kJhpZw9oVvS3Hq+i8h64X6IoU0XT9u
sfc/DHQudaVy+FAbWAKjGMaX1crBpP8qHZtqPlermb9K+vMlLczgs8Ve5Y4NIUDp
pzEmqzuDWJjtZP9x+OaegSxBMavQ2mZXPKIeC1laOX98364YNBT6fGCzcXd9YW4Z
ToUVZeRRy9ustIxbvvrGrSkiKtJe7VWdKc50XOTG2KOkk8Qn8I/CTP6HsISj559j
FJ4ofK8AuxM2B4DXh1LTDHbYdMjGvW+XbusI4l4W/7TLV9foz9FspnijZyh5MPdc
Dwg3bIC410zOatuWgQXHvuvku/G8cJKopn4o41Y155CMKoa8bxV90RSenTTxt26M
JAeVKCbEX23fTHKxlQgTfYz1jeRTq1Ux4ooUTt7jT3tImtyxduK0cDVtyyVHPysv
eGZgPaR4zN4IvtZs7QXiav3rQrCHzfrTKzIMKGViwFkHNRqgJBtxETy7rwX6Kc9A
0tJ7S5D9o6QxlwoFvwwPf5UbCA6t8BSmKf4XH+KmoOLKr3Lvq3PhGDl5HyIx7F7s
HkydpGm1b69ouCkr7DUxR0qd71rplRH6Y+tfN39IDF/5ludBc9UmoUQXaXZKyAM4
rPzWay466qufler7Y59Vfch4oDX+5D07n2jsfqFau4cwJbtkZMC3HpvvxwWVuT8l
KVXne7p3f8dRFOJHKSZQuIg0m3UmfVZ6WXR/bAkbceWG6nFEwXtnpJYar1FjOAlw
uODgaVTmnkwk3yAeazFLRh4J/++bwYjnFJRdHsjCHmSIofp04LwDL9HJNMYRTWlR
a0Kd3Qaq0OK8D8M2Uk+EgIpyyh/lNOuXDw3iP57mO7+EtVyI55g2RfFvii8qdLuH
6D+ccERSj9goPlg//U+jxID8HUJz5eg8GneRRnOqOpUPK8YLBCAPyTWDQb9Hnitk
ahv1woljQ3eFc1DfBOXXkW99ufofjfm4hq2kDbwmaNxbfc/gPU37/1AjdRXDkRQD
WfoaNN5VlTyAQt8CsNS5KUjCNVK32OIWcIWC6P2yvHpYsVDbgXQI/G8Ug34KWyHl
qu9XCW4U61XNO5dXztDa+andioU2hApNwVNE0VXVqwbmQi+XvS0VkPpe3iyIW6LK
Fi4GdJlTRm/Wj6g0QtR06EPHuuROzvmIzwre9iggJ/m6RoaPCssQ2ZSzZWXyI8rU
nLBCroSexWLE2QMJ5nQyGkulBJbEzlNQQLD3kckYBreadWAqU51nseVheKuOBCmG
u7hozXSVx6ZHDg4qjdfW9Vd1wrUCjv9DKwFPKllRVP4lhAZJDBbasVvP1AKCgqUw
zgfcIdgELLjLgW/ZIuauHj9apqdpTjVHjfqGBuiB4eYoV/7aMTR6ah11fhwll+im
dDfvU1D0Fe1UmrmAR8QZw3hlk3yw3ERFMNpcVGph3WYQ7vidJqOvhBN0G2WY83x6
ULaHS0JMkGGITIPpjk12htM8pja2SquebNR+TfUHQMRwbSIJjY3va8AmZZKtPP2m
2J96w8NHhS/NmYw/tUTDMSJeyxBcZfAH6/L36aAH9dl8azhpxvOl0fFMaMu5a9Gp
MxAPZbNF7DI9hJnP0Wb5G4DypOZ0vneyVDleLyl+MCo4AYzW5lgJiKlfhWGC+Hv3
NxV5siRFvKT5EUOKWrWVhdHQ1Nrr5jKv8w2PdgSgs02RdMvV8H9g0IVhJi/b/5eW
Cz/KjM16kkX5isdEBEKmUVE2r0cziRFcT9R6YTJc2mmOD8BVCFmltO6YqCUk/4k8
j5wCcvkgpgKNDM0UqSpVIig0TrzAnt+aDGFc7AYTQjS7XXyVfciB3u1UKAOrA/BE
wl8JUgNrhiRDzPFH50IVHxzoenJ3c0z9RLSslV7o173UvXRpFiTpnrpb9xQ9n/Cu
OVvhwb8tFt/ek8S14fNlVqSnRkY64e09E/tTInWTcecwlAd/sVT1elaW3AaL4QGU
u57M1rseUACNalcOBjlKeiQw+m5se+b2c9ELc237bBVkYUoNKUeWRnjEaOwmuBw6
ShUya6A3OU+mcg4MH2Qo+aHVt6JrGSZxrKUJVDV2/TM0ZRy2m80+Rx9oT22/YHr2
cWyyW3KDP7aQhRESIIHOauyk1KBw1yikwM27iqEIn4gaUIyI8rWUVCKbFZzPnOG0
xcSSwbC+tCzKZdZz/Kok/vHitESOYy4akAYWouvg3kBHKLhvNHogjn3AALbpDSlw
kIe6JQuhpbNVMxSHoRmhMQKO+V34ThUE6B8lQaaJBm9A8QKXFpS3bYlMKuR5KwZG
mQDK6fX2tXQf1RTVJ27qaPjilbr8O2LeMh7v5Ju1A74EqOzjpcG0WBWTLpXVqMFU
yhGniM1OERVdN765hCMb5VPmbQG4id06U0nccJ9UwXPOdNatf5JuecMkk0gPXK1g
xzaWEF1hDcxlvDfhZTS4prm0R5502h2Gk5VhdVsg/eet9GmvEHvXHQh1gjuDwRAV
GyuWyVm1INIOc/WxCEnbSDJHr5qpVSvtYjJKN4GARPjZl2HPC1AkqyjZ/yCxxoIC
bgPACvDbk6QM3/6sr78XpwWZwHUxIGVuFYna6hEQ1/7Y86Fqmfo0SvCFs8aGVLPZ
LwO0NeX2+Okxd2ebtEN4XtUDmTDb2HgqZzjtMDLMi/PdmO8HSfpU7UlNLorVxTay
K7oZEm1MV6ohj2QJkmiqtTHki2M6XKLuidPtZGYqyb8/ugl/IqSIPQ4MNgJH+qDb
6kuya6HQ1VmTcuqW6o6dYcWDDFkMdQcirUZ8WL3/KZaWdQbPrjlDpOE9IIs2g6Tf
nhlUhtwF3IqGGk9F0TuuAZkpzLlYuZbULxvFwwQ+PGcDZSBst98Vv6mDzhDvMKeD
ckUkBbhoyt4KFT2NJ3h3hLxvcUKFdUGBnp3fGguvTulDxiC1v6nUJkzDsp+pwsC5
5rBrwAqJNdQljE4jU9sNZwZlPP6NYXVha097MI0S8pY2QCBId2owSZbK8gdLyGjV
bPCFOAhvCnmsHhWOsdPOrm45fmOBUSADaoPt+edTsvgVWOEvYjYvuydQX7Rt8uwe
A1DS66zUCV4XreuqtnRRncdAaEz86+IoIKrieS/nQX589YulyVTywdJt+8Il3dF3
jPCky9XTjViOZn2TzEblvIKol2o2Rf4nkZr6vbq941CRm/C8HOd1pK/ZU18RkvIy
rgRqM6zBRc5fSCoGGZU983xxXgiGHrDpL1yllgicosghmG0/DN9VNFJoaTXBlMGt
BrJYIM3E/ifW8pNAZHWR8SWDCcGW3/YSE4go3WBPRp+FqKNchfowyA9iP5Fq1CEg
SNELpFCkZF3aMd3abvLeDaC4KnVqLAozhBwYa8Mry8ck4h2n2jv5fs+ELlqxXHn6
p/Rzb17aLPKlwsHpyVEVi9VPETSHQtWOnoJP2WiZC+ljzOiXlW9WmtbpqHyq71Pf
uzRFW0IEM6Fh9qMPtgOQRcUALbrZ+gzs5sFl/pTeoSh4/hs9DooxCUJXiHV8zgmD
DdLjsjXHzj7/2sCaey5zWAdVl5cF/JmopsAcWlO/uEtGvzg6kD012DQDwotrSFd8
twidlmFw84ZPMKmQC+n1ydwooH1IteMkWIF+TuTVVqZKPinzZvYzw5geZXO+o2KE
/0FbktPm++3iVQbFBJA9vrHV+EDDHAXs+V+JZGNBLLx0SlQnwC+MZpZ3C/2H3Bin
P5K9Dr3ina7yEOUQC88VE1mJXKkEJ7NAxMaZAYVS8Sg+HNK99hDecbVCriySgkAF
ysHT3owghoAIbNRWwm9sXU+669eCnKWdCuYn5dlv02X3CNgge8D0hbY052OWosOy
IEuDeIZhnpnPQ5tP82ziiBjn0bOB8pHFZpmKcBHwgTdAt2DkhaSOeB5KZ7XWVUFW
2uwC/U0kkeZDctQhf/0B+D391TshTMVgUpcRoqT/wu7rb2kz3E5rfGfoqxcNiAbv
Dk69qKfHUEkcfjhqKwlHokbaPAood5mghaqqTo5B1YW00fL4ivYwEvoxToc9sbb/
6bksotv/STw89dHkaH34lRAIlcj6kpnxLJ6WSbYXJVd4o7Qx7htw2XDXOUhYktwV
4UUtDL0a8BxzeDLrGytN+fOcTFIv1P+bfe32dAIzF/1W6FwHDwXvwkwmRQEYc/Mi
2UPF7Ke9xjt12bH7Ngmg6TfPItpNczAEncBxIfpnoiLm5R11do4skHCZJ4TJFhSG
14m9Dc/VIDWVSe4hKOfE/AUibeMj5xhaJnQrf7ZvmbE2daU1UMOEbI/e7hvlJmiD
PaWCPqD0TdRCf8NFqJQwQ23LfaJjOb8xaBkv7kMVis+exzCgQiavCBq9YUMYPt8r
lZP+rfgz9s75NkDIi7EPmU8k5g25A1I0i6E5A8LazsY/UUTOo74v5485jbL8Mp6c
1YktL5G8qJUrNSgbYN6Caicix3GPV5dwj2ffUFP4SM8F4XdFogWrNj1x5jNt6u6G
X1D0QX+63gTpJmEsfTD1j1l8XnDaqypo6GUNZPmLIc/YQcGL9yUouzhIz2vYLAzX
pdglOvRxqPp2Xahgzq0XNd0MOszJXMyM8RuZV05iw7w0U72IOKPXDYUCH1Cb6Veh
lATh7/VLr3m4Cbc8cCasYZ/ZwngFW5pdGtZrVdwnYpv153/YIFqKzs815HxYppns
2klenOhJZxWqXEJaqTGldkzbjCsfT1RX6nmiD6Ig2FlubPX8TzIjgh1P99g7tbTl
10g0OnXx9udNyBB3BfaB8rSVEgoArvoi3J1zWa8XpNPdFsKqFmOigFM2eQdvvAZH
lN88QCv+Pla9lcx4l7iz1RNZ/vxBxxaIif0KCezVp3KqRlSQo/QI0pEwGPu3M7zO
mEl3IdW5NgsAx25b3I1FzK3ZzL7DpD8B+kXgU6ZI75n1h4Y8fFACLfX3OZqQqiXN
8QTWN/wxp8YiNCsOI6ej5Wu98C0zhF3dgEexn4kQI3Ox1abJT2PkBEFyJceUYrzG
0YxtdbZfaMfivSe6mFrN/6pP938WLxDrDvHy+81HbX7QRiKOzzHCCEByTxqv7K8M
xVgCiQxmGpT7ncioIiycKPVaJPfapCAvyI31KfXLQw54YYRCUODAf8ryApjXxvSR
AniIuKCWSz8uSxv6khPCzWrkWAga8JZpuGEiY5UuApcQCMoRcEXZnqdqyEgp8WAX
eyqGOR0aI369L0b4W53TEfGlnkbO2vbS/GB/BQFy78N50glL4SWtPtsg/1lrFs7E
CYKpNtzgh2LZIHeVr9EAz8/ngs6NEMqvvTtCi/jF61Yzw8n1uMMlRBBhs+Jmn6Rd
CXhH+92tOvd+QW1J6ibsAqXkO98dMWyTifhoKsX/J8IMVuICrZVzviuDx4FT1eqO
E13KITmbiw9Zc2IGeVDqRvQxmd5KJak7oqQ0MPiJtmMPA+Mi0vM9HFBQW+i0j/Wz
2E8Az6vCKlNzTITKZsiUZHiVmCrgoxrprbt/dTlXVucqjFjYGsHi5zdxQ2sAe0rT
/ugKBx66umvqFb9M7WSeWz+PLW2AUJrAeHb9w+xKPLYwJq+gRYAU6tGyy/t45bfZ
oiO9nBrZPvHB3xdUMaKf+iP17wS/aj9Rdi14REHPb8A4n2fpvMB2M18iMhRGR5UY
JSfmruamBGx1jThRfDOLIMX+7z77qv6nb01ok12JYZ9BTnImtyIU3y0Xui9Pv21u
zAExcllJaq97CbveK4cNPe0fO1rXOwcd/8hDP7YOugh8FKR6r+91bJ6+sG7SFn4c
XtoLevoKh5s9wmMfG4WIQSiz05RDUoi8ObmBcWmPVT9SGpL/vPpv0cJgEjPmWni4
EhlDuYbMR+/fzx6n8nMDte3Vjj6/2eq8htaiwqfSj/5x1gCic0W/8febnS0+wsVn
hX8ZysQPd6frdaX9VrcG4RyF9XF3sOQv6mRKczlDtpzkgkydJ/xKtUAYYbwwpQIS
RXNeLExymH/cdodJPUjAT7CbZLgsnujOadlCr+p7tvzciZxB11d5w72gbXQreYvd
3GqB5cUhuavRSuGPtnUHLW/b0JGEvqwD/UNoNkuewNOxhGcbhnTK4/9aqABJkOPJ
SDxN9QiDtQYqDe4ir36ykQajuFLsMQyYoGvKs13n0/L3ss619eWAedssNl+dea1u
LYpUL3uMLiGZMtRJZ+A9SJUwF6IGmC2c+Gm/3flcJ4VUmvVmrZMOoXQT3Q2CRJHV
86isLdxPxCne53JKRZkapmkKZILYByRRuVcRk6ItAFFsDBFHKqg2g7WgOEKAyfrz
wtUJLwoA4QY3onV4WBvYbNJPyWkIb8yqU8c8gL8McvV+JiYJkrj29+guaAWls436
8jOU0Mf3JHTDmTxQ9Ri43UiJvOPAP4DRWwKPFs4zPzy/ufl+Ct7z42pSJzxYVo+J
O745lpWXEEufANH0Y4FJ9SuJz2IMAb972XNTTn3ourlzUudqSvgqb2Q9jILgtwpt
VMRm/aUQPO3SmUSjSAMN8IlFWULTpdU8+CACZ28+XMrb8GiEb6zG4SZIlJeC2f0T
ZOsYN7iLQwk6TjsOfJTcThIdvK/7lj9j1ysLkFGJydahN8LY6nOeMkvaZjI8bMqQ
v9KMe7gQBGnkjPYE8lSq186ctTiYjGQP3b30YGr6JvtJ2zNGOWuOFBpzHPP/40Kl
nROsGB8zIxaMElcky1sbzBfcDEom5WmEE6DoqlVgncu3OhzHaRLA0FcLki6mFm1z
BWNtGUR8WVXR9tvDG7HBYKshOgd1dlxmszvBkjj0GznKhntYVDYg4wUdqrBKtwod
rD2WArl45JP1pD5jBRuqPOFF9udjyaMNBVHzgbOuqvd+slt1VghbQvZk3Q885IIV
dEYsimI8+Awx6swQYjARQCxp1ktTAU/b4BaaS7wGZE0x7u9avJtL1TSThpWoxpUB
uL8Y4fNJ58R1yR5zS8ZrMFSvi58qsXpTipIWDxCltzbTnjJhtDj99O+VvasY5BsQ
E05nbJh4QeFs8QB3ArawkwC0CubCkxtnxeVWZcCfDJlfRZl0cascfYSo6texA6l0
LHH8nAbUw8E96kZARfZFHFVgyTCwhOoQwG/Gw97xz7Zx/iTKUD4agG8AU6IsCYQA
xxqc95QsWTq8dfXC38DHVtvBl8FogWiBuhE11oaAKb1StPEzQIX6pM7AiTowpPoE
kxYyNd1H/A2OJ7U8SOABogKA04x21d5U3K/qL9pFYE1c+rU+pOtTy9GOf7eBFbQV
g/vxP8bq13SSvW9wLn2Xa6AkHjGGv8i7h1cyibzHL4CQU1XrIlo0JpRCIZVinC7X
/VGFwBW/7hsSMRYii35oJI7tv3I39T+5mW8J0ISRG9a0WRoBOWyW+lKoarnwS3Zi
UT/l9vLmvpDcFhgEscvJye6PKfoqrxI6S+zgu/QTCT7TS+gW3tqSIDcFZ7ZjYFsb
RQuWzn0etjFiqWe7TtSmVJuEot9tAoGhKQPlWKi3khRTeYJgzjjQRJRc2IoixAYq
virnYoIY5cEPUuVERt8bmFvQAf1HohrAfjcTQvzO28iQqOlrVmvGgtq3TFS6c6E1
4qXodkHTR0AHfSfE1A4xTMpsumzZ479uCFO+BBXo2rrnQEn0vH0f2WYuYvnKGPZy
byTR41cuEv7cva1cfRsUnvOPz69ZjiPWj/+g6sEVA0KV4v+a2cJ5/JqOLhCNV1OF
tt4jUZ/o5qGKLy1TYSL4OKgeQbJiMFxMEeJVnTmoHXH/4S5XZZu00za5oK8QQjWT
xpj4itQn4U75uj8F0I0ZdH4YAdcYUw9v0F6mr591F8QhtkvMWNk0TX7/7210xyEq
2EBGlpL+ACKIPNE8UUNVmo9vK46UoBM6Z4IxiD4ia3AzSE5SKRqXmpk9OQFO5aXz
GAn0T6+BdOfmmrHJ8vL52db3VGO9y1411LB2oMjWQ6kGXtCThmgBwT6Wh1M4fej7
v8+9mvEQdiFSqAt8Xjzr1b8bGiOhg/c2eNOAa5ryfg8HSCom0It81KF+fR3zkQMC
9w6lesuDOruqHjw0qlYX6l15smSywhXGXwMn1ux9jGWc3dJX9Q7IWRkVuy8Lsp4H
VPhvIH/Su9oFKmsbSN+6G/cCE7wg65mCkPaCL+RwXMCua1ujc38ZwhFVv9CPseIF
o8V+a7RhDEmxeEXpwStk+5GBmTVFebC+Ryi0F1cTCs3lhl67LZvz10qq8c/BARTQ
8V9SVOoaFXzVBz4OSqRG7AIHGA6dACUeRQh3Xgd+VZgtd/XoX2mkCy1B9ljjrfce
9jMBlCM8cRFIr+FrpxUGeIoJMgWtii6V8lYjnaTgJn6XnoU8q8JpVG0bbv9KzKBk
VwZcWPdFN4EeXlzyDqqStJmO4cY6hHHXH/CoFf409vnP29l475P6JH1YG3sEQh40
LLtENy45b+lKiFcHvAsWXAVao3/0Zan0xMCESX+I5vD8EiXofsGIJOMRILXYF29+
Vi6JjCzjboZnM5sfe2sz3PIiGzdedZAip0LmQQ4uvMQ9jFKbQ0kV+ZLpraBKQz2J
5wb7B086K9HtJVJsk3W3jHSjNIjoGe+db9EEruOyZ0hsCHkQHYCLobUqce4YpAnM
GOHx60iWCkSn84qh61ME0i2Oksgg/vQ8KlEtFLFGI+918PaM4T9jC9onL/7kMrNh
R+copkzbt+h474c2zCWc3UajmXCLVpNAageQ0GcBH5IVcDyRNKRmdacg2ufm7jPo
cM3vW+uYOHfNNnbis2mRkSsJTEirBnIKDr19paK5F4Cjbu/kvBLj0AH3WJmF6Y1Y
Lb8ju83OMivlQVASPTsANaRaTPsflNWxeEho7xcg4Zfzes24n6fdf1aix+v2gcou
OffXvic3VACtQoMCB8vIVeNuFWH7sBoQAT7ve4qKHu/Ljd/rVIEVzQ8UviEmvY4R
Vpkh0TC/QgGjgWVFIjFOGkpEfCdz33UKc0JcwBB2pl7rPmE7d4tAOZPP8iElVY74
lUCoMbrzGKf16CkFwvXGOiTlzTK9ycQz7hw2HhDCh/zvgo20opJCUbd73lS/DLOo
4FJzaU4ZELrVE9xCitaaa4OetkMxxkQPhACUzOray59FJgQx5cTs1u/p1jL3+kq2
x+3uQeLw07Ec8Thhk6fRzfUHDvujjsXcN1bR8oOGUq33rNxPzCse4jcGoeUXf1e4
rVVlwHCaUtMG2/+NmNVt4SGXGwYK+u8d34n0NfspnPWn3qt+bhsK/lM+ad/rVTYx
zIpyq6wdgcVvkUzarjeWgy5F0v9eDlkWRCpa5lGpXVF3isRYYsIwmvQ5S3Aa44Rv
8mOy35XgInco7DajbumA0h6atR2zrSk1vSyPYJ1XYxfkd4rJVM2HQJ5DLmFHVS1M
2XTaOJtepsE2zNxazG7TQn/KXwc9hEdRYDJ0e/oQNHFw4rb7OzwpGfeHr4UuPmFH
9h/awsdRuEUwkUF3HUsZyQXkonnkInxYh8uXJxcbRbQti3dm67TQNPfYB7HOJqrN
RI3L4ghWCqTcU94XC/8chpCByOa4CLqOywzOZMEcWafweTEQohHEKPxEBt9uMcvx
L8N5WlJ8ftLm7iDSdRDLaPEcsh/mmLglQjHwup8Ycii2LpmqSqDUfWLHEWXEvEXD
6Htl6UZYGbf7uUkJU+LwZIFA0CNzcrFfabIpt0P0mDMv7XkhYzxHIetWU9knOQM1
rlh3YbkMXGvfNMtm8I662wSorOq8qVlL6NUs8IMa2G2kWCuLQOk1TbjVdZGOK/GD
cptnbBQhQ4eGdmN5KweyOXHLOxFQ1ZxB6fp1L+LG1ZNMKr3xjFK+OlOH3qPJtKje
Yw1pfwmD5ej8+fCcF5Oy9FyDI8okMV7iCqpg8L+xlaSEYNm7hLblb7R3UDSO/xjx
ZL6dZZ7ZEQqX2cTNpbrLO3MK+J4ue8uE0tMpxAM+Nrre/GsXO0VNTATzYkxxrEun
wkdkyO0nFu+Xx7omLhoeee/QtQKMR6Dw8bOb4/mIg3lLcD/kZNYXP1YgdG1IVnmm
X8yHSIEgPXDIUfi6fqXrtnYWSEsjpYaCVllAgf+n8zQ4LKyNLH6t27iUhySWew2O
kjKD3aJmeX/Mm5VQXKIAzjE59e7yu7SVtTn4tspi5j3rk7+hEniF3m5+huRj5Ltc
o06y0GtL5fJpHrSVFI7Cm1KhWkqtcMZ4l4gsD2dUiEKnjNR7ybrrfPx4o7b2nDtz
GRYoZQRZazj8ZTYoAqw/U3jXOL+nY5ngNmeZiY+aSJi3QOe5nUBIvxPao8PcTc4u
Xxf8TT9immCTB6mMcpAIctEsC0b71gZnTPTE896f4KwkX8VWZiWKM8mrD5a890Dm
2v2UIh0saYVtVh76ICd7B1CGrcvq0nQyzBX4Il0WqzUn0vo6PqxqqPcCQRXWX/bI
0i220x09axZUTr2EcR9CB16Ek5PV2MD19WL6/BSeaBJn+T1ppmcpDdj5rFQ6K9w3
qvpZDOur/0PmPx+HXyyA6VfwCgGspho9AyCmfGNJSoUBkRZeUczzuuNCjs+dxqPY
EpvhxP94Ph4mevlI2wCE60inXz3Qkoxq6a9aOgXNc+2flLjMZL8fF73KI18w/6Xa
fEm8P6Q8QrYg/53eg0fJ1NP/diHYR4kI33XKNFLmiOCsvx5jQ9wZzvVsELqblQxK
dvkWnSMwsO9IHxWRwmWbA6vxlyPiirciU6AuYdC0dT+ve+S+Wu6/OFWxxPR+hauO
ZUOtQRALbQnsyIs0O0RRJw14Kx5l3SceL6Yq1+Ysi5zITQpFWOIgfRZmZE9gMpqH
ycr5ySo0EDra2VCoTrXIYgWrxFGzKdWbIUyuieiPDlbqQdZa2jUEdvYlypjSiWUt
ASoiOygkMfuy/tDI9McrpqQo+kZ+WVwDvYtciTnQDEdXBIG5ooOYWc6j8ZG7Q3gJ
pGjFKEWyZnFsqY6OVfOagEp97xudHAGD1HibUlLUsyZ46h9+TIGJYzNycM1uMZaM
ZP+1tUo2i2fAF/wp2r+9izMYzE7Q1wch8GZrhQMpQCndHsutWkIc7UZ5/XM1XIaX
pJvBpgS1fSpdLkjpHugYzKvd22hCYSWtFDmivh2YSAwRadq3XQkZVlGrPjLLw8qw
Ht8D6wdASCpw6iBrnStukjBVzdsMU7e2TiqTQoLS1g/KYvy9mcEiZVM418lnSPbt
2OUUAzLHZCImQA2ROmfCjkMy8T/N12aeyQFwtrF1g50H2xVgvXQwyw7hESzsWA5Z
sPnQ4ThWkpwVD8me5d2TGer+r8jqvTefeuWSwryLAAto0zbcl/3S4nP8ks/E8uim
jK1EGmE9JoiZNV3ANkpOJglr52OPpesQ1GWCKk7OusiEXPbLmQvgVin9sC9g8Mj0
K2X+B7ry/iqg6kGT1M9rNf3RHNP9OntxBqP14o2/ZeavApP9RqBgvC+iapX+z58/
lskjADZbcpmllXkau+P52cR1jDwaZthW02RoxpTso1xtjDjrULW7n/dUwlL04aku
2YdAR5kSnsCkWCbMbKSyKu8nx7DLmrV9gEN98pGZcP4LC6WtH5eMuV/GtKUZaS5p
mmrBKmXryiXCCm29kmlwcKYK4JH9wgDHuhdmpRYLXFb9qZTwtj9NdXTNgKGdvQvI
I2C/8Sm6e4nZIdtelrCxg+XzsSB/hHBqzD+6jJ6yhW+1eSiaaNMlgvcj9ltw9Hds
Uxrf7/EFB3ztUJ0MzjjKheSp/xc7Rhn8NrisFrZ4E/hREkHf/Oio/VN3Td1JzEkQ
FPxX2gz+H2lotBjCdXVbKe9fQoW+Vt2yLa0hFIIUFPIAdPmpDXnFuksKMoNO2xdq
yICF4V79MF+qeyvjVhdrA9N126x8UnSSk3QOJn/griMteZFJB/vnOxhxYBIqcuKy
qa3VOMRG/7n9ZmMO1t/CYVbQaWuh8GQpSEdFicNV0Qi6v0Adu+Jx5LZbYLVu6YGv
hrVGrZYWksj/Yhv40PpvEP7ttNPW3NaULiK1aM2hdbLD9TIgZaQWV6ai9O69/ekI
rh27sTzCgqzoeQYoCZTqb90LZCJNioBdeAuKR8PkaV5k5u46hV1ys5zvT30eO2oF
e20re4UBJWREnaRTwbHtmUFGhGRGR9fDhIrfTIaCoEbtqvpuDRlELcwsFrvA1YWe
T95BjJr7/eWv8b7uydqHBnmxA739xB6/yFdDkO1yXiCvNNp1iuR0vREwzZov2eMi
g73nbpP4GOf4aFFOWcSRN5Fl2DhfIUTM0AUePVSF+V1ZOOoj+YXVoMseJonnOf9s
5Up1mdCy8fi36KVjBDHFZLhaKf0/3TehG7TT/TFYB+Kd635xai+rxqWZ3qTIJ+IJ
w0PLKxp/AMFiokgDp2G6jQNxMJuq3PVkdBBiq2y6pERYWexmJXgkLDq5y2Wnmpp5
puyuxuAW4n3262RHJDoUB081emJQ2EN4E0Frzs3w1tAEcM2Fl4osDU+Rd6XEynUc
ICB9sQkJIpX+XxTGyBLEC2NvJJDZC6UKw1khWPGCctnn07/TADXzYi+57atS2bD9
QxLtCETrEs9+EAu/tNwmEaPR4ELcmuPVdTdLSzMWGBYS1ZejUToSlYI0/TbubTIj
3zYP88SywaucNoVGb0E94tkk1EGJ45cuJzkKFhf/BWoHFX3eabFyN8DZb2IDTloW
2al+6S6zPyitTMU6q4CCGFGCBwBF4iEo5jWG2ztlmhA454vO605RQYpPZxGHt3NU
hIgLcQxnXLNgeYPCXKekVs/B19iOrHJkrKJNNGtWGINtuTCOZSDGWoE7B29mOmPM
3/RyuYXFdKNHztR75OER0XXVXlUHQ6EvrP1eQbEtXOy1ev8eKySplOKWW5PDQdVx
my2MucjVUetZTEYGnXgl0FbPiQiEWZ5kKvjLpMfTICdVLTXDNQNCnW8v5Wp0nGx4
PjnIkmdVe802QrpujfxGs0nKtYBEAOwjwxX/m0tk8SDpPL45Lt50RqIVI40KFolO
9DOKvdcTSisPZ7DKze16Z4DgQ2ec2V2pRqzrfL6UKsF4scibLIv02sQxxtyVe3S0
IXThE0mXS6ocU4Xhk4FWdG7mYx2Ft3XNS63vUAFekZyTs5sf8PRwnkewyZNr5W2u
QYXyh6BB/lnBPB/0eNX4xzpV97bhfeDupKxgoaE3eIAld42k+I5KHm/AXWb+GKO3
3pjkhh8RI4FUVBr0M74I62iIElv5wPbBhqZdPtp8B7Gpedcj8ooJoFKVFcEDooti
DYS0U36TONARd/ghTlZHYcBMhk+BXEcITNlB8ia2pwWIFWl/e8QJ+EIrhxXnh5cI
sBHaDjd55X2FEx0EvV82Yvcxw10/upAhGb3oE9rR3lHwXMdhzjN8JcU9bj25Tp6q
qU7LMWd9dxOJA7naK0CJtoGx20F5S5+7J0Yt8BhWasTW1wAn9LLN39y6NgfBtwt6
dFsm/gAyGp2AP/F9vzJbP8RZ2fj9Bjy1H2J0CUWy9BhFAlmnNKioKRjLfKv2Rcfm
+mxxFCwRaMZ2L8wZK8Cr04rauDl7+rJxdofip/Ucg8QUOtgQZ68vlUG/if76pEqJ
aPJCcs/KyfLi3lrpgt5Lo07XOVjszoTjFpzdgWozmQ/zXLn0So6vpzdhNQe3F+w5
vuRomw8EwJBfBEFXv4AzsFs5lpyg8rXj8w704vebCwUR56YB5iwcZvhfCiuKEOPP
63FhdImM9RUshMQrvjeJu3zlN2KlznUchSBn199Jxk4zS5BPcEEDET7l59/ZDv6i
vBMZrkIs+S1hQHUz7SrgDVmVF0APciA0AsJSMbk84qQ=
`protect END_PROTECTED
