`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMY0mcfeTUydGN6bm1Uum85+Bh+nhaXtgWQ0/KcmNmyZv6dbEoI1F52Az1Sl/kIh
PXDng54wT3SDAVzq4QIFOrrgVX7bgErM+hBRAYTvJQYsyTwLMt23EZLp8VJGKdfM
6q4PzwsvAVKTthgkkxqcmLBL3CA+31ALYVUUd0i2I0F0ETIFjsrXQ2Cbsi/CuLJ2
+BiazAQyOWZnuAsMC4cwx9OdbXMZDwhTl/TeuB/He9ICVjd/0bEPGkdS+0Q6o8Ex
Damu1+/PydKJBSzBx6W9CbUNu9wr2jYx90cYW13IVGjPGVpwLrQ5qNcCq38db+6j
KRBGOmPb7191XwyE3p/1gAKfmIGAV/wKwV48SNSjYi78B2eYsJ/Ul8VbNeqyOx7T
f/+cRFQIjFf0cBw4VwWka9pL/78ox4LWZrKpDS8ekw17KqKMmoVddxfK8eyBUNij
ZqT8eW+B571Y0YDFIeCVmDB0iiTeHAHA0f8cBQR0XKuRRW/99NzDVm1I1GX299wH
mSq6a7Ka9PkxEbch5FpaPZFk2KnNQ1eG0EDQMo0sDthnDqD6h54HhwNLM/yrY1bF
RixjRYH8pJT+PBj2G1nNjq8LtSj4knN6Vryz9fa3Fl1PxCsjz9SPlPWo/frlsw65
8rDohcd255oFWOZf68CwFLwEIsduHOachCuGHJ/Jceu83zFSYetoK3aRXyAqYZmh
V8vzZuTJd5s9a3DSfR5/aZIfQXLpolTScr9NneGSMtY2gyZN6vKSXSCDea9Gs5w3
4X5F3MsY41SNlq088HJu/bz6NghBnHbAVis8C4cDU4Z5P1ZPAPRxQYCJcVPkxllT
R+BwMJfSv2icspl9oodlIbmyaA3Pas2d1u4XUz+BtdpL1C14OmT9xHQrssu7vwix
hBr48Huk2TCj4FHkxWnibFwwn5CkBoK5JoDVHfOg/wMJhEtgSyihvSe9ZBZW7t9C
86mUZHwCuTvllIyHsVGKmS8gt90HpaEifOfZUzFA8ZXMLxL4BlE37ndon/uc20Rc
+NQWEIFQntrqw1/6ejt4K+GfovKWc5xWXtOVM2yrzidHyY8KNRYkbxH8hra5Nxop
eeupWjmjDpz7s0muEThRh+X9drHiQuG8UNBVyCpnRPAvBiLlB9068xhaYc2wiBRh
uj+59/4FZsV7nOh6DMIZeKJDT4SrXPJRj+W2hADru8ABJbl0zgJmYaVk7QuMqrg6
j82yBQer3q+DTEkmbLzHSCIP+E+6wsliwjiV/WDlX424ml5Mbezi+3p9Vu3NPXbm
O+qOwxyHouB+PZqItuwfl3UNoRGyP4BnF/FXz0/fpUScGerSY5VKeDtnWRULi3VJ
1s9HKt62bZnHKnftfgk0AHc0vDruTIOwDnVoei+pMB6Be+TAcBrHIloyZMIl4LjM
C/ChvLEtg8uPC9sN1knaGxmTKDxaAQecbfLdB//u9y42ZWz7oSmqy4RFw5f2ze1Y
2ZHNZ/+WjlOxKe4wrb+Z1lu6/nbPnj/k4Emq4W7nS72OvTtQslSCzaTVADp/3t7q
6Dvy4EHsyZERIUcuJdsfI3SG5lTLiuqvp3jpm2U8TmPWiZLA1JcglHGkq55eJYM8
hdpRLodEImdm80XEPDAyQeq3r02xnBvxoYSOWBQsnhzkRwtgu2ol+MoVmBemuI/s
sbysXLbv+D7+fAycKxgBnGJwGHXx0mphtXaNvpzpWrnZp2yFiw9t5SoqqVyUwA0m
1YqnLg30RJVf+nqeQwdDYAucokPTj4Z3uWlk2XYRaxoa0/epLfu+7uABWjigSdB+
VgjdV+6Yz1rMxX4uDblVRV+ZGqhWx7/V//2QdkB6TR/WIRcwX2yG5QbURPar2v2q
2JPXoRymXCvRv7FIIs29IH3/VQd11lCv+h3CqVDzM5nyroFKFYXOwL8SbOv+s/+k
NJS6FF8wcUxE9ATZKsYEel2u2tlWqvavK8Szv6K0mxwgACUcwOgv3FKDK6yGjXzO
lD20qumFTINYiK2s67VWDcL34hd476SN756XJ2NAIKO1ppKynAowpR/gcFMydrp2
vw6gg8pNMtk5YJqOGUWcI8EwRW8qwByfmY7wDfeTHHoDizsBZr+N74onVlnyOW+E
DuRZDe5MvPv9TYZ8ACp3JJ9rGDNLtMD/sinqbeHB4lokEQH/Li/1IwOfa9HhAoEs
r5UIY2Dl1DR+Hpezxg9Sonf21lXAHAPEgwxjpDzu3yPymDfYk0MhtRV29BEo7jHn
26t2iC5XK4wU2hoKXrD4iKkCUbcqrqLGbVcFUmN2GTi27s7+fKdpvfwZL1Vj72GI
Yg8m8pP3bn1YNTOt8ELgkzToK+jffNvg89Od90ZdxER9oXuen9SwSSnAHwHkiTzN
UCqqbwcFNH7tOJSYxrPvaflYlXAp8qKaRQbsBQ/nYw4MM/RafxhscAKyQn89oTDX
BIHhcjafMTXnpSzi6vOMyNOxatREruQpgEngYnWHo+wxJkYqX4nU453faJieQDn2
83RODunNDjm7axzrONtQlghTLGPoZIAO08Rnoi7WSwx5JM/f76FKJUhbthIWHyhv
7VeZHHHH6ovOQFisfprEh5U/HfKFeyTSOBwswYQWTKoyYcIeDmuOFFtxGvJynRDl
pJ7F4ar/vEJUgbnOs6WzTb43r/JYaz++v02Cz9cQ/HMdeZ97THikkQn4Ums/5sBj
a7IjzKFLrn/SnuRHofOxoHjZX3hZkdVyPrNDU7JGFI7PU6JEj/KzeAnl4QPb0KdI
7nD8M+VoSfHiFkKljZnxumVIXUqCegESxMoP/25MvJchLierj1MIPuNoIyRKAhxZ
/8/N/9cmODZ/TXhRmzgi7nLlebGX1dOz19xOUn3KHnjShZxYxlFiRX/t88HmqWsK
9+/XhzMQ+Bc5zbE3P7+YJsy+4Rd0Jb37B/pYsAqoGAs816SRn8N2hlY8S2jIRk9T
BPDPvc0RU8mTxrVXVUW2eG5tvROJED+tN2xWRPuyPMmnBxIqnSZhm2Mo1DOuHiYl
KZULwf5aOaQCXNB/dTdIQ8/ZVJrYfY7niDt8UgFSHwyGGWDRU+i0Iw6cZcjZJBY+
6IDs7SuIVtlRxvGvTCpASAHTVCEkb72bZdPJN/Hd2X1rLWi437NjxwL8/43HGpZx
ZT6tVHOFgYFwY3oKh3xcS+tRKzs8I4Coq7+wX+xbwRmfDBbWSH5RWQb04dG8rtWb
JWq7EBgtgBLXz6EzpKmUUXQY2dg14UMRYbdldmkhdIVGhkYhNh3Av0XIBHMvfCPi
cEPvkBnxeT3lDrOQNANlhJzpYj+YTe8qhjYjnJDrvIC6273NXQrncunVHSoQgE8m
NB8eLoOsMnZlDl/bDuZUKSIigJWnxDHZfk8qQICjAhTqI+u8zxoM3ZDm3cz8435f
FBt3RM9eu6B25KIZM2OFpz9PhxgpOTaNk09HnDD1/R+ejmF4bpJ8r7PZujAAadM9
h1JwwyG4rrI3ZQQgbWdhrovYKMXGoyZ6emouCjruyp/0B5vNx9hAXVp7FWg5oZLu
7yblV+Er9PzSOAQk52WZeZin33dlCAeYzGCYopPrtqLdMpli6BBes4VdCAUhwzZD
GWg5msyVIJkNZZ/DMGj87M760xFmZA/T1QpSnrn6w/W8rekYuycszzrDjmW08ein
Na7rnZ/ZejmvBEANBt9+2FA0xs9OsIkMRirWjaUp/K4IxkxExmxaAnYHfpVnjBDq
eXNp8RvSbZoImV+QmyBzamt5rhzG/njoSnBVkoCd1i1E5PCNkJGA2nbas/f3diIW
738b/xJZYFVn86IP4Hg2WdKhPdHUwFkAcp0GDaI4fwHgajVowR/KxcFUeQm7G318
Mi2UjiDbhbhhZmxhFT2EPjac0c15HKASpoSst4svmjZwt9MCt1SEHKkgHhHl9nl1
unrv/DqQkdf+23CKqkltOBMum1E4lJcc+7pHzkfiTyrMQ8p71wlAHZoqDHA8ACA3
LEr++IDJLq3SAHh72dRx5Na8UN/tC3IY0i/wllT5L187J9jPMwfonWR/7okl6R1k
P7XViFaVrUEECFXWRbsyQjJChiSCL1QqbZo7LXKpT7s+gqrIERE7yGGJLJokWcok
M+ZQrkf5V6oe/YxO0oQC/KzZ+83PevcFiKSfrb3gse4Xb5ILKvE08a6Gk9wavIEq
iQTn2Ls673/IlmnjtXXxlDVyJ1PRatUXhlXknlQlB2RY8Bo/q8GXzDWEu2do1I2N
39oUBtjstwdvqqhy8ZLUKsRQ19N4QTj7DuJzbNtotGZECF3zp4BCjJdd52qJBsDS
t5Y7+JG48stNtj7pjF+tluuela5Twn1WNiM/1USd9VAYfPjxJfqyZLUnxeUdU/Iy
2Asm5s0i1YiwyBEtP2OOegjTy5KGVNGHR6QJYfSTbY4=
`protect END_PROTECTED
