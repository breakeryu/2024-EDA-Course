`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgGtIhqbGlBn5fHlaOip/TNDbMSp6hrTz2MpKGE7T4M3yW8B9+cf1VR0CGPWn67i
DBf4WK1jBB1kNwD6Mwh/kIRHwbuHfvL2HIHvqlZdkkcqTd0IG/q/rpeUOT7Stocy
kus2kKNGcnB7U/dF3DUAEAaugkIaEiEWHcLw+DvktHHLH6xqSffow/Gh2hn9acAb
QiBCdUZy1d0bsonUnU07bBeRkgBxJEqmAPcQl7D6Mfe57RUNfxk0Lwdyz/W90E4v
FfHrQfPlMlITlkI3PUN/elt7G+RuLbIrOu15E3U6b51BfiKcRPh11ggOj5OQKpZl
iCJJHx1eR9ojhSEjpX59qYYBmKzIGLHERbI9JJybZizNxpSvm9NcHkQDV1sVoW+U
YKxocZHCtHJFXuufs8bcDlu3bxz3Np0PgSy3kTXxtWY=
`protect END_PROTECTED
