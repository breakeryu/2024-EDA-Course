`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6zwoUwGYB4OCRlZWuHzY35Zdm+JHVegx2WxKEz7K6fxa6nIWIwsuWHW1C1ciR3j
AjmmzZqpbYrncD7gazCQTT8MvJUQOsW02u5ZH0Uq9h59R5ATzIp2EbWZ8llcXBbb
1NSaVQ5MpXEy5m42ysSvFsz5vQgLMnllBfHd7pHGl7T+jOKopmNhtx+UQuJlgGMB
1bDwjhdqO1gJFArFWG6Sen+pruqpOQ4v9L2CJprM6sq0n2QFId/LNzF2wiFDAfuV
y0NbrUGUb2RLvNLPetv2zpey9rhZ85YurQU4cojto9ELWQGR3M+6skzQmGgZ3BjC
H+E6IQ6E5si+cVRj90KivOJhFTxEcqMHvlopl5NbYepwBC/dRTQHyAplpkSgrS13
yKR6+ThJ3xk4h7DMYzJfvz13NAiSCkte8/Wn0HPk2X4VwFA7w8m8OYGlJdbLkvvx
PxGJyjYZ9NkqlNOrs+P0RvvlQ50yPeWAFtKUdEPyGk08HcG/epBoymvzKzscNeVO
klDhYBWnFvl4RaKbyutLvc8y4xtXDwRWKi2t7gtehseS2N7L4SSA0f42sivRRuqQ
a3qadsUoxpg1c+AwLTdIFnlVO1kLiqV3SzUDHnmwxHAOC3oto3rn8SAFgGCoJkG6
2XG+eu1pBgmWgPKs2v4gNRul4IdRWBuFGCGC71NUz6kvQWKkF+a9J9l8FlVcR/lW
t+3u9unYPvIJSI7E8yF1/KjLGHL45afVDmyBwntM39rphpG7jQKMTzOu6Rf6z5IM
+gtuuxX1eXdnv5nn7PoziGMnGhjFCAPizznldqLwFcYz1I3/+Bd3a5MVbpo0dkpu
jGYhJpR/A7YJA/PMCi2CdJRdqbPW/wT3+UV1AZGK+scUFe00zRstkXG/tZFH+6g9
9wgtyYsuq5uTNVTFWGeG4bbvrlsNHQ7op93agd4a0hiWV2q8QZbokdg83vjpDM0/
xMk6//TeHPdCizxwKYRts663VIEv9eV2TgulsHU9ocosPHXd09I7O0fvZkA+6x7X
0F5nQZzBiaJaGJAs0eF5tHDbfWvlrJ1HFx0De1SyLSg+ejL3a6gDKdlh394YzBDO
5k9ux9unTnLNgUKuNC3m6HSARGmw085jSAMwvBSsg5M8ECaO7LBSlQ5J4jMUbEp3
Z5QPAM/W4hT7dE/ITEsnSxDNgUR+jl+2z4jBEV9w5q2cGFgttNTgOQZi4e4GXs8i
D0fXsP/NXEn15Ug+3p9qfKV8csC7Y5c2B2LkxdrF+cwZeJ9WMsVBZKRJnutm2D/I
MzL3rkhqRW+DcFNReGurGGvk85+XproU7us0kzGZKllRlzve3nWt/PIX1RIO2Y/y
Kx8MY4R2qXCrZZ9sVCzqpe0JC7gXWxSCKwD0TC12h2CxYOD5ucPgocl2xKy3WXAS
6OxupG5VhyzRoEuE7JHDZ8Uno10Jv4z8Gln4az9ipLwi+rMzZWVrH0hPwkS3aXtN
6fpdUgpcwlbMytU2BseXul/Oy3ETJlQtHqI9Y2UcDijiDQxxlqRvgQWInhODiDEv
by0jIOSk3yhwxZ83/shigy8WxosVoiWh0NSNMo+8oFGgh+3eWLOY43W1pY5Af0Iw
DTr8JiVAXGkgVLO8WsN/ADFyzP5hVzlwqXuhsoMd2us=
`protect END_PROTECTED
