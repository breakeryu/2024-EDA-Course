`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Os5SLla41gH7stiyw2LaTcHgyMoAd9MhdOBaMAaDPseLYJsFZ7nTIvyfd4e++BG2
T6prGrmLd0r2iFhKAZA09szkbLEbJtxdLI6pnQkwcWMYrERSfCR2l2bjKH1WMZn+
xemrkQWRprOj5E904ENIY7PV4jP22SYZy9+PAeuH6n1DcbqqSF2zg9eaYhhD9YxB
4bEhCmiaWSvl/IytdvzYZFyFDjIcKp2Y/PFw6ubD5ihrcjZ0ryhjwK//exiq78fu
pS9FaVzlEC3GrsCsUlf8JiziwMPR/60tHcze1yqPXdydKI0nRWgMDCACWiHeEd55
9hXH3+jK5SN0xGLe8nPGNzFl/vdTDq+0h4zlE976rOSfjtpcIcdgLNVBBOxu/8Eq
Inn98RRirSHOio+mML8f+C83gT+kPDSjjr4mKhJPtXs7GwOPzA5HShYOV9jGNhNw
7QE5rbVNRUzMOh/IjHtPK+VsbdgGTfKp+8XR/ibu1+syJ+K8P3M6XRQeEAdkQcoN
BDrMicNFbnEzJg/OjAaMPGK3i0F82RRScA1vfdJBtf9Sy5iyCNzebnYNxbKv94U+
SGqnBBtXyibf12ZilNDVWZpsLMZC2v/S8n+yViafRWFgxNYhdrllLIRkpW3hHvls
G/q8uzpbvKcVhX++uF5cSiJt4iDmWzwjoHJ01EWC9sBOc4ssx9577C4M9ZMsKf8e
IERVndWLysUDKrrQwK4nCDMsa7XZUw5DdfNcR6s/KU/3ZTymtdZjePMzgqycTvkL
m388XgQ+HIXGMaGoVpCoXW+w8HmYNJ6mUzDfYor7kMDUZbn+Cgah4QxQTKdwiZRX
QIn/nq90YYV4ZBa1pVsG2KoCvCHbCu/kEuJmws25ANnvFsO+6yPXJJmqp9xUDeKr
CzsqXqgBUSj95hk2UIDqGdbbrT1AChKOKWkdFeWPukbFYEvnbXbropJTcbDeF4ZY
FD9S9OnK4oacnKuZFHSFN68XBtoMGcUG+Y9YekOqaoVqXvBDs39LntMNoV25sZyD
zaeuQkFxfNQz/Z3a0yM2acO7iL/jb+5sr6uFqS5SfizcGnthKoSt2RdzoAPxRQQx
8aganJjADtzq4hXg960uWobgpJqhWEj5brYEcGaBjxOVsyQFGVosaX4q6yCAnip5
xuIMD/TNRukh8t2H5sR26QrowEaiRXvuPx608cMQQCq6xiWR7TrpZDqECXdrfHKJ
4Kf20+yN14zF2xc04pR1lyZYnAjgzkexbj8oi+w3ZZqeiv0AEJYAtWtAMEQTrQyr
jUWDjTiQp7f4Arrh2xu1X8AjivkCQSOASNKQJT332aYwEUgN33GipsXoMsH9xE4Q
Zv0JymgvDIAMOa6i9hKB4vE+GWyxR3cNJU8khS2kEF5ir/pmPiCekE8WQYePlUHG
i9sMfWPmLJaLHeneJZCuPkXcVzR60ZE0ntkzxX4IsA62eAsyb19BFhWTGab4OhJA
`protect END_PROTECTED
