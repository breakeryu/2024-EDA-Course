`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2CARmrwDqj+FH4N5iHvNfXb5qkUmRS/eWIHUuT9qs4tBRgK1Ga8a6Jurute0uGe
Y+QNLAksj8AwqbhlT4LGV2k/Ebgm/xIUgM5BNKQsxuicEUd4n0kd7v7FZmJ3G1Ma
TslC8ijED3xYdJ8fK5JLQiPaMvMUmFFNWu68yV/47qss+tJOOrxTYUy0Bk2FIYDy
2M5kpC+K+39iEJ2CHMEmaXlujOkd4oIjCGfHeQOy5pS1enRJEAiIqR+C78PyP6Fo
vPKZe9MjXyFtOvN5hnZvFHwNZEQh/h3cXndgTOoAr8YtSZPnSLIifx7eVISOzyzu
ZlCFWzdDa59DVbsorI35xRLz0iNjpVfF4I5h64ol2PYFZwAn+D4NwrYMifAcz2wU
jVDNlwsTcOTBy2qmkhLr1dl17Z6NbjgkRMVij/4cZd2Ux6aNtMXR5TpBQkOGGtIP
h5rFZR+OZflW4W3aeZZncO25NRvuySUnODnUysZIUfu/3m4bViFvWkVZVv/RNWAl
8ctEYECF+5P7jKy9c2TfWDWnxzYTcBIY5Gg9ntoUYnjTNtPj2CU7+9rfuPoRwj/Y
7rtyJ78+VB2/hiG/Eb1x9KnHjbGfTZtP2czx+3kSU68XaLdQnKP7T4TmVdsdQ7FK
8T5bqpFB+Cj7tUdthi8zLdXhRXf13m3zIaNuSlOPL2HlTEbbw/7mV/VlV19cvKIE
Y/KjwRkGqUOqju7dhevMMzEfxZbiDDUdaCaICCIZ954yCh88WhlM+YQntMRolq01
BRZJBj6RKE9Z8fz2tI0KO7eS7iZ7rHhQb4HvFnmfvMqEv93Y2QjdoTydj4iMzxm2
aD9e96EUO/ExQLYXEu3so3K8pXDDH0F8T+xGApEjJKZ/lg0WKCl/hHKnMdd/Sb4c
wv7XwJXjIWXjdeEr77gRktbKQxs23FQbpZ3r2pQGz2ao7KKXgZD6O2GX6nrNyY+B
I5MpAq6FMDAyH5d2bVEvsGquiK8mnW/pgRhv6kOw7yXHl+wCr7UNJoiuzs2h09f9
T8OZmO0kqA9xkAEtk9+k7xC6FtPQtAKfw+l5gYVzd/M4CwFf609Dvhqq9nYAnXNT
Hpob4Nux5aRPwqirRgir+CpBRDGTCjz4PMjFjlEGfWSoZV9FoXyFjlUMwanSGhFi
asrov0UQ1U67WKD2OwAws+3FD/EJElEhIMBAwuoP7Q+B3CUxDj8lrtdMMZtpOc7z
5YWY1StWgTsjeNa37nDM75JYHzG4+azLhMRGmaqbtv0kuxDhkriUBLsGufyVS9HB
QJH8faO5oGgZSldNM1LCp4a+Jajn91l/Gd1lWN05GB2ZPt2xldKLlr9CPsNcEMI0
E6ECReOIMgUcjs7jnGA0jTvF70wrIfmeh1w+jBJfDQeS8W6qMYZSf5zTZEkWwC7B
rCDiGP166ovRwnsK2Zts1kHG9bU90qjMqFbA+Ta0sWmFEhYAFyTlgsDEev2ZHsFO
bodK2+s99Pgiy8FSNe9eCf4gZCvSLx4pWPYhlaj2GeZSqjI4g6WDyykhJdwa29nP
MBtiOcYIfrWOFeBhw2BirvxulHjW1swxK4kkucwdD5t2kekaYvXxmlfxPSt9LSvG
nEuL6OEDtxVDtOZP9islsHLsKI2a5PfXN5A3TWo9Xj/rtg2pRqghnU0ig8Tj+6mQ
dKn0jkomDDXM2R/HEf0nrwf4LEKk+qhD0EotfyQOu2VLUMlaJ8N1pbSwazVAdoTx
BAa0cHUdY7l17AJT/7oGPCeGpFxsvY4LcDEuLGBaZjeDiG0ZGPu2PvzjPeVKCpJP
By7SeHXDscPX93ZtH1DjuuOBbbn2CPAXGrqH6Wdffj5IIcjyvQEcfjEOczUY6APN
QBi7Vly3TcCz7ebxJSiNXgjXGUl9UZhC5vSPCHeeiQZaov0EPv7+eUOp/SG8OhdD
QQXf/826UkXEpkrejL7Gvi2wbclSsFV5ESrG1+NRjMeHpv93nmstB8XWAx1T4htf
Zgfy3YI3fwQkmT8bZfdI9BmkKIV1ZUnUc0I/d+fNmcigw9mx3hPc1NrAA9voQcJt
8p9tful18jI+/SNgqM3jXDlJ02IF8U1o9qWmQBMtyHthmvLeCP27Phcg0v+9VGhq
8XwqYq3oLC7N1PcuxSqqPh3eUpd+7MTEl83teOcmGaRmuJQgEyh4DJIvRuT4Zl/j
GE39T5wuVr0RFpr/jqQNPCAHPEkuLq0l93XEAl6HqoMaZ91id0UJ/z+xUw6fMfAV
ODCvociUrqEH40/O7pYGXW4zL7zXO4rSlTomjFxP3CZ0UpFkbN1rAVvSXdDYcfHc
7Cn/zPFQq0kp09sFPUPzOV3KkPjh0BgN2G8dbOTO+ivVPOqbMO+1Nh2blKps9AXr
d9RpxB96Hj8yAgqCjfwY9Y/BJmPNJF9qRN91mFSD/PcQcG3wUkPH1o3P4FRxgeUa
0/oxLP/fI3alQsXCfTFb7Qv9eCwBTPldE87LUCp5AXTgYVapKcPBtGIP2tL28B5D
bVcs5SU0ZUcchBb1TiEAYUqqqFuTRneYIT0Xpm5r9i8vGbZj/7LKWc9a5i9chz45
IuLLFwEMoLxrJaOc6FAten7HCElsqlnrFlr1OTl6xcecu18XvSbWFdU4kIBCE2lc
AsuBVGyDQsakQ1CiJCYf6TCLM6JhoCcQVYPezNMOL7Rdgc3LtE+VGDZ2/peCyqFr
jEddeSU9GlwCvWaPf4O0/dTFxaJP4Isgtgn6jwYkId9X6W7ZXZbU4EDARU54qqO7
t5VxeHbH93DhIMiyrKBmdUIa5dp1V4/Ou4dELLTO7QgJsMjTBUmbZq5oIHLFNdnG
gpjs4PKpbJaQcKGnKlWOR3mmxQ943/e6qoWS57OBASkQ7FzT8KuEG65ClZdyR4RK
vJsulKTPuZbJnQ00q6xsXx7lO7wP5SMIPpDuu12R3furo/rPoxhvTtsd0/U7YHPc
mI4buX4ljxgkLv2R0Hsu5IAXHb28F1i+qLYAldjpUYXz223y6S1kFqIGDCJg48Jc
jEY0okrhjp5hjthrVmAT3XT3EADdFfIHY1DqsMnRye4YrXuYPmFO3zF/0b5tOVj4
48qGj5iVPdGmVXaTXLAoQLDHnfMiE9allDvyAVyzGhHX1B8L2qPuIozJo495U88h
uAq3ZZGs6XGQjsHd/AGNcxb3Gcd5XIhckiGJPgBlCaVE1QZMcdQivLZxkvx/3JFV
o8ihukLW9ZDPSi8DJkuHOEwgyJWEoQyfZUANwMhqAALt7aC8lTtCTK2jfYRGZGZC
TiPtDDP6p6PD92K7MYbt+DUQm+wSSn6qTysdZHoIYNmxe/+il9P/gqrz06p8z/wo
+NiWIlUSkJdoTpHmKlJf3erYuoGGHUOMjTOYTkTuqbQzuzyGSrv88OvrUdWAyYbi
40aDbgounNCvpT1M+QK3rPKWv/a6Wk4TK2p0bUkMlpF7Oy46wCSKzb6aKSapHe4p
V/FrVQWEEwUjEAR/mCuF70sSB/seujP/eTtZ6TWtPWgzrej9oDuOnyt9Rzm6RIW5
Ji02FF3nMmGGMsB95714H4pxwVKDtsI6dlGO1ikZ8pBXaax83c0k1lBVlELTFUA9
sFWN/qsMToP4v/ZUBfzyMGP/1/1E/VroboHO2DJULqToY3JCGfdy0vjSt2OMPDQv
ZVmMSICp2sqwDbEXk9O/O28npNAbaV6AbcwUzii66hGrNpkgkibd6lHtz5ashVuR
5U4j7vuKeM6w5AnP+PdYiw==
`protect END_PROTECTED
