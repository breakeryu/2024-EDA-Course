`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qP84PidV4dDdMAAVbN7qq6k94VyRMUzXeWkoh3Sojt8frGJDU9G844pTnYu8k96y
DBD0ZZ6AEFYHkcw/mAUcovPHO8XEoE5sofpj3E+SaUdEmql2k9OlySROoOJo6vpE
KaBLS3h8ecIymzT5WXU5hDzn0NO6T4meip9JgZciHUWg+Zf8M//CveMTabo8ZlcU
mmxewAy4LoNNTU1MF+UX4w==
`protect END_PROTECTED
