`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1RhHPm269M7KtzkG/Mx04D5nJSfr/bSYsfFBidvSeD6UzbKTvdkC7grauWIYP8KG
2jNIZCNUqSQnRVocl/tTIt9the7+dtqbjJdANmAN9iOcgzEJ9CMN2S0HTfSHTexj
xeYlDDCYwnpYiWH3enxlLMKvqHX/6kLi1An2vOve5kJzbgCFhSMUj3uPRRfRbUWA
LDw0r0LblhxOlj26dAd52phVUCgvMTqg1VweYCGAU6lz5JamR3/rLrK7V+13Jq3B
bkM5j0E4iO84aHRLKAwaxVqVc73Lom73SY3GlMFE5o1si/1wiPwTwI8xDBo+TPmG
Ts50SnMIn5UFkinEhrFd7kDX+05GOLSqZjTu+tub0ZvJsDh7fK4Tnvqqfxo6FrP7
muQYBkpmDFxwm4JYzK4Jz3LzBL8/ORZNIJO6kcKrd9g8Y3HiYU8IBpi5NT9wuKJI
RsvVQjxaPuHl+S60cfG2qEHmNEI9uGlUPuUjg2KoApCMSDcqOkooKHusJZ0Omvrw
qRvZCilNDhlezd9TRn/PWZqbNqPqskzGDYGwl9WgN5sw3LiQ8lTJ1fSj8NuM8tAc
/VfOxPnPnXUt+hLthUrtM7f4qrM1g7QCyjjoPYaPoLeGFaM7qShBWo6RcIqL1C7l
x9tQvA5P2syAfjpmey4hy0nT5x499g8xGc7IA53w68Ek9f2u/ltd8Zr2FcsKmwDm
Syg6CWVcKlwpasOd0TUGHYr4Zi+igtiR0qTwwtf4S8hNRPDu1s5ETqdqME2lY6hV
UNRVj8ds7AbPopDR1iKuOawVcL6raLTyspmdMzs9t3X0Ll1LcvvQC5zUCjapZlIo
6UhfiC1XpAIo8aadiFxvsmp9tpdFJHQVZjElLOMIwXSXYSrLdCARNU6TQAYDGwK4
EZZbMbhMHlKKogCHe9UuqkCJFkA7LhCgxRTt7Wiu2KqKtFXV5z5FSbejKOBVjeAm
ge6lH6ZbK5RH3IEN54hn0gXT90si2X+8uuy3N2W5I/BlgohcVeY7YSrvCPPM7RVM
MwsQecJYSBW28pC2JgxqylbpUH+qY2fX8WC1PMHJR+mCB0HL6rmChNg2jVrpuJf4
2ijDxXcvR4hvfqBSTq7CAUh6Zvdq/Iaeykp6b3ey2jKUPVndLdmr/DRqESBIUzpN
ca3AHNvMFYm2uCw+oJTlf3UvgSCZKDHil6a4tL7dPvqocZI6UivaUPPcN+BUvA2J
iOxsPuG2XvGlG/t1SlCMHsGJmq1uuN92Xde1s9w+l9u88CpKm5CWVxo54q1Av2zq
IRKCb7OaIQBDMpVSp4l1zuMcV2SnY3JYyfng7GlQNZHo905HTfqh2YyZePWCVt3S
I8AJsgJSJ2G/J0shvbce5mWzdJeOxDp9pIVb8+iNU4g0H+rUqCWms6jlw8ZEz6d6
QFwkkBg4QSB3buQAlwgznvYvSN0S0mLYCXtMQhPbOYDVUvTZwUZtVlLn/a19XMV0
Fqoqp8nFrdNdnV+EQBmwfKjHaOsx8n2jEBtmy1f04JPjyVqXNVU89gCoxXK5Kr7B
fBvdNIaSWh9K1LLoZTJghX+xdfjs2uZL5Nm5m6jRluV/loTcn+yXzyySlMWzOuXi
t338GfMthRFaSraE7eoXw+86v7JG34AMZDwrdN5RNclwCoJXOnbrRlCeWPLXj50Q
+/qFjt/sMN037sLqzpeTMzw4a50HgEwR1UMzmY4eVnsnAaehCjE3kWrI6FsXP2ao
z5mhlAyhUmITKrNP0JK/ZkhZ3HjguvIO8cLMkOFtQZ2StHwRUVKp9xUjPg/5cMbu
TtmcVOvswyZJdRnIKHm9NQoQI9TR57VTbx4Jg6gknt/Nu4JZf0b3nSXT1afs/Q4b
DYXXT/WL+szwk/eMTTWukrmsBWB/aiqX3S+BU6y9xucyVFJeedCLOr7tdgojeer7
jM/ZjIFUONEz0drraM+Tu8Oth2CLN3OCwddxGoorNxuNe2TTIsWzAQPkvOzzMwng
lWnyDgyerjB1KRUDoQd4uelJJFWz9SZ2mrb4XHYaLtDZ8ZRaP4H2dIyCIqukOOZS
+ie1gvCt0Gwg20JK3NaCqj5VQUxy1YbgQbA+1iK201LwDgqJEX/tKPCeNOrD6ZBq
KqsltF2iOwowjyojmXVRwtKTf8j7q2BJgMtyscj2rwR6DmON5/+gEuwUR/W8GdC5
Mt3vXPU+3GOYQEj7xZw1EFbfJMYt1G5kI2NWOaeFn8hDIldaNwqHrvO4fpDREUXc
v4rV7wXAHC01zFfSEZKPndIvXrcs0URyidzddMvm40syl/rupkqr+EqAD4g9ipzw
0G1sd3LsavS6l22eWrK5V2/8+PiVKObLK//c1Za9fsUOVck/kP4+RjYRWkA+Iz25
vnE0NBp7SUPRAr/2aGZcbHzEONkVI5igfogARxxOdTi5l3cwO9yvDYZoWJ6uDsAl
9eF91mZkTnoQMgVZDo75WLEukc5GibAYNpcGxbFT8i468C6/ROesZmMOLq/3jXv9
6omzLI5Twpzd3pZpPdM/Omvpy4QA2xnlVqERqcHNkFWorXrAaTWtg30drogbg6rn
zTODVWjOEqyli8H0yYr+MD62znBBFCcBJLowbr0xCVXXd1E95WcWeGPWZytTlR4H
Eg60p8OwcMk+IWHh8qw3vcJ/iF6e3lslmTQ1qf+OjIHUK8J5P2+ITB/plb11iD+S
AeQfetmL33FmyfRXCZk4ji38W1zie8/0pMMeEJEJY7dbOCvEhaUi5Z/yzt+5yNg5
u9NKr1IrOEq8cJAWlcEAvOur11T5mrYLBfj6fYmHF1ZXHFH2uYWPjpH02/L/xMGa
3MYzKcFh0q7toqlkiIh+LKy0q8E13CF55LnB2pBi4D/ThWbKVX0KQBanyzbIkEEe
ErHLV2uCZ8gTICJi3dTYh27Zeav+XyH40KQtuf08A6N17UlD5Jn+x6IcbYi/M8HP
UsiV0C/eFZzkCsK0YLjP2VB0cZjSBzUGUgYs+hzkBEEP4cxmsWvCwZ8/hG71wp8/
mj9aeuiOwYQPgBgxGDyArgKJGasDW1jItAKOcbULzH1tn1jySK9t7Jutjpin3fna
3E18wVjcWOsexkDAF8z7Xy/4oBjaskElLceTGALdfX4sHrwjux+/3z6za63ZZw+7
xGJDFLmfrCJuJDzIdo4ehO3cMcb64rbS5UIVmuKh1vSbCdrxG3wMotHq1ojq7QXP
JBvHCBGRAckAZifh0iD82eyESRpf2MiWIY035Tewc0rIGRNoXlf4+tkrUaHqzalF
p66IcsdV1oPlNhhkpVOw6S/yAkJ5+sLeV9QdUJkcWWw4mC9uXpTFejuWLxyQA2U0
62YeL/wd9PaJC6qVZfl60VClX8MJeV4zCbmLa1DP891oFwsAtTvQ03feAJsV7XRP
RT+a7VmHSZTjWEzI7s11YPw4LT1x26LvKO0TNw1tXFJegTuz4pmgMdACtaIK3tnu
MH59emtUouRH2zrvwBIbnLDWJkIFihxP6b/ABBJM4NsAX+aHA588g9roHsFbh3a8
CX7VA90jAFLyi1lZQgEbfMAAgUSePoxNZL0zSEddEFfZ1Yez59Ax8xo3RSyOowFw
PrjN790SvMMQ7tlATB12QtnVdE2IKvbzG5MJx5bcsinHIdjDNWxh8vMtpz0vaZ+G
5PS8lnYDlseVboVFmhWfVA==
`protect END_PROTECTED
