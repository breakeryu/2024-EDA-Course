`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgS7yVBslwcDbu4fUJMKMIrGETTCUTRJqMRhWlDiTE+Le5So+pxWoJs4pKRBNjFy
eaS6PdgUiPVqCNuHgflhHTH3m/2rvtHa55TfzY5q+IQrMgOznn4V/Fz9R56I8tbn
0sqlel0awIXGVLTC6GBFQ3EhI7F7rTLmkB9RmUUOgnFFi9tkDilsNq5WbiDuQLKo
Ck94k+nx7F3X4r0XCKCMVG7vjLYjXozrLdV9A9Ig5ve6w/pqU2a0/A14dTf+BVnZ
MRBK/E6KhyrrnDuvBvinU0gNLo1+LhbSQrtDJp106IyxC5J/DdpDCwCSW+3URQbQ
q33XwW/tVl8HSTwNHmkL8PpT7Y1axxeXEKu4Wpb2Q+vtnzr8LkmeDkXef5omVoOQ
ddeO4r9nsT9raI/LIvOT1uIgIPn1BAhhen6nAhnhTDWmaVujnQsM4oRNvWfKS9wh
8MkNKX2GnGMPnIP5/Gs5v/xD4CK8S59ExQeE40DRUBd0t7Q1nRRJNrCudAPlxteY
O6uDRh8LNbxKZCcgqpXKwn535Ypof7TU2XErkkpJpypnUCuKSSQBMG2HGqwzhcQ8
NLKDzNmiii2HnzT+4MQ1tHQfRQxdewAn3/fGpsgt0H6s8deSOGEsz9XaMcMz3VW3
IeFhQyoE5ZMokEo3JF2P8+1vERAweQjDGZlP8TgSd9LgV80l7ZlgesyJIvqQEL1m
qKzXNTBrLNgaa4us++gW8cCxqRDYEk/3E4pHKKulxGAYo6C0gee9vzidmVDhzUDs
Pv0zJRO9r3DIUVC2urjKnWA6Cj9hcBEoLnpScm0pwClL4tMOXC+isIxQBbo8rNaw
S5U/VqwnFpwEDn1ZBSr3ZJcz7FdQSN78VIpjYDIkwrzPwGuqpblaKbje1SnE87hZ
4wjlzyOp0yGLYiRsgpRol2j0J3Xm5L08pzof5dX3XOp5Wn+nycUOSX/7L7nhY37K
BmYp0TeI3Hz8He1nAGukNFjQZYyBp9UF4rlV9Wi7TWQT+Vy03vb1EHsmNMVs9Zaq
C4/CK9iNRnghrmxFYXBlXxxJCDq92L6cmWnsoZpv6Gd7gI6VCHaKKKWX5KOEsgvR
va+0cVPiQuWRJdeKTMZXDpULVGlwC1FBt8981UuZ9zilG4DcxpGXAP1iORo7jpdd
9HYE/PrCCNohgQ1+M1tuBl2wO6oxG7B+yubVSpmd0+fwmL72F682zEoH33ymENyX
WRNL8jFG0d3YZD4ko5LO+TI5ze1tkIfHBsiqinYkmnIcPB3UTwxe6lZ+cjlATz8K
D1/siZh56c23x2r8IWfGwvCe3UsO7nWjpQI4LIP203NjcNa2JeD9Kx+lQUd+dAHF
v3eSmbpun9f1NEGDp4Wt7HWzOTJVaolAvaiUHI6q3WvNCAfcz5Ld9tRuatwJw2HB
6cWjc9vkB86OxPmvgSriksDmJqnyDbr1G9DzL0knoCY4G6vnjJG8i7USlaedfizv
sba8gfNmyG1Ukaqe8QBABSnTAryCrC8hd72ndvIPUwDtgpABIvMFPZ1/99jeTviH
nFJKnu4SBr2eIdXzPrHlMexQN5HZusUuZ8VPCXE9x0DC8t72S4Tnzb7Fgt+dvkUV
j7LIPLg1qhBnJJnm4Wljt2RMSx6NOuJcKbUXr1QEgjiz8RxzEusfCbTljvA3ZAcF
W2VfAD/5jWtkaovHN5b5VGTgL5XLNtsW7Kqu7Ykc3af9Hl+9rTATYdpMMvUi5VrI
o/KWbl5zuAgrAL0XHwBdSUL8RZFhX0v78l5KiJBX0VoG7Hx8JVpXXUiL7kt/11zw
cIGfwz84cv75nO5n6850oWX5xMxb8bPXbqbHIayguCYWCVHu0vrt4UbL2MEc5/kG
yUIia3qPdYFKWFMdnRoBoEKUbjU218nHLznIrV9OLuHYqJ0qHyA1+HCyJ7BUanWx
wWLdstUJMdfDApBCehMJCW9jh3nwiVfXSfEDIShJuWHOBduVnpJuRRk/FHPGP8Vw
3j2o8QbeILKQx++kyH7kWzbq8jDekUX/L4S2+nav2b/b23L2N9f1f8jJYSc2Fqk1
QNmmhLaeC8mcrL3hS1s73QIuUn/Hor7NHbQ1ubS2CbChg81BvgTbX51eWLV8S1TI
ADLOC1q7YDQblBIJCYmQ+5nxGtr7/B69nz2f8DTs86TYzq7/oIsZP5iHXq/Tzqw0
wD0iZSKAGCCm291+JLLYDdbVzeNRib0Bk+4ne38g95nrSJvQvTVBygqHETOQni67
+xQuPjZYaW5eJ59/lGsgq3FTVXIaPMSC5NPviuiGejWf+ZmI9GWXMC2eNYi9lSXk
kEVG9wxKg1sewEo4sSkSw1AVJLShBG9VX5SOWYnTCMt86ooZrPswxSnzUrQciPgU
a4FA0dE1U09Qzbq/apdmGyt4JG+6U+7+FIZL1wtzYzVdYHGb3hfklsoByO7DwfkT
28t5X5DR/Ux+pL96VX+NsT8u5WH4porYBsPB0CaUu026Jonx/wR+dzOriJp87H7W
0HJ+u8pmt5jUvmWcSUzCxuZjOayxa8w2W0qOFIyU+XbyLB1s7vW/aACgJoRf0olJ
/bXaglMYK3v8KPFp8gAwT3iHg5dAXD0ATleNhzGNb2DnBJiZcojs1psMaxggR4wn
UkNjKLhv5PI62ALePa8obytC1axJkWXNV28S0Et4lPnOvoHnDZ3ODpDIBuWzH8kf
g6Eyluo9a3VOEelm5gn6oJ5TFW3HsbSExOiY4aQEgPcbahwBI4H9AWZzPS6Coodk
jspKw4TwgGMAIyBilliyFxotgmjLhkTrf6uZSwM61CYY8KTZoadOkLFvX+7xC4HW
zLtku+NWCQKcXwdzSPHy/s3E1dE605zFdiDsm1ZAqjYtjhT9T9EEsptnL/Pj6C/A
U2Bed2L26gX7+NBjaLvTro+Vp0H7scALgIqkvYar0hBKdsniQKBp9Qnb3A0XYKEL
BKY8mVvcJLVgHlUAQ3G+v7i3ljjo6EM6Mm4/xEEOBVmQ6Gof/8MaW2LpiN+XLM1i
D6YqqKTzEhWA7wBwIZ9UQ52oOeCxiod6H9ur8oIs7NCla9zywQ4jq7HqG9f8jiwZ
4TXZ7jQQMm1uEoOmYigZUtvO1pu1XniDr5W8gfgOumYB/+AXfVnCkQe+DywmcGds
e2z6/rIdcQ7oIdFhrHRAROR5sfZd70p2Tw+P4epAEmI+GboA2OQof8WGaSfdL7r4
6M5zsANwLRY927DCLPwOegigYWvGou8MmVCzpPWFFrS6Z+O+ZJOI1CEfas1kxoZt
lH8kvV7Tl7exUM+jJSEcY87LDtyU67lYo4E6v/vojHBNA+XFshZCYUM1P9xy41P8
lJRiQiSMtsu579wTiU7eZc0oQBSvgZJ0DQNg+s70zKGgd6KUMGgHDOPy4qAIElTP
ibRQ3ozdLtD778h2wxlAAmwtHYJ8dVqxjdLLFRfYlR5TncHPvIcDfqIB3Pv8AcgB
XlNm/5uvXAAst/K+0IRb5o6wPIYhA3VGkWan1PllWYZjHA5WtE2LwYXMn+0PPv2c
ESwTDk2jam9E54Z8mlD+GXy1wUqWFgFwLBUOqXsRDIFKQWm04dtGq8PmsZi2SfTL
i8XvxEVPbGp91tlswej5SR+K/miPLK5+W5UZF96uBPdRChuJ/MQvmosW3iBIqj6i
wNuSPjOks3y9rMJ2igJuViKDypDcKPNu2A4zVt6k6OYaPAAq0Nvz05XIpkuHQhCT
krVR6gvGFdzK0HV97/Yhh/GtOAVJ14Xwnz/rc2LW5PGRQIXFSQ/oaBGCWe86sWY5
V+hQOWN7bJKnuF6JeqAfDhA0yQZ0JIQhhVZsan9znUmq0Ec979PEDvZXiLCBdOFN
s+rwGvkzKqnCFcR9Ra9YWdccMAn2QN+kWnTYKC2hMRWRu9TKGmPfWy2mhwM0huPI
lsWvkjZJM6U1+Pby80/YDwWVQTx3MdTDCZ5uD0HHcTiRHU+QRvPHxfKYLhbZ0oP4
cuibC3LoMFO+v3VUq26OAY9DrXpA5OWTvBkZqnj67aKnkl0orByNgBCGFG4jRPS0
bb0EsQsXWopWZptWTQeEZBjdKL8qVtdzDBqXr5hqgwcVNl9bWaydMBoAtUnTPL21
oTWLC32Eb8RZVg/bqgDDUzLqLf8MjehcpsyWmophrpCmR+uDjEQblqAbcQ2vK4ad
Cf+tl7aGP3Evu6gp4i6DwUufc+iV5serhmGCrd906QWBO2YOFZr3IavgiEX52z2X
pDv3QGH+42G00BI5xkeQBUA8ZbJ1hlPcma+iV0QceLk2HqD31jhvQtKH9ak3CNvt
LjOnZgFWwXqGBs3Iy5RGgmTJN5FDIXA6ihznWzY9JD+xSQjl9fKFNv8KTIjy1R3K
DEdEA5wFYELfPHZgeVKwQPQfI3U4Mi/rUp6iwqY39MIzkPd8k0UA1iLlzBD4KOpR
LeW+ZhUSMIUSx5ix7n6M4DBj0oM+IOb1kiZHaXDc0+WEmDKSgagF21a4sQLn9NbB
w9gZYPyUG0ZM+6BJU/S+8VsF14zQIm11Zs0bwNgslJN41YTY5tPgJT1yMOGuQEJQ
MXkVFx1g0FOdZCNkzFzwKfW5qvoLl3P8XalzzV0t4mDmWt8Ak3jrUJ5v6KeQOhap
oiDDlEBJdExtP/9zP/hiIgcwYTliViAiZ8rgweal1/DDYjytryRfvbG8TDK9T7zb
CaB6d4INimZ+LVbsZRzGnc0bMWTI4CNw59tZBIDRllmhm+KzyFxoOZMFmOrb+8Nc
A/8XJNbS7OCIYQyvzIwvkDy1KZFlbqihiuwwTfbtq/Qvacsmv1JxD4GNus/s7yo6
Dvq3frZRx/RvIxj1gDjJWnSm+heQBlCPwRkjzaPy/Os/Gv2MipUwmyPCjObcSMDL
e1+MIqDzvmLdBuMRQhv8eq+y/2/YHCNU57HgEfWq9WDH/N4TvqSF4RBZtI78tyea
fA9U5HEFmLdTfSsXeMkuBAEM3T3Zw38Ayfqe9fjjL6rA3uwuY0VqaCVOShKmkwQY
gAKpsDNJ3XBdWRUt0ax7Q8vtjK18ipGhWf6+e99/3kuL2NfcLmw+KDDFprMG+flK
RiMr9/PvXxlcMbndMo0Tomt7ZTyqgCDU2nUQ/TT0aOpRC4BN6+TktBjxuchPGh/L
b10YivYoATDHTyqquMk2mtlqY/K5TUpHAmA0yxw3GWqjIfgoY75bnfg4+T5Fqztv
91cJL2k3UDuDlvoTHEaMoQaXO3ZVKJTMnwly86bqFpPz+6zMYEPFMdISfd5swpEc
BXo24vDJ4xZMjDrCkZNqDKQsrvW5jddF7imjTJUOOdY3HnrYUIN1l7rzIQXaPW6b
DkNv2IZgJlGoX6lVafvofrrnDC3N0HHSjnsNBDcN2kDnYZMP+gJaZ/E1nWG8PmZc
shheHFdIq0oOHPGoIWt8SLirthwr+4qMDPlwjFX0OFCGSFRjiTmjfdC6QvPlFK24
mgP244inFHNR7Q8QsgeoJLwuJcVjDyi+3rhVAQEWbR4L8AeHDB/lPFHPnTAsuYxA
RcMpBXyAVLRHmelWhlPVtWTeWlixQIf970jsOX6LEetM9W+u4nILsne5ai3x1zuH
sE1Gd825LvwffGMonDugwabNOudAvJgseotUpgtxlTpzSMMPk7AGm2lt0cuszgc7
57tgov74fSUUFAn6ABuOmvBcpOpl36ph5ZbFaWW9ql1urewKPTEgztQe28gHgm9B
jmxhCA70UwRedSmT4Kdp+OdsGvezFtmlmL9Oao+M/ULXYGYO3hkkUVOWZmFCttWg
EaigCYTX7Qc6bxrkNW2C0Q4KJjTqMYp5dZcGoT2UVAHH3560OhAsP9DCe4l37/OL
8OmcgdLfpFdJG5QrQ1j+4BxhqWcIFWwg803lWpI9qQARdO5zCFmvDQuKz/itTz+D
TAE3KBuUoZDagusrXd0AYpwqM/MjCCn58rk5TKi0LqE6yLfAx7sMBXZ2uN13UgVd
egCm0KMKM+38KNWxXEHMXV+fbaQMm7rUuWPKtWUHdb0wD+oKum4lsMjEkhJRYXma
LnixlXcTCL27v+27Yt0BBUG4Gfuye3xtwvlgZS8xlU+d4Ehzlpr/zl5rCES1tbge
+LaylQTthcf33UHkoHCrkLWJ6ifjGAVUtRKC/T1QsilzRHQ+2y4QjfDgKcXWtqbG
gNIfOUj70SjR9uRGEKGbz26kUwFv/lRfp9npjbB0R0GKLlWaitaKzqZ1PicdPjV9
zHu5DlSBNtkOEn42hDx8yBTkGi/nfLX80gTNjIfsvP2BZhS/KFyqPmVF1c+AQTTx
B9b4Yoxom+0vWzCLDLS2o5+pFbOd6f8QYXVIk186NxfvkxXd81rmpm8QxT4yk0RI
Cd7r53vSXIJzKi17Ye++A5bD6KTwLG5JZPd1l3kPHC7AtX6lSNEiEqRbsmJPNR+t
PO0g6NTN9dY+NDaDiiI936J2vIViWVsMuMg4/hz2d1jqj/QSiEv+nwYp62iMRn7A
aPTH20QTkcxQ+bZ7HHYbrFdHuzD2+H4siYYciwQFJDnHwxs1O9/PMiqyYibJjpLy
ODkoiLMlFEuG+OYG5TedpSe5NnMbwpmP3poRDN1u2S8PlydLDSusa6qRurK90C7R
zkFREIfc0uQsQJ7HwDMj0TlSrpu2ttPjM9BWXxJ/QzG4UoXPCOL3hvbUAl0OBaPo
oQpByD8MIEeUA0HTJnv8Ns50yvFagDg/MZmR3lj+42vomjhSIWj+RGpuOCHlG1A2
crQwxskkfMa9ha/jGHfHGa6KNyaONav/LC5BqdfqdOHh9wPiWP3Wmw2mM4GDzRe2
kI/UpnsQwUW8boQe6suKpmqETambmqMKbjDPbVbaz4ZGSD1+GDO2O1EIRT9NXqNr
1vMAbWEibspL2wVrRvcQ4ytmxh9lewk3QwIR/rAqG1D83PqexjQ2Psmxt6HU3+KD
WEQjp0DveSLVXPu31K56Zrbi26hsI1MAEgETJ873g+stOTxGbVH+ZiTpSHJLG13s
cgRJSdpQlG+Vu7MkYs9bv3J2x75t/59Dn8EwkqLP7E1wLFKyVZxSYeEFdFdF3OkO
hXXpkRcYbdkg22Os5nEAPOf8Fs4/GiEDG/C4I38oMoQQHByoTqIa2SmTFd3e2R1B
n00FZn7lxdV8WmV5v9zob4izezlUIaZ+s/GlduUI8UetoOS/FjqNJ1DwK+nj0SMh
cex1ACdMDViBh8ClDkxo3D6kfslnbaxbSXm5e/1v6Bs9NKGuUUNiPZIT7ihwhLFe
xTkiTpQy4F2O+z9he5I5wBYqapEXQtNJYND1KcHJL/JEXCeePgarf32Q7SjMCio+
SuvMoMHSDkLl4j7BHrO/qQh5x4v5RvTwjobGkLZh//9hji6JSq95Ps6O/pMrmBqv
vlZw+BtOQb7S6mpLp1C6HrZRvPolJy6Ag1QyF3+EzsdSvgFoZeBAoyz28QiTfmc7
2WpE2FM4KQL4m+aNuE+FJLfK0p5SPgvA7gyHtTwURWY4UX+NoGjec0JXJzLVtXZQ
0U3LF8xewzaeVpu5PK5G1uSrwN8n9rGN44atqrudQ3684YoEbXz5FZIFm5JZ7Q4+
V5sjm4Y+C66O9O+jIv+o7+VuA/1GW+ardpvU16zddo8I0HxhrvQtrWi4lp/08nxw
kNRQDvfEVn3sH42j4ZYWAgubWgTn1oc9jyCnUcQlKryUFdAZJM7G9E/u2+kz9WZT
PTJfJ3mPOOVXvRnhYIKOsjHuxXQUZVv0qk57O2UxvNNEWC/AiVnAglA5iFsTHhbe
aGHm+jvWWfzSfCaM4S0qOfqcQi8ZCg2UIM4AEp5hiDtkxcPMCgJbuuc9Zc5eIOcV
d17VCVLylbyC+0ZEsKtUKF/jKVDzk8gpFyWPQRnm0gXCniUwqThJz48qQgp43/67
6Z5VBE4AU4U1T44SOTjxBhDd15g8pH8+VL/KnNmlgVkpinma3SXvVTfsXxOZK1aP
T8xS2ylVeb6DqD2VdVRjGdkOgEGRyPEKyAuIn5vREepUs6IoXZf6llOKOli8mgEt
azKPvrwdfYTc6IUSiwSU5jNk1KN3s1bgPEp9W7vg7Gs2MrcDRAZCi4wvbcTzM0UE
VLyhz3DPybRlygmSfHn12aXdLXvyDEAcjX4bcvujnY66MlkKmUt9jxBk0wr4h6rr
JnfYZvirfk6aw08OvWKbqydQM/5PN3LZGRuzDzFBGS0cf8T0qTvza/d+w/WlNg+J
SfcmZnDtfpRFriGSAjGkQ1dM7oZxHIhW0zPrSby405i3hxKLzzUQtaaDwtpbhIJc
MWeYfgDRiCq4KE3w82GBAVNiDf+0y8L6bYDBnPpjsbrqNRH/YjdgUf7diUxH6Rp6
4y/QBxYnnAUmSVfIUxPLOsbeG+fuI15H61kZuDX0bPhfVtRPA3eRg4VSdN2Y3YtK
bTiPKcDlam1yS3dJaog6pKA0UqpBQj4fDRX/JvhP1RzLuyDheaectscf+Tr3WvDm
qxK3cia52o0RnV3cXIIQ29sCzUqM/PhWOBsdtbPnTeqsknSllrSPB1DkGAYJNgv0
KDtXocd9d5kOWbyNoeWTLy8huQHu+d5BPL3ojGEAIzgSjvJUX04kPGeiuYad3mXu
O6iAazd5Sa1ISMTWM2ey0nsPkqVuR+JDqazvj6hgkVgYe5mDYITtE6m6SxPBB7g8
zmh7Zhsm36Zxm9I+b1wk2m4HqvINccKHRUSdYgHyyiTfGEaI6F8rJYEXtS8U3u5Y
hjSSwUOur4TY/AhTOoirNunH/2Ke7b72NnH098LoSupFxIMabCDEfh23Gaz1vW56
pCz4RLqO5JZLPFvhogbl1w4xuhgKfeqPLOQnfOXuaxKkfxVSTO2ojWVieIDb5Dse
UWg4VLzFdK4/7EPXzqZw9pLujLqrqH70SavDrbJQGZ9Hy8pNPlNKWbSyuXP7CtSK
jmxmBsKlnGYW1iZ7LpnxIx0mazlNOyR54vCSMo1Eex7lW7PLgek+FspFH28J6HVK
68sa+anRJmjVJqVlDiPq7K7psAH+kDQgePDsd3yM9OmfwV5jMYE3dXqq+ackMrDg
xtU+tiIdMNtNu+gacWqVCRXisGqPGh6GBpeIuTwmLk4IbIms/HICFv3fnpURxR5e
Uz8ocvdCe/EA+fVQY+4OqbkdS4kGyGP2LH0FCh2pgqyuPaE5UbsmiFm8A2IP0KDW
I3ig36ybJxAohlqmhVFmEL9j0ObdSN8baldr63Z2BefiDkWq63i+vGATYgf+RqrH
yI+OXfUmKAABw3mQlvDrbE4ZD+s/3XxRdVZolDfz9xYdtetzPpRCmfmajcuIFgfN
Fr5IY+Rk8e/k3yFwKCJs3QJIQXt4dhJg2Y59JbXX7tgfREDl2rhjT0oOStYSFBq9
/kaAoN/Gm6yRiNhEuIyOdiGyh8mZkLoHQKpOS26L0P5sPy1+CidxpynnlPVBWz8O
UW8K0fZXhactpWdmsTwE0atMclS+I+rLGCjcZo/3lAsyhX6GJ6jUcxnh/6ZFWOE9
ARxcbdri7RaAn0st0thp3rnFk5SJDTCCDq3QbDCH41g44GaX/SjhpSFeaXXLortY
Z8CxqZ6YkJQ9EG7yvuOAq0jHWYP4wLiyL7w7mx8seKtX80/m9y+HwJf7ebeOZjWf
MqC3jnJaPAG8dyjD29DBswup4R1Dgfb8AgjJaFkgDBY3bxL+GFh9DeAKTx9cjYlC
Yf+mPzboTiTCxzAzaHSUVKW8TOYusGyiF/2J+rQ8Kl1J6QsYX8H683CcBUEVLp+0
yyKbZCUCMjuakhy1GxcYH/o+lua4y7z5rXrURKGnHE2vePRiGzUwNvhqbyp6dskh
P9k4mb0BKUMGFt3v/bD894oxX6VExnWoRQb9zweBYtnJbyeUFC1oSFNQR/ewwZKW
tdEzx+xN/gCBMRuDzKAo5tt/aaXfEFxt5cfg4jGIC2ESBfmhglUVqncR9TmLDhJF
uh4zVROtJ78bHw5FlFoWmamKaRRapbRNUnYTd6qoSZqgay407BqSgfsH+lslCv8Z
MdZ7Di7j/Rhuw9mw6qX0O2mCJLjeCqWJihMCEaF6YQaMp57gCT9If+9d4CDgsbMl
OrmqxfQZ4t4WzIEiVAH3Hg5UHq3VVUfWfapVlizj4RthvJo5bDh3Z9EB29Ehi3Zp
EXQE2HK7Z9hO7yv2/IVcMyXONQK4kKTJy4QBzn07EqiAYnS7tvq526D0uN3Xuq+/
GWRhEbUTmPc7vyXdDKLoYXJ/mUv60H5UqLW0IOEjhJhA3e95cdajkwihP9o4RO8u
SGjJII+7F9A/ZhzIV5FDbAaRSrnZa3AKdF6ybfTF7X9LjY4R0Ta695S3L/9JQ8bB
dahB1g6xWyUuUpcJ6IS2UAt09oOQMPL/aSgVZA04xiRQsr9Z57Szw0+z22Uc31nW
+2o+kpr5Ds1bJWsXCkjHiPXywdYoy1ERl/djQBQQQKc/m9yd3iQwBvmqy6DAhMH+
uvyREYuwN4UgLNjo516kD0AE13eTCE+SEd0Ltl7bbwyjlAmmBHM6xaDarmUWSt0d
RY1C/0jyiEveEXxKOqh1VIpTY5TjP2kHL7ELqS0KWJaOODMT76m8CKWRm5pra8O6
G3os8DkVd2KW4LDzCuZxDwUPN+UhHR9laPqyOTNN3nn7HuS3Nd/Vao+xbixuZwzo
8yGpHc2ojc+0Vqgj3fJhEiqEeDMFX7yqLHALbo784Jg1b41/icTibg+CeaN1VNxT
Ssj1AoVq/oNjgQ7GyD/wnGHcQvHLvhNoTAtZTVckXYp/tmcT72knYcWzvV35cbXF
263fwt6FlHeZ78p2dol8kTj858cHIz1s+p1+17v/TO4vH7HjRRVNNN8JPhvZXhzZ
DySP5pKD2Eycc3vjbKvyHmiFItauSYkOjqWbrZxBBZrQZzxclTXhsGohPoQjdwBD
4kExC/MMMtFCTpxyxwLiuu3bqk+n9RCQq4rfgP0rEyT3euJh8F0Y9AjOsSkRYoB8
6BGzb1L86KDinYqS3oowFgmhZ4xnKmOtpyQ3GfdnhKG1QMtxrKu1ymvuBSoSBXmu
ooWxznLQ6dU9ez/3T6UP+oYEXBDOU0H4x7FEDTWYL096/8Z2p7NPAENb/pJ9CZQO
TdvgVLsY6oa2VwjdrxX9/TJIto1g4u1y8ERWjzJ7vjxhpFSseZyOOCkTQTyvmZ+/
1GUdYpJiqaqC/vfnkogTNHFT6wX2U90+5h2wnVR9YexNK1/C0SINDPTFoAOVMv5F
A9FvB5EOJuSINfM+n9OeXEgSPKWC1/a2H7Bjkmu0o36kFzprjIMySvDiDvz2nWPX
TL94YO8uR/l786Y0MG8fyq+GotX9uKuxBjxCT1WIZEy4Ho0LOhr1CTJDLd+ki25F
O6012f+KDmdcbwP6cdRH23XAcdkI+9V2qyKe54oSYH3oq+DnOPGIymUW4LLu8mEa
1xp3yREh0uHO//AAUA7wn180RD9HCx8mc6wN9+5rBOYiGp30gBeOnVSkHqdVo9ti
44U/dHF6F1WvpKf+EqOuqEduMQq5oaKqtJrXXe1RzGAMaufACtXA/bzQFwNjjcLI
qSDMiUxPXmJ4s6h6u3ANO8YKsKlP2oBNeFLNblkXH+1YfRuJ3uIXxLF2RxjoBtvT
LUVRbDF4Fj3ey0x40XKar1EpYMPSEucwv64zDpmcgEWR5LqS0ijXkZRhYbMHO3Ve
XwUgs0vFsp4eoFsMzVlBmYzQxr++06Q12u7ufhcdphldzFwCD3sqIpM3/HgKGox5
opZXhwYVnPV73jA7XiTJDV5kIuZc60Utg+JxsgV7GL4GWzyAwHrPDeYNDxbbnv29
tSqKMtj1m4fIryEbPgDnqJ2PUQSdkHqG5EPuBQUZv4o96yrJg0YbGnVlJLoZSw5V
52D0as+aGxRVms29achzAdgGh03vmmkFvfMzhlIE3bsm2tsJid9i1vORjcnFFDdU
mC9ji4cAJbcrULOWybT7FS2ewDODCIzl/9BZOZWXTAC2MwWo/Vo4spe59+aC5GE5
e9bv1Uqry+gCLh703MZrY2j3HuhXh/2QLAQguoFBY+M9CF8folD350wbk43QjVqz
SRfAFtOIVfR91EXdRHz1B4JqxlvbIfQwEAYJl1rIe2wv1wyfNpKU9c0ZohNYAgQN
2eu/EbKvebcyvSQtV5FPh5/HsjBBs1NrK29zJbOyJ6/wQK9ajbCajd0kCYIjbXhB
fY4GSHdwaerHDzK7lGjIvXRdHbCJPwyiqrGCrLGPycyAip+IkFRQZnKfdD+DPUI8
z/XIY//XOcVKAKPyQWrH9p1MXQ2UFDEDJIneKsJ1hM8mX1rA55dIbcsod7AhQTk2
Q0qw3LXDf+pMBdtUaoxtX/G5ZqjYgkjl1zAPPEU4dysc3J9tVNTzivGlRuOLZiHz
W2B53lS8Aom30vv7KZEXqDMJ31VWiJViUU4nAXVU9Gl+c0keBO35iaB41V83yYWM
KXXxuNevMfACdNz6DuDk0JwLFY6fi6Jwi3h3B69DXDOf+dT5jEGhKQVShgypa7wb
/t+D/KdhLn5lDdPWt7cuQ1qGU5i//iL5YjNl2iIuQrV2qwuIeosEwfrzAdIpmY5p
bMDOmb0ji+bmN3bpIc9qF+9s3AGvaXcD6+hpD3qx7BiKTojaynfjr2rtBZ3IFMGZ
1A4laVhUTI2P9UdBUU9RbCu0UsfMOJ7v2ZAhAa6ePsesr968A6YeSjve4BPtIUcd
mRWeWuHyl1zHclI9Ia4hAmNG8GgkiyvdbQnG8dU9jNbp5fKomZB8IHHQ0oLGzGJ0
2zsV1MbLFFqIJ5ZlGVrvV5TMgN30/v/3hoVf/vHM7i3TlArtTS8om4Jr/Hm6GxCv
dEFXj8fQuJu0yYmECRSO8DpMmdPfe6lG4WAAlFypNCxt7Mo1/oRKFOjkZEkUnkrJ
7yYOeZLLVW0p+TG2wq9sjVIw0kcloCq0yhHcaDNkMOSUKoilRqt8rzJponMh14SW
9fLSslKwR+1cAWyxre4q+rEmwWptL5hqMJ5x3fNJOvJHdifU8Fh6WPEVARIxdAx+
L7jSFC/ek/NTzDbJvulyNFEcG7aC+v6CWxmHsRc0or8KtJl+40z1Kjwab7DYzjmM
GoQnHqF0Ek52VpH2ewXqPTaj1edEJu8KGOkHWFCAz9jlfbQJ5VeLpsKBPYnDCdcV
FlqyZFo6bsq06jJDcIlKn81LwKub/D+V7iRMFObYQJBSUjMGN91ZUJ2pF6LygF9P
3TD/suLOjQHxtbDpzOlqiwoOdofcH7FpKqJ1ezInkelts4+FqoIUruWwyv3lpLf5
fV4V9OrnSRLLerCwPNKLUOJpY2l5xG+8vB/qdhoViLWPvDqpnSZJYKEmgSaK/c0K
GW8KdO8P20y2rGetQqgoeEd5/6XDffTnoHYB6jSgFcVLcw3aUUiTIi/uaygyevFJ
1lpQyze1nwyEFg68UUWDXeG4raixpd3xXjdsT/lfJRfgdX0Jpc08Q6SoDA+Dwahh
krgEV7g88zBlRSZNQujbhDw9Wj0TBnEUnplOOfl5GbTgQx9Ln+GJzTCdPk5ovFKA
S684mJNex1CXFGziEAU2y8dsqlcAxjPvFDlOldc95HOhJGzTGkN/lzzZUg49R5gN
F127eF1Ijh18Voo0pFDkcUCzP6DuGJ+ZgBOzI6X0u52uMdcAyGhhVX19TIFvO1pp
EYlzAOIQMkWQd+Lzr3QB9lXzAFHBP5qAo8h5yci1v5NaOCsuitVnbPGrPmG7NpW/
uFrYRJ5fW+ygv8IXlV7InGaGhaPdQ35aeSVoCFXaQRNL97V754TyetoFpznhmQNJ
821Tjk0lLnaTUmnZQkYFmU8Z+S3A3wmVTzgGX6LFHQ0BNSSj4rGnrhmSMz2NGvoa
DY+e6kZu8s8xFVhbbiaqV81LDCdPUO6YDzxomHbQwIgBvt0v1/nZMOyFQlK9VbLd
mRj9z+0BVUzNLzVUZNSDF46XAEovM2vWumcpimC2omIgCDwP06l0mxJIOpugLjtJ
WCRtvwG45I+39bPDTB94OHFiJQc6ThROk4/MArb2qNYbyHYpp78SAUdgwRqA8c77
f4i8qnA99LTeUvw4KMXKutp0WMXip/Osl9ro8XLJngYGp49AJlUbqTJsR/pSr33g
AkwuIUkBl5t78BZsFwYggYo820h/opNANYlsMWPQsPkS739hrS8DkY/3MkVZ3c/0
MspxKOR2Zp5BLrNf+8s5eB+lxDwcDXwakoorPtDKirh+anDe+akxiJUjVa9kg5XH
AexsvZ+qATewH6ZFWqwCz1IYY2jO/1QF/43bQnJ8Ps7YGQmNGW5JciQIX+P5SNSz
QvSrnjXBrAYPohX0e/fdzfeRsOnjxr1zsxlnyhdUqVrGGBBb8r7gaa5SiyORGAlE
xPtp0WLC9feduFWbF8DlIHj4MpF53PkAZR8jwHuSXw+UY/omWHlFENy47oHwwlTj
7Aw+55mydys4MX68eUd78ZJvjOEDyioIvwWmrVTUC+JQTmOwcRASMqDjr01Uys97
1gktIZfqeazt5+Zs026w73oZzErNpjmnHLIpQdMSSxKQbibhY0ckr3Z8JDMIBUq6
edIxSeb/PbFmkXsMih/nq3eCERVEF8Vgir7S3f01kGlJGjEjMfHlFho+qkeBv+3C
y963FYdGYUMIdfn75vp43l8AuDlBA6jMb8u+vE6KYYI85hTPly8voSGYbpmcIpJC
pj9UJ5m8JahUr1fMUiWfIGdEDtQqA4pe/+3Qz3J/lVvgCA++YEHrETjpQQEhHv2Y
q71RLM1ouI3Opq6ntyixdkvxKN1d4jZl6kW1lq1wDWFQ23zR/k46UJGFjMBJED2A
YdUPxSaS/LpSs4JXL492t+E0eouUy7HRZV6woUVZ7/AjTifYptYAx7rG8kscgwRI
AuQPIBhYOKl7MqUw1ll6uiAWQB1xdkImK554FxqE7b1z4HYz4y1JWz6rNvzhhPx8
Y9FOt+glO3fiu2ybUOHfhayfXnqH7lEvQ25YBtZLDFUK3TkzMqek1uAMtvJ/Hiu5
xxo/MMrMmGRwKSkDlDuRPXAm4BZZzOXWQ0JzWtjJssxdgflck+G8/j/IY+aPzwjH
X7UrjsU7FPyYwZbRzcd4D8tQeEQaTs4PDj9gbc/KDOMaDV/lLci4aHBodljyqr5t
rd4qWjrRA3UrW+pwI2xovjA+wQJgVv4HQ6uOAxBruWsQbJ7d+cnrI7GeSWckB2vJ
//7dwxn20PNVX1DRvYxAVbrGy0KfBKzOd5IHrvmg/c2SChmAPCYpqcN5z1Rj/SJg
49fbAByJNoogFwK2zCjgGemuQ4U6RS4/zTZdfZiriQs4rLl4lii2QAsKoblzjZmh
hV5Ain85l+/yGogIP+oHbYVmXan9mMv4Dx6HSqG5hUz+Xjiv9aORFs9nBsKpaxea
YQtUDRZwqPehkf7FoICgRmsStO7Cm+LQ6Elj+1DvFlpdFOdr8f86g+yVVFtauIcU
kLuRomfScP0x20YhbiCYzkQlaP9mHuUzZK6slDsl3p6Z3HAdJPosfVsplisRx4h+
fb+qp4e5I3adZ44t/esjj1He15B9yaTmYxF814464F/XZ2bBvW+nSCGpOPPvAXuV
OoU+8lbt8dxdY83i/YxdxScgTHToOwaedS3bf4Zn5nNwCnaQAQ7WT7mOhtsDno6V
XgbjwH7VIIS4+0RmOXDza+3POd+LZn3ZR9glwK2EzoXxO+s7MT1iBiGGwX+Mu3E1
JrR7otBA2uSwP7QQlPqOmQ0D/RACsgpfyuCr9yUd1haKgpRhXYJRrjwPP07xDsP4
a6zSTWnhzaJRt3k+ay632Tb412n/mwqC09xTxW7g1xIVl/UbyPe/iCMUw+RCC2K4
S2+kV1/srky+UrmsQSqytT4CHS9GBtPOIR6D5RnYbH9UlgcMUfWo1+3lr1U/2F6k
oeu9/PyeCVZUTaEsSx4zQ2UA/J4U/e53jL4sUhoFiIGBjdzEf1FstzHhjbH1LNH9
Be14HxRruwX+lnF8P2duVrkH+u/kzLCJyGP52Si1uWNsuL5ncIpPK+2VDc44rtqR
c6r3UrQtubgv5A3eAJlmbvm+OraG3fkuTFjI1QLpqCv18F7cneNZSi8NBrNFWewW
yThKibWqvAhk1puFGPwR4SW8apwxPaDx1MC2OF0sT3c2jY5kiRBH5l/fEXWZBDg2
k4dOs6uw85ey4Zy7iTmteDq2AGxmlkeiei/Yllo6B3I1s4R4qm7AXEjDY3V4A7HW
+hKAaaprbHhXlitbmJlgRtsUdCbtoQD3ZvXhlkZyEH2bG4sDa+n6OjjlfHH5Ji2/
LMFcIOcKkTQgaOasywyIkMX2VWvdrcHTrnaVlcoWJlRV+T4Uf9iiK7AUQizRi0rH
kzAunmph8Amkm8N791DMQTxTblJZ46ksXobqrELOJtDQbtw+KvD9Pwaf8VGcQYXa
rNW3CPNBjKd08lVKH1XHJULLklaSnYP/4jlTW2SVMFaAUL2sFYXzP86GcGDk37ST
I9JWy2UCkPZ9IGxXWSuJKhTzA67RZnVrYDNnhvYzmC5J2NEDEgKlvYdoHB4FU4Qa
7Dumy4/+NC8Z9rZSHsQ4Grdfg8o1iniudETwbHVypleXdstGw2QPNFpYReXoqigO
ppOF6U0IlykAF9M+zLcfScJ9kK8enRToHxg0PCVY8PS00CFI76o2zRzjZ8vsfjuI
MlY0hiI36xQvhFXqCS7RWMyDFsxwuu3B5+mRQlQLG90WHdekfPDxJYhHKZutG4YW
qPoFxPuNnrq30I6UriGRSZItGYPi0Bx28fxrB4Cdpos1yCD2xHkWhoHG6w7grclC
K/AcZJSyyGq0ZPmqYH5C1fKy7vhklhpPYkCAFaUwL1jfKOy5AcD+yTm8Zkj98H+Y
pOEoHw4ZpbK9aayGJMpi8Ikl3uLXMRdG6KUXtVt11liAXV7I0FayVCOZ0VMtTBbT
cYKUNQjKjNqGFbB1aNQWfQnLbP37UOhgZhCK1rkBRchLe2FGjicnm8aWqnYKja7V
q/LO1tSAQc11dHgQEib0l4hdHnHMsCGyavPEt79MSm6HBgHJa2wwLr1gJQ8k8Ocx
xnbG4Ksy4c00CizqYB+Y4TiSBgNReidzdFRH9EZa/IePTYsAxWKKjnCiyzUalC6q
FxrXE7y/Xbk2cXAAr44VUqGssuZEv3k1Vd1DwwMP/BsNhHeyFr0vJVoHL4HtD8qY
n5mvHIpGfX7zoyKWD7iGSQLUIeWwuVQy+SemFHeaDbhtoZx9OvFKZ9xvHep7X58M
mJzl/II6E5KZ1m0DnHiZMWFZK+EC0oVW4VfZ12FoDZoPL2UUiPbLiZBIjIjGx2V9
Puu/vDu3ONYwUZMqqf7A6+qJxFoPlHi/2s4l7F1WijrkWAG/fwakA6TokXvVFNnI
UvR493IMGF/fDkb7WrYgzafCNoa5mQpXUXWB+sN+7NsjWdSy0oqzrBVqF4a8buqg
CFDC9g4z/NWwqfHuXG8ybf1WMTPlO0X7g7qJXoB+2Bp6esMKIR622i0zXK84SbhB
DJ5RvBbqJ/bqSFOF8uVwVfsEDVMTmczqI0tueLcsNLXfwYSidy1nh/DBF8ZrpyYG
84tFkrhNNiKNGhb9JTtLhfl3OkAyeKiH0h1LmyHRtWVGgZucVzFEt6vyrYy3HEtg
s9PG7ffI0Jrsxc2DvWj5rOmtdb+VPhWpE6C6JjnigNfqybgvoX1g+sNet+2TT3Ps
nltIsRa2ViLJisKbC+W/t9yDUlqwWFF0UAfklXnZMGs6mQNDaaY4tYtT4dGvIwUp
+kSMpb79J7S+hBVtKP8YLCwQCQHaotiJi59Qaw6HRyku5aze05a5MmWL+660P4IF
hvY74ZjhXYiNE2LM5JbJltWx+CEcOrUzTfaX6WdNnnUMJH/pwxVDUsHPwurn2BC3
ALE5/kSPLvkMs/Fi/zokPNm8Nz7ErtGMkPwkzB3x1/CjtMoZruEx66aZFgxQ+B5b
YD4AvhglXM5rvD3RTn9paFJdeAWVeswzW2o7kvsZmkLVY5gvjD9v6RrceCOvyUDD
thGRfsvOY/YFuRkMO4XoIZVnkHw0VTijMjpDRc76g8Suo7iis/EhDQ6dV4Ly5Onz
+iaS0Rnzi5iqiQK7hELi8ud2SmPVa22IC6cZEC/WdUFbCuI+HfZE3M2ak7/S8Vsk
PposSSl4ZVOb0bFgG970uGP9kUcIerNNrPdmGf/ip8j8n0F6hyubPD+rZTfdF3vg
q+vCNAMyt0P7aYtyZ2F3afAeWhxzIV+LH/6boLZ693UaI5VCPVfRLnOEqS8ABQ28
VILLo0D8s7BK2HGYTXixneETRHusPHo8C81PRwJAsy33Qd2R3mJWwQCYmg89loao
W0YwnbwLExOZQWsnYrWlhjE03dkxy2kE87unYoeLRusFxsn+1DnAygqW0iSghty2
15CGw5bgfsYb1hu63lHldpmKORRkLq+LxVzXqvDoCtm/bURA8z9cKohVugFKuk9V
bqsluRPNPkaFmJASwGlUai7WGOHtZF2OvpiYEvNMS1kTtN1KKQbo7zR07gQkN+yl
L11HADcnCSGctFi7vx1SssoBMcTrzZF5FqhtE1eX5XDJGXCUJMIuELHCBDeXMnhE
KgIvZOvCV6h5nZSmBGTAdzXqw1VZzL36GI+i0IFj7iY/hE1eSxmN1tyF4p0E22YR
RQRilCpquIk9QJJ0JrBs8Ny6PW4PQcbCmfmB2/bKR3BZLADm9LE9U3s3DT0dnbn3
QDmKM3vq344ydaxoxSXLc+xpp/EmL0SbNQuZ3HsGkKv5ah69JGM3O3idgeQgW8LR
ULSmaPfvA7XiwKFTeZ6N9La6ah2ILw4iaSG1Uq3vtlrxCZ3ckvtP/jJpawFiC77z
CSEgmb1m1b1r2zQVGdfTEQtzg0MAJvhvqkZB39t6CuoReZIVk2lwAEmcJpHbYSPM
hVmC3bXiFgMPRuClDcB+HKLFOiTU+DXw0wjOkPwdRmOvfci6SEwzMl4j9kn/uoi7
Z/SoWo6jKiAXVSEMDY4W6YVx/KikU7BerAv7FzFj588cH3nhAgvvsbsTk5zQyRye
7UWnrUpxRrEcIMROXIQG40+6F34844LlpYl23Nbo5DXi7QhC2vHAJOAwFYf9Q6pV
82iibdUHMaTYN6gn1J5zC9Ws/AT7r/c+uIE9TN8Dh/fOMHuey0Ne+jUJQlY8GJwA
xZA13Wms0kIO2QcTdee0+ZLkwsgGLpEew1ZX89I7SwQUrtjxJzYB4K8T3z0Q/Clr
JjLie5UdAX0pVjVmFosPSoFCfPFERvXGCvdDwDD+Yd2YVSRoy0z0Ut8jgLihT7sL
RkSnMszaEl6boWWXI9t4L52ISDo3X+b+E2qUvJ7of9jmns9AqhT79h0tbipMZl1z
L2RGfBuC1HdaN/P0MEUQqTfuw7S8mIwuLZOnnetfVrRYvSRGPVVn3FE3LtY9cpnc
fQx+trvBmjjGiqhDoTQBYuPAeT4x8bJ/fR3c4L/ru3M/UCHl5vI6zZjYc9vPW1et
zB4SM7ZPUIHCEFMiDeOdxls9xE7MBoIW5E/wmR+BD39v/S3g4Z3XwI4KHa9BlDxt
8xhQCHPFcqvM97tW8mwDZ7nunV/QUTXySpTSjFKcw8n83I4c5WHgP/zDCbuv5PjV
TdbZnUGT5txUXH1MuVab9x0HLvFcs+GNl1XEWD4vzZDJZcDbghQpldo0kzWA96vo
HBEnKgBeJZT3pQIlnh7FVkbfoht+4izof5qAfY1gTyqhz4k6brq4t2L0nYbMMNoa
o8TfhVlr5JLUqfJRXgFjNpoLPxd4/tdHsWWuzPuVIeXRiCImXk1XzsdAysDbuWZd
jWGU74OpfAY8v4KKIv6fmEEnZ2VWDSOs5CAoto3noihNEzM2Tm35XRtc+Eq0MstQ
FXHnn5NKJh3M4/l2gwlyphKBMZbI9s7m9VE1ZzAQ2rkSkhNI3UG9cqeZffPFOuy+
S+yPXgG8HMbyneSN+X4p/ZfUlYYNrmlYprajwosHKkYef4EkdodfxuTLzrxq5ZsT
3uoql4H9uo9l2mlrDJkK5Fg/lD9Eu4gwcKq2aRIHLl8QGznADhfCWUys24mEiowo
H/6pb7DwSElSUkpTC4jSCb1czDUmlrM9IMww5lDpjWJX3LBb0yYda1yGl89mPUx7
oXig8GJ/AxOOOvTj4ONxt09d7Q4Mro/ijB0zn2bo9quBvT2u547Cy1MKJCqY16mm
6VEq8ONE4JeDFLgM85javmNYFfJhaSRGyVNvyjwbSaJO7jdYgrUijtEciV/1/8o8
xIcNZI9fbeJY4HdLjvlPaTRpq64jB8bEqtKrpu+qsbXr829mgCbs8c/nLuA9gDDL
M9PLmUVWXy9OttVYKBD4Abw/E0to79j2JIClOm1HFZtJybPcIzCwA7jBT2jwcpef
9yzaZs7cQsYu253Ht4TVQ/mrnfBCloene8yJe2Fj3c6SqHZULNc+j3RTc/bryMWM
I3UilgwwZK+JZkLddIq9xhai2ohfVLpMxjUlsSNiMK7RAeHdM9V2ba7p7YlK0W/H
Gis0LKpZR2uYFhF8SS87xsEkwFE6YxxVj49kQllqlmuzGN1buP/QuaQdL6h1ofJm
4AkURTFClNHT22rzqCPaBaRAFfHLUzwOq1AFc3MICtLfwkr/o/pBiK3qw3tVQcBo
o/3gvU0JFh8l8ZAz7ScxwaQePdcv/uVxyv4xXp2Tr7yM4bKZEAz/khwDlnr7WFuL
YQLadMJ7S0RmjBox04TPrm49uHLY7Hu6W0yFrmrGGu5k2MFKute5fQPLfH8zyIDz
OY5XRgCbRbY4hxfwoywe4haoimSn+EHUYLQ9SJUKwd0rnYLljbSRnly15+48IXVx
4ydK7SDd4HmjNlHyYr+mlocPupwy+WhAnTnJRUNBjV6Nu2XQrtkKGjZv8p8//TZk
RQ8CG7SvYpgVsPMRccImqoTJnv2heC49XOSXUj6HH4Jmv4klDCBzNTLfIo1SArk5
hbAQrfs7GLNKvzVmMI1kkm8yNfuaS8WuzSss3b+CuxOJCzoMLnCeXmD+2Pp039ch
EGEQ+WtJ9LM40o9yHHfBs9FK9G/7cSkBuf37UBZtNbhw/ICwdp2xhctmV+Pfrtiq
Y8ArGqtqZKlLRvNl127Zg0iKquhsfisKGbn7uO/gzbd4eIUqkS+KhPLJ9LarHjn4
xZwlfB2s9sa/n/LVBGvqmaW/UR7WG0QDz5qS9s2ESxX9KqbtYZfSnMHNHByRYn1Q
7V8/J8Flq3VMUK51mCtBWWQlXu9lLOx0ERCbs2gwcJyvv0ej7ObsfOiHniERTJPm
3r6MnEVtjU1dB1GwNMt5/VrLkUEo6O10jT1Pw9fJTI4ZqtMtgsbFYHLcS0R2Ktx5
p0ZVQZWbfF6J6Zt4GgjKwLH3+CNvsRFsob08sDnQKoHjQYHAqlDWcgrLhZOT7awp
c1p5/SlcsgosGNpDypjqDy+tfs05j6/9jKOWw7spt3fLd5jhnKOgE4cXcb+5RNZV
X6a3y1zG6jHsFkF9XNsGPb8L3ObppjwISKSui15LEWqFFWMT/CyeqkyWkmJXfOpS
sKi+j8vzgxLd7bHuT6uYAz9FA/JEGuHrrdl8YbluTkGjlQs7RDxO6crprHihsZ+O
K/6TRfSXA1Ipii5j24joQbCSqbQDtg5mq0Get5twXFT+LUJEtRUff6z2G7pPSPKj
/yU0gQq0BsvNoFeo4jTczv8KKLK3hDM62WckBP1UXMrEu4/73UQEIymB3ooGaNs4
XTC1rRqujS5MM8zV/h5OnaLBkkfklKv3NuNQCOwVgvwOpUswpGkMQXlLLkYDrtXW
CPNEfcdtRgs/zwtqeE/bzBE2oZaZ8++ZW+nMpvtx7KUniuNv1sclfTWBwiq3UsGo
Kj3XK4seL3/v7697rCDi0M10O+ztH1s4O+zqfwI1Dxx4EZKyLJdNo69NDAylcsPU
Y/yBBpDO7qWbzXvD4hglusvIy8OQ+NVqD5dJPGqGujKi8LOrWHLhuLrHJgVDdqMP
c8Ct8IcTVwpmeUXdaJFrTEKD1lFNR0Cd75Y7nhdYclwpKC+vIhofrDA3a3JXJZDT
D51EU2DSPIJB/H28J55q5uIHEBTXXMAU0HwiYeM9VSaue52PnzajEUk484zkPeSh
VpTVavgR/r4HvcX5qY6JxvHRzGFzXOfxmWbgoAsReYm8t800/vRRft7FVwpR0pQc
/ejLdDi8uzq/AvyADb1cFerqk0jN3KlFNl37sSqZQvy3tByezqnqUy7phl7XMj2d
STY9dYTWg7I5ssp7GPomfYXMCSUMv1S48xM5yfbTB6ErK/n0rp7ICGTzySk4L2C8
rfFt7JUfAGBO77vCOWzrfTiHe9/2y3Dp0SvtDo0DkUwbnx15ynLDK0IiuUGdbwpP
UTLl+vH1x/BB9SyfG8WQDyigqWeLPhlG0ym0MVAci2QPOlVcHDUF2vr625kLvq+G
Aebaj25D+G9k8w70hQmRg1zlSQsEAicuty0V0szdu74+1XxT63CZLnIF8BBxpKYs
aR2JhE8jhLzCCyK/tqRWTY5LqO9StqBcKIZWZ9JyllUMzsbyC9e5fvKXEtV6cKz1
FQJI7/mac5f/ZYbzmGWaS7UVY/YVnBcfZH9LPMIgI73UB5MLW5m9onB67JEAZQQ6
3PArjOqoRu7dBTygnjrJCOK8nXDq6M6yMuQ7i2z3U06iorV3cqYGyg0Q2CtGCyQZ
yW7VUQaXsoWhEF5zZ/9l7ugpFOoRYXZPM3a9eNnpS/scH8wXfpxBJ2Iq9j2y5Ybn
fiDFz/ZOg6lIiYRnIXgZ7YDtLRh9hNrqHPWcWHNiStWHIr6WfVswcDWguzN2/ePx
HP3gNR9PwxCpVJlD7ye+6xBvqaS6RejnbhqBzKa8onACfPjFztho+tbionHk1s8a
RliW2JUrhRMzs1wE6+Uf2vuYEJ3d/ZQCVtM0QswSJly0wol1G3fymTuMOY3/SzXh
0dxZDEae3gBW71a2v38iH5ArKHSRUyYUYBvA+epoVhIBHeZWL/zZ/7cLoI0gnOcY
4sg4PUN53HgrnrpZTk+2Nk9asZ6Yv5+OqEbZ696t4eJuiYeShuz4rMnZQ8RekfO4
V+hFDVyIDyz8w0nnDCfZK/ItScpQ8LFA6yrhotC2dAg5156yh5GG546EZuOrOQS8
lxXxtpJQDzuAvhnCZi2X4wKaEW8LQQaDf2nbZY3LoK4t00AXrUrfUQZKwSz1YAEu
oqxawHvmjE6tk/vEVZgrTnB38FMP31G7T08B2E/X+6+oRCMtR7S6a3LtIDJuWvym
ye2b4ofO81TVWCwC6/axc2KByb1IEJIzCBxto5xVTsL4/W4VkVZNhEmwMz43KRvT
aXU0o9p9cCNZVoKfxrlqGqubUwYDz/GB/GktkFxTWp05mcmV0RjjQGWjjp4cQVci
Edxe7deVeYW/BFK7YrkBw23ZF9wzzNRG9VymJ0e/DvFYJN2XtjFaZasF0IfpCwCT
0ve2vCPrlRvZWZ68oYU/DP+J1bcItm152Se7KYg/65tJJuLQYfqgDjyPha2JwtPB
u8pxiXAvjI/LFw4nBE19HpwdsMiyJbI5/QrW+aHqeb6UQL4hNYMouYwGQ2zLahLN
JoIZmiCP6i77vASrM2rQVR4UZvOZJiD26Xn+EyLJFQEw+bGzLulJc5/mQfgg+i4C
bYgdFSnbQysQOeZrve7ude8flhVwoYcl9I48snfrOu/tNA6QbWnTloNxaoRwBeo7
QyrKKq0pJ6oaY58e5CPeqPANuWt4ql56jXjzBOmWShssLfQbbdEw7agLkJ4vwe6D
pny7UJFpLtJUfxX4cV3tvOZ8SBxZAD/UFx/IopxJTTXcQhA37+QSl+L9ZmIOP31a
RL0XhOmsLEZ3659LF0baHXxBPksPyoYPEajWzY6yvERmqpI9jXL7Z7M2rJ1CT6wk
v98fRtD2HDHuTLvBmtesz7Wf+a9B8dUBqvAMmHmqJVtidPSAbMzmOfzCa+UTCNYq
ufFZ9/nTRyTNkYjgi6skhj6yl0WSz2xhhyK41EFi9FYmiRceCQpTCBoOU/6oGRga
TLmxTOs7Y3tGppEVuoJwzgeNbgEeqB5D2s4D1+B/a+jDHoa1KsSs4buJKfvUzMA7
UCoBe32CP8zGoHU8SOumlbQ4V/GMAjCeWUYu+BLGiI1xN8j5BF0PZdv/7+O1U71K
H1GrO7JmZx9lKRcPwWYdbIZ2YntYy6cSWx0+NuFt/I24Cbtl7DnvZETKqPcd42O1
6J1frAILHu3FDg5ytKu8SLiuWzOmco/DJ2Xs+lg69J4cmgVCtz6MI4M4abMnzIsC
nqX6tkrFJh4Wqg7wE5SV2BULVARsthpmFHLjz8gKAKGqJpSsgSt/KrTuVm7OGw1m
EkJdRH7RTmQW67iE1nZbVhj+BDGiiTfl2gU8is/oh9XuEwNgoBjeNVJ/gCxb5Qns
c7K6n6QT/XY6hClm1nN0NczxYWNf05CwjaSFuIZ14LHXBHD8GFfJT6rqMUDD2iah
TDdaJ/4g8y/OT7fyBPhQEebGJZ5U9bJrKwsUultecYnQRgRiI95a6Jcr4u+QA+aU
oi05EvxuFXYv+K1Um1eDrlD0Ua5qO2hTzZBuS4nB6SFx91v2zZQjOHTBkfVyDBlk
KEFlHSEaDvKrQsIUgjAjgTsop/xiUH6pEGeHy5i05OxMvllSwXDld4LFO+fznJmn
IB+50A9rCWjBhUkmVpuhSSNFWa5nVicU7QDWO0HGsRZ+YFaCMuNGFAuHFhQJWswL
4oJ+bKij/ms7YOAgd9afXY2dZv4jmmZyqOfgWBn7qzgiAB5W1t7zE7rbtO6zrVH0
cznM5Ij7z2TVwol6KtGvrvu4X8P18uv+g4DUHztQajX/gzzWdt9fcsvG9ZXGntkH
DP1AeJSRpnsxAd+hqHVou6tkUcvj/hq/M7WujVa2t+b9cmZ/S+plT6uoD3R56jRj
phN1723yAcY+o6z7wh5Cdf4skUNaLHkr0dEy3xugzyMPir5xk8ndEKQ0J5LktiJX
XHPdLfwPV8AC7RZXidt64eCv5nXwW+4yLXJK82HfVgr6rqzFZIvtQ9wKbqTYg3cm
vzOlM8zdZux33wd5J5lL7C8vJ+7mpKdukWDsLFSerxnDI9mBiWYEg7Jbt/APXE0c
E2F41zR4TUzSj/t1Tsg8a205MHFbTDXUAcyPs/vh/BQC7cPQvGkP38IJCZF3woc4
CrP4l5Ku96kfrzFeWE0mjwubzaLCdQ/YR8CkqzSY7vb8Oargquu+oljJDGYOI7HT
QWoOnKwGQK9c6es2MvnYnyp0DWxXJKpqxRWbe79YyZQ3akJ65+ObKeABnWiM7yRS
4jBbPzpCFM/Hx3mj/qFr0twXNJi6V6XutNK0prKsHT0d44+HGYZjq8YAr4m85qGX
r7+EWzSVUEFFSZ0b2D/hr7OClK3mRNRoLyIqSrtOWOVyoEeFDr/3JML5hF7uiaB/
Cq4e7yy6cvaB6F72BL3H2apDvQaeii7xi6Y/wu507T2FqBERm78LeSt4yyb9/tL/
mj1Dg9gF44nG/teZZOab8mRKd8x6Omuoi1u4DIiEEjl30KjEb071eoVS6Sq0RmSa
PP1Xf7QGZiuLmrkSY8YjR4m4YQl4TMZsRx1B8zqsCiOWA5Bh3D9mu5uF/mhC1yFk
YRIkM1aLAmVbSUjv5CXW9T/EIZQxYLUrCeT3pX6Axoa3K1UwGJOL45DdOeDMHCZ8
2BSAZ1tszbOiKULa7L2yQOC0WXGNVIRUnswTB5IIhKgWNsd3k/Jc7y5lkBROwQ5M
by0fOkPgbEaWJfhhOTN+GbLfAtrM7lNPJHM2EedZFuyISYg0eHbYMTrdLuyVtBkJ
JzoaCCCj/AIMBtlx+Sqx7Gn6qxLih/++Gx6di0qJ83SH7m39/5Ytw7Tsag9uKEVF
q29j/ogG1TTHYgFH1WHkDsi/el4PdBFQvg/uH5vzFfJBw8hDclId4RjFshqHlqBl
NiURUdNCYnit2bkoXIPvQFrjUCqe4HWvjf6rROUR168b82t9ZaSZEVyKbHUTbtng
vTd7MBt7+JySgGz5icpH2qtDveSyJPzjjV6joQfhtgKhEcVzU+uzuIL/7wIrRQp2
VP4kJ8NgkPtrKAVm4aNaGg9YR2kedQYF6Nq58zGnmU8U96YxoDZuZaNwUZq6mB4W
1JRF6K8AO4Bsd9Syf4Ga1Bz33kGLOrSn9j/FiUscxftt9Kor+AQNevd34GmoWtYE
lZhbacl+nl4F099qJUwhEEzVxgsVjX4jSmuxBl3T6YHJvgvJsvzFWo1jSvZE5eUA
N0LREJyLgjWTYoRVBtMJ3LrwiFaTxKFExpUwlhzzmnzLf8/zHk5xsF4K+jTLfMdx
Rjq8PTqm4iGTV3XZgp70N41d4xFgPDKnq4h0rvaTEGhfAxaGBUcOOsnOBywy+L3P
aU7+VlDumC8TBQxU2vRTCWBRt16AxEdfaAd5/Zb6yq6W6PZIrs87UIctGejti2Af
/d6LsdajSe9D8pKYJdPPsfD6lF473XoZKXSTVGULMjeNhRLpv72l6JE+uBpavuiW
TkSkflpAJpUVcFGINVIn21J7z4atQ1p2vcpr8btvKgB3Id8PM7wFaUwO4IW45RQM
V8z1NepClNw0gTVBwaS8kAZA9lsg6zYcthTA34HJbOuLYy9XPpkQZm7/F+fwrP6m
jFZZKmISo70JGNWFNt5f9T6daI1kt7CuuBPgWUg35M0N8U9vum/RDVqjbacGp86e
AwJDCuepEfutHwZBje7bpWfgGT4tm1N7QChJD1t/4H0lQ8T+n7xftf944XZxxKY9
if862KDkI9dF91SgcIx9MQhpWuoiISXycQiWC7WYGos+CpDmAuXH8ulMdh3WCQmR
ozn2U+XryFih9carteSI0NOiYI7SM7LyG/V6KC+LeXUUMuQj4+5eg9W1QrkclwO/
YdgJs/4dwOFiVwIymVMOHoBxUhGRRFEKMlVwy0Jgxq+S2gsPrtO6ey/GCw+XjlMR
9R1OmYBIlBsrZRIs4MTX+MaSFJNY2B+rWYrGStalbjM/VVrATL+WP8Ra/oNFvlua
64oD4PwBNAKRo2J4FpxlqNkdJWHgaOPG4QSx9sndMRsaXlY5Nbj1n3c939B251Q1
TrUAp2wVYuY21O+1z3oWsie0JddvFnJXYkq0E4QyD6bP3ZcyBGY/qiInHSyOplih
S+X6jjdZonaDzF9X2/uzkfvJ5l2vzHWrEmyHjjJ5/Nzq07kCkbhSzMvJwa5WntVm
sUQrBn1sJDFGAkiWQvKaeOR9zNl6BAlteeqCfipr5XTAK4ofg4tCbSs76iLSv+3E
E/VhJv/TU5vymWuZXVOD2mgKDSBKTcpVn+AocrWFyL/RQdneYacP7cORGRfsEjps
CLb+nDccg20lgOsQpqoMwg/OYPjs/Comto7q31Zv0y/15q0NB4+DDcms2OC4fsn/
0LEBuWOOvsoItGG5qb3lasHWz1ASZUOuXr221kmYcbJw6rkgBrqBqoJNt9McWh1O
4AfVOUuo7E2NDhXEfvpLQokMLyfci0kwv3zZNy/vHn6gCp7QbejQzs5UvmiW0Wpn
6Ev04Qy4My1GONrNFRylAYJcdu7YDD2TMkQf0yCGV4f5RfjVCfVz1N2TIWmVcEXy
zX/ZvLtcHNBDd/VUmo67f8eT4DnYKoU8DpIMnYKtFtq5hDZQ3dJglBbdQlYXV6kt
HuoDFQi/HEtIP36JWA1O4xJ7Ep+IMPtbTS54y+pFqhIk5BG7g47nfNkN0OASs0bL
t+GIppq6L0t1Ho1VhVaG8o1zEGFAm3hcK6j84YItz8QFn6JQN8QwYl5xMCM6DTt8
PWMHB1FPkjQA3usuEvp7DY1WT4KN6DTGThEX2rynj45AP5uoxUP1iznRIyZAKKOf
oNCBy39TG8/nU9mthxE1chmKijZ65SE4bxW3xXFN5ya/QDJY7qvX4Rm44oj0PWyD
jksT/b5WFhwrAAR4c6eDnk0AJ0Tx6q9khiMSlwUmVPDhr6oD6Lw63ulUAf2aRhR1
dd6b/yxpEo7Jd7BbX2eDVPwK2QKB9fPGbFHvWYG6vrgPzZpnokQ7Sx7sxL5DnVuK
HOnAOe50racojooEMxEUqQJhmNiPz+9xHvgIhh7jWEbIn+Koy7CRDdZzCsTE+8M9
QFhGB22RNtnU20njVi1mphWgAqKsaf5aqHSdlBLoF0jf5bIVUjtKcx0l6zaRWTST
X5fe3ecy9UGSJ+G6PR7PAIBe9YJSGoFM3B5DVTe8ObXmK3rf7Ctz9x7HxxjwqKea
CwWkdDfRypZDX208Pdb13KMPKmQfXm9Ex6VE04bYdq7k0kqiElWnWYmSaA/52R2m
G3VC8GIUSe/rsMJCXjk0/RTq+FYD+IWk0gwAQsdpgYOUUh4pFEeE8hsT/K7Ls6LU
zByUySj7xzbuj5LGwUeHLA2yH5FzKD59f/Aw8U7c+KfAps35D7yKr66D1R+hmKoh
rGY38EXdgRepHj6ZxZ9lMV7iNUqSQuXqaWiHdWqh2VZlCGZK1JasFmZUmffDzFJf
cfohu7zcRLGtf4KCxoF/SIZXIoZ3drnlmtuwAP351GzmSQK5F+ENA6SZidfoeG7Q
azB0AfcPS/jmmrRZ4dGjZT2Q/WSEegPolTOJ/CEaGu5sbcxqTIWwvND9NK8Ihz4m
UPD0niocNfTyTIxUPlU62zz65KSjK/TIr/3hZ2btCQZoGenPRn5AiXz0cNQ2iKuy
4VCmxWx7BAzQh7FJBuZj8P3Ib8jOxKlVBMHgNdnpGgN9LK63S52LaXPglanbKlRg
QjOPws8vZX7t3gkb0gzd2mDgUsQ2TaC6jS3WVtDTsZtLgLcY/hkCaZtJb0yQOxBH
KniU050ypQaU9J9maK/6o0Iq37QJvOP++GdGy42RYH3nRsP4jhEIarEuJhp+D4mW
lb6Gz8xcpgBj1Ltnt/hBsc/UUPSB2bfAQI/NhrAANWA7K+IRZvyljg0RX4mR5V+V
8ce+P+mz/MUo0p+dNVVG/teeEjB1BUG4taRsJWhS5ads0WgQRc04oTbxHTL/Df2n
rF/0fnt5t4ZcJyVaMeHwdu+Q/b0xVhtFkIbrvdGooMuSeNwaKvau7oMg8SvW5gSm
HuluMK7DuamVag5S3Aa72vJOLtWG7jBdfTrbjTR4G9QTHKj1ItFfMyYY08Qz6quX
7t2KoQWUIZGc6HKnVOroYAht5+jtm43+wugN7kqK0zkHe6IImUtrEnVkRQ+D6lUZ
wDBbXOTvFQy/42/TeCKSMmryakkMIlu0KXOncc+JX9Dd6aCIovYZZpUM2+tpJkFS
eJu5zh68ZotPTxuxn29dhEO7kGI5FVnVMJX1xMjpIucoX1Go7rVv3Y1jYuLqbHcC
9wYdPnQFuqeZivj++rmU3QpcO3OoEfn75kOit4/4KduTndy/PKQybBPySpT1xmcs
ycftle0NfiQYXv6cWcD3yB8fCtgavq0Ft/6d2lRW0LXwpfdaZQcc+Kq8V0/WpSpx
2hlZzGQsfFbhTwQwAtW598wxwrP7qRaWNXIhDS0++csh0lSzpgtiRX4Wxc35PsL6
0yJ32waAyWDCQINLMTS1iYigo+zK8gYk1bCEiS4FqDb6wPXDHst1P8k80gSu5/nd
U0g4EC50l58pf23n2j25XIR1ToZd+dOEgbapPyrfj2JFqxZukzZjhAGVfPO8Sy8W
BfpH8sBcJFWk2++1Hhrnx2T/vogtFHcKbwoq0MYNP32Dz75b5PS/uO6CRYh+YnMo
vo2LvXRufnX3IzVwS6XBxKwg/eYPCXXhb5OmHNnAJu713VtqC3vZxINc9llfcYMf
xkmqQTcoCT+YwemNNRSwbr6DBue0HYzq2Gg/RNdOhJunxhej6VW0qFfniABV+2uL
8CnKA9v98GkaA3uOmtVcUMJuIzuUEeGDPLueyABghXHXoCNO0iNukBBG1Kc9M6rn
6Rm/KzrS1x5NRkAGosswmGHnidmrl3+FsUn2sIzzvqfBB7ZAjpFYkUbARdGlC7KA
9cszbG09CY3bTwUR1NKsJFm3Axm4BalVronM7edHz47HvhDVdfTYB9vQm+lkEpcL
QbPW8VNLrnQ0uOMJyOmV2V7SAdrW1fagtiuCLPFZYGWKU1mA9+djr1sVrC0LQoMP
wU6Q0Y5QN8AtSjFhTPqG3PvqjNF3JU9W7F1LQSUnFROSye268Z/Iw/E/FjT0SShw
OMN0KxZ46QLT9t46vLwig1pkpDxAlmkln9TxRpBiSf0+sMklPt4BOhe1cGJDoYRQ
Ocaidh7HdkFZwUxQV8ABM8KepWbeMpiiBJiO/U4+mtCJPGeC6eNiM0m0pwWRMHlv
XIo4ooOkZY5e9b0yMuv3G5M0L/kT5ir54BM70NYlXufVJRx+qPc32QcLZvkc95fZ
NPzFjL0QfTbRdI5wJ4JaO2xahzCmhBRfluzkkPc6ed2NfyrC7xIgA/RJGJzf8FvQ
A3fcB8twNGT/N4JNJaGOVohsLTLYpvZ+V2RPk1x7kMu1AuwNW4ks89hN60jqinQ6
xDlQCpydVIum65miOeVhwTqJpScWwpux2kvCho7mMpnwTqooodxSKEMEO0mVghxC
Uh122zi2Vn5QzHzMq8yKUYhiUk4wgktldKZ3fLm3TWQYoM8WwVQNDRyoc0Aoa4ak
vruTRpqSekOp+sX9wXuM6jbWXFBxH9YgK3Kvm51Wu6KeVCd5wBMSHXwMLaTFxOPR
G7nU9MEL9cvFeM3rMFQ8KcF7+kkHXtXSiK0w/Mb2SdZLn21B578S1+4/JYyhT1K/
hKN4sRQ99yRbPf7b7l/8GPpWnwD1rENANk9Sm8dG15C2LgNBRWRHCW0iXESccXYK
7mX9qdeioEcGnbpAuf+VMKs3mjG85jyqQiWWtOqxdr4gmjS+gFD6AnwNmfiCH73M
WrdCm5H3MLBupozeT1+gGjcsgzHFUMH0+XypIzSFFO7+/nR9kvZGpHp0+31Y8IyK
zA5fIOiYk4uETRXac3uFWyG2p1YtII9jJ8/4O4bMhDdiHxqLS7KPcGNuHMWgz6G6
92YdLPCv8BYPmhtXsBHqGMvN8iFMh+sSE9PZoT+Re42tWR7+0tghG/fuQmPA46i5
hE6JvvpXYWImQbG+cy++4isY5zcxhFnss3zKZ1HcjAumOTTvPbd2+ZSMTn/CR62/
DdzbfPtn/c70hdjBNYtUYXIQRbO4Tw0QTSxM0GtcttOO/CcnynV/GGGrO9J7eNep
6C9ibYu8JL8iEaI1pnVkMX5xaDR48tTLp0Ei3SsPRcgj5dRMkedW76LBsS6ru42q
04DeRcBFfx9YbHI7uMizjKZpbGgtDHKdRnf9s9QLXGMK8yLGNQJTwGksprd+CMR8
6JiJCUs6CL+Fll8qL/iYQgTl/lsUBMvQWqC8lzqY0sPHtVQoBNCVPZtrZ8TVmZ26
sNcBtGMIjI7Cn5DDC4XyxKWZJCol7JxxdtxrXtIFkIwCqoLIt0kURsdCZ88O63h0
yVG0g2EUojaqHXnU9XCbwcKeDQLVnX2sRzQjgEfREDY0kpmE2YSemQgYGA9n5qty
AJX91e2ElfHijU4UnbapnXHQFWipLPAgmWyBS0a+Vyzhey93xceJe0tzvBL9LE8g
x2yVXmn6ym6v5d87TDRLWnpNdV9/0/xO2oOedPgfL/x1VCnlfCGSFJZv0CKOZTU0
gle4/M/lxNVqojvB62UXOAKeeHuM4JePJmJvgYg+2VPmoWv7ZXVr5vEK9RP1xTFo
j27XPoXJ44svW5fww6lkGlY5qKytNodce5bfKTUFZM1yZABmhTR25JBkg4D29JVH
A7Sk1XfS2m7+KHi0nvnBDUGyfJpMr8yO1Py3/obQRhYt9V7cY61RBk5zlzKg7X9T
ogwVAApcVsYb0oQG3Kw/QihNpM33aJbNiMFau4CZnvhxI81FigCztgF4oq7Y+fAr
zzj6vEpp7PbhbXtI+Hlpxj1ANOB33o9Lsx491LSD+21w4tDygGaihydhHpERCTDW
Ig/vsXvH7fMVM+Ugeqo6S9o9l+h8bStxhHendenyp8dByHNXshlQIECC4RcikKGx
mMNHt8e9CUwVELOQnkN7PvIwp1Xhoq+uFWuVrCsLct0XWX5ZuOy7pauEsQ+vAzyC
aDzC65usmD44yqdq8kSRA/BXna/6yjtgHGwfIODIQAOiwVEK6eZQYE42+ink10kq
+R1RQ6weXMKqxvQ/ZFSD9Mb5Zl8r62GluGHqK4ghF77zhHEkTzYeWznl1zHZU/Nk
oEPWLMroCNvRGclYjIdHB/qcJu1cau31qRD1koKdkLSkHA7oHexfkCjlpgV84rN5
Og0ZLlVZ7bh07JyKoaH5VygIAO63TDiEwYplPdlKn1w9A9Uj7A46r/v8B+KftkAG
vkDlrw/mgyuOMWwAC+GDa+OX7SqLo3u23YXqs3gvspNPN5zQq4pgCQrVWi4pWLjG
9w5drjiJKHV8K1tTs4aRfPSb1cNPWeQD76ZGnG3Vy+z0WapcgiLd+EzCZfHSa7NK
5H8G86dSdLGhUOhRAXrtJjRXIqk7s/BjHJGiKS6pt8gUpeoJ5dz8dDzRSxaPAyqu
n/wZFTvkSTABy47ae2Nspq/dHikqxo0f2A4HQCUX8B1nr3AUiPvL6WT0WQ1pMnEn
33DCNONu+DjaYjAPvoxtdAVCtgQyT5FXByrD8jJWZzUlWae7WuBRWzC4rO4vx104
8VZ58XGDqXWMNxqShxhsYVjjiIuUXKe5Hk1QZ+H/rCLWALzhvoeMAWRcdquNcCak
bizxv1+7286Xu6nZhhIqRw6a+r+oKA6nHFdvTj+tm2ejZcNK78cdbSgXo0OruImt
K1px/Y/zP/WS5PQqiaOBHghv5Ov837vEd6oipqGJbM2Lz+RtpP3nT7qaVq8kV++f
BWrCFfSB7jGdo6bXjXs7xxolUYnQveMTfVHCkk8/bw67QP9cMDuujv34KusgsVda
JcLngshhQHMIcV9cqicZ88GZkPRvOaP+jKK7p/Sk3bKIBmA7sKNrIt69YO8TPQPM
s5LHeo2CwpsTO6r3PsB75vQBEntAFhNHP4VM+/ERePiZVn1wILeldT5iWqCNsgB6
lX214NdO138BWxY7EglOl6eCYcCeUZxaxtpibxfm6lYT+jOkNshdxkjtkIieLykV
v2Oh4x5FsgdEQ5tlPoPqci1sxz5rdf4Kib95aEgnxRgfTe19Y3vZ4Am2pRgCbu1b
YHkttBF4gevukjkqlfmOHHrvdtcZKzra9BM9dfXOjQ91RwhvbwsC1pw3aizLNAm2
Obyc/w+XsVwwvhYKZBcPJt2ARHOxaoTibu01rjrj/CAzDfdyt9wR9BzW7L19/LtS
GA4zo69LUmWkX703+fv9S/6C0M+ain2H1IG00N2oPlSYX444bCIEDImLEX/svVOy
SHwtgs7PmLrsFdf9Mf0ajvacNlRcxz+V2IkadXMOzM4h5D9UFp2q72psRVZdH3eD
aOBaZd+6lRM2obdYQW7ytKPS5VeZ92W6Eg7XB3qGuivEXpzxHdNJq0EQ0ix4JoUT
pB8RnWiRjHTviL6A0NW9QInOtIMG7xqWUyTjYauKcY+mvIaWBt4bZhBQRwA5jSTi
jim9bTht2y23dPs10NnS7UucDBT2QW2RiZcLxi+ePnPBPE+So8gNVFK+Na67enBW
8vPBL2RrvWqgnWSZO7hK+O9Wl1q7POKL+Vs4fpqD9xtjT7WIrgAVN+eqisVApp/c
fHvCV/LjWIwlLpPsX7vzXuPHCMmvGl5B8LJZwDalFxJgGS0g4MkLFYaCSSW1cHWv
qCn8MTVWIvqX62cKW8wRFMhtPWfAJ7Iwwnokq44CjhpvA83b5O2GqlZn/yxiXVTH
aIvhLz7hEK89FETp6Bu5yXkhla4IHaDAfXKTjx6SdIRmJjewnBr0AQwirEnt36qd
TvsxQSQCs/n7MIBfH2HjiwB4Izbj0ojTh2AJf9msucM37wStha9Jo5lDyvS7vKBP
fmUaq96+O+wJ1IdPAVD6Z9YI34FJxfS4keFZOw4Ay6PJl8yurm5C58OsDY3EjTu0
c7L+tKPovdLmjFZA49RPGJpd3CYXoj6AdT7gig6RMEfzkPMqKNX3S2ltP+/YITg1
uGKsEI70GFwCtQNOtJlj2Q64iafgUvAuzUa4kpzSK2nvaHZ63gFq7fqGlfORPtL5
23KmlL6+pKZjUYE/J6Y1wvo8Mo8AQ8OwkVzZzKwTJe9c8goVJ3F4KDSLq+0QWmKY
0b3pbkO7OxNE9lzEZM7d6pNNnxwMZquC72kpu9hSsm82q5cKqX7qLonVkpXYfTAr
2V0GYPya+5ZtBPGcgQxLugXZsk723zOKQxeLKAY5bWCHvAGFzcMvCO2YujNfoFmj
VCqxKr5HV+1FWWK6GAszo+AGqR8i3S6yPzeGmT1BC/dOLv2n0Dufdg2nCeYcM5GU
HEX6qbcuaLzqnYYQqxqVcFv5t7DAovdrGTbEGF0p+vp9USgyVGWEC7cIpLzL0Cq9
TI5yOIZyXQAwcRmL/sMN8avXU+fejwth40NoWRhXwAQQG/rmJxxsCOCpi6Y7v2Xh
Pr1cNlrESxoEzosTSCcS35L/qV+wxfqz7EwtM1DmcZpExTQ9rQSXsPSFIt+fsaO8
nZLV9zbLH8OkVabycTycQc42UVYrKD3Oa57HVgC5iOceYOjrE/+B1i3f9K2bSvP1
4eWuuSm1+WxWQdYnpwEfMgEqJGJ2WyG/jwVqJL+qTQnHnm5FMozCGXQw2J4EdrLw
VZcxeM6bIlNanxzpKgG8ZKVcNtRuArvpXusx0KdudD1QFPyVTAuDOLcf2SaJMSZa
7E22KzBmFz3xPj3/B3Sp2D00wxkg7d92u/HrOqwtR0QKH3MjAmU2M+ZTbJoGWuOO
Oxsdo+Nhuc355BBaykIaT3QL3tT8bWu0Rapt8Ve0r84tq1r7QV/+mbLEmyB46Xdy
zKwjz81hdRM2Hh3qVbPjFS8Coz4TCpHSu3ydCdpWhuWCvRcw/3d5s0PZc2plw8E6
PR6rhhcdzlGrt0A4R5+oVeqeaDAJ1lGE7ZBdCTOeYF8rfp8fXuJcaGK+1ZuhFMjB
E2apBrPdLXr/9H58zFip5BqzqyrEMLUtzk6+6u1TZwXeqN2gqhMPVLWWKkhI7UEp
elzutZXM7/JtG9IBLYywo2I5zggZUoe7DjDS3pn2SI3nzciagtYoeq/Sc6QwWe6U
gQUIdijdQlRIm4pDJrbcf9vG3ATKL5WQ08mWosZihJFdGOkb4YwlGeEl9FDMYp5q
fB1UMzCBQWEvM4SU950N6CNgKM+wQfBNnnKSRLBEC14Nuex2e9LW1nNYkXd4NEg/
1HbIHNKgvo5bJOm4/OgL3bDaFJ2ZwWIwaG0UO8Jh0xCtopTp5ovU4X/OhWD+kI7/
xrrKOoQo2Fl0OUu/afYf+vYQegr8MrGo5oiYmFglkWC/yEBkycBfboaldPJNjGbP
2AuRfxXj5dhWSFOMdWqWdZa2fe7/VxfsMjic+nPlqWwjKDO/tP/b2ZACJWmZ6Gpr
JoQsgn1hGWTGH1hhwcE3yVd8UDdT1pOy2cX0pLfOC4ymCdWZcAckGB5PMvDIi/iY
S+vSBeEIFxZVymgP/pIbNrcrr5OxusrEseIneDua/n7QMQ+jKy7zcYwO+DFZxc0j
VpdJGqykZgJnweh3wNi+q3s5MF1Z1fX3D+Um8xTE6aEl6h05BClHF4c1RfM7VSR9
7RPWseEr8VSVzGYEmm/vDmALK1RATDlj22gVSKKJeSitE2eBGzqMZPGr17vzidHB
IQ+U6zRQ+Ysia2WPKcLUUy8yj5nQMfvS6yyYTgNVmPLYttzSe8+6jwYD+jmDz6IW
6c5fbGdoVSNlOH29WCgRoi+EynBwXx7bn5pG82yg0XrLEFLUl5CkIJqqEj2rRHL+
X5kbe8vMFHdyPcMtiKpktgR3mzxcYKQ9c5vs3+Qwc3jZJuNSte7KGV1vmd3adPA9
UIZAA9nYh8TmuY3YmKZoraNvVLqJZWVS0PgAIZNwYwfTR8M/W5FHvQOhuAZZqmm8
dcMQW8BsUtkE3Rf8MaNnbkNVr8UX4rQ/DKLstGmdTrAkibaWXXd+563sAyiFPVfR
NvYK7U/ej2t7E8cg+v7wd6rCVxtRImz61zykcLMrOId5w4zeEz69ZSnl1pTCeFjs
RsNKdcJfMQ3+xD1TqcP4dqkGTc0X88SEz7xyUkhJynsJEWt5aRLVJUEz53JUqsz2
I0NbKuCgzBMw0jIcAEGuBbMkui6Y+mI/A7JxDVNxGBqxWXeypUOfx/RnTfibZEAL
7agohcb8qpG1wija66C0H6EB77cKxHAHpS06KR0AdR6vtjqGQlsovae91LG+Q/vN
aAAPhAs1FxjbO4yMxGhZPZsx/Rn83naZi1gN6438Wv8nlsW9cPUWFIgRrECuHNrK
RG6uTyX2FATuXlvXUkPCbTdxciGmsuqs2XfOsJY9gBzmmryc4o67M9fYf/4bGkiV
Am0vIxjjhpwAPZdZmt94mlQ+CUlMslY37oL9X3J5L6xo7SMRVtYdYmxp319ERVCS
y7cEaEJoThO2X+51pg43ZZDAvw+c/PVJyeLZXbVV3yP1oDw4Wevixd48lqGhhTn6
oIAgfK2NDpqWrmhfncYq0n3wsBo0yJObcS2xF+Rri02n+TbFwr+1I57ogHCd/gpT
rv3aGItg0XFXAR/qjHBg6fDZYWi3+nrzy4v5th7GAksHv8VOItLy8S4Ymsv5GVE6
kKAACcPEkUYoGwORgLnoFEysN0Q2LFEdRr2+Pi3bEX1vhY+BWgS+OSGgCiQfA7PC
zUwmvLfJsgMR1USOgMHFIaHzdYYoQSGAJvdONY4Vi49+fzbDvwqvet5IVU+3RNla
ElXywA5jfCWgj5wAYybwJjvbCD42/7VppZP9ySH1KNn1xMoDeAOEenlnzYhG2fjw
MzWMqP8xPFJ0JtFeRb939s8gNS1up/i0Gexo64u4VynBccr8Tu6hRk4O0PpbUCBD
7bICalSk85BFZVjpaMLyPyOheBm3TjLGuJxQZZFNZEeUludKvdbtt34ili7TpVsB
krkqQVP+dAgzR5MqR7icnufF+dnp9f8StdTQktu/ExqskCd+N5EzMzUMUHe5wwgN
1AHHlZEHgzonGYWBY4rSEG18B2FiySwe96VVzLGIeQfdybpelssVC5rp5HAAs3E4
e9sEHZYNr7mg14mRIvjt0/yTM/Xx0BA2ssf8BxhtE+waNio12DHNqUTwfPQxO2z5
n/F1b11XiHFIH5Nnmud0y/IgosJCn3Gu0UetQIUB1BieKue6Hfkj4Qf7G1gVhYMH
fXbNOoUxN1V4vqwbuiRAxxNsKqT+7iof72X8BmZZOvUzKKDwZT9P032WvOydFmBN
OI7UedKUR4DIv2XjRc4yMVsMxqKVG+bZR5nw+PMOp3Fk/ej+wM1O0YT2u7GDbtyH
2q2HxXy2diC9gzAHRbSVSxtAlyKb2ClXOMqI0LH80IjX7bJzHp6l+ibeIvTK88y8
uINIgdkmd2QaXUoO9h5Ads0mTTYRWOUo697NTh9b3bZO8JsGcJkAT68gYRjcWcID
fNKIBdbY3eow6QIQy4ARFwBHQrDOnAF6F/mgFnSXQC5xkI6LWHDXI0RhTgHL6Zsz
2mFG/zdRGYJ3cF+HrLVMm7Q6b2PVVjwM5NemTPrYYlsDMpttVrLQzH1wHS95AqQH
YIm2uoa9rJ5cWxIovsVGW46uIKCECRQzb1otB/2WzfEi9C8bAX/Rssrniltpi0S1
ghw9tHiWdkW/4ClZAKSEDYdb2jh0TbmIzpTlKxThx5rA8ZISyFp3J5W9UvYOAk5K
Py34lLFrq087IpPf3ouRwmOlti2mQfbPS/DG2F9uv/PfHc4dXplOrO4jvolV7f4y
ZVt9ObmRrtPedVoR+3X0gTUowMtcCXTkYGozMeBEK9MPPwNSXg52PRc+BAaDvaQd
EHfElXUMjS+nPF38+HFv+i9y0A2SjbsakM/2Z14Wz+bs3uTcHPAvke2uE1qpUt2p
VekCj4p3feqF78XqSxQIPmgJQj9FL26Rtv8yvtkxpLG/m5amrVhIOMumBzUGuEeK
SZ85Ke9uG5sKHGDDfzdskbvU0mGYrz7ijcSey1uL18MEcFz92vSQR7eKryCEhlZW
WZ1goVO2YuFlHhxMYhRZ/r+DcoMpjpKceo/Jl+nn9v7BHBT3Nnwpbs1K8+xfvdKU
vHN19Fbm0fMgv092ci0/A+cx2JODnWKmIWG27ESxHJVuJnMTGgOUhzuPAKvFzCpW
5RovfkWaYjBcAYtqtD7W2FymL9l/LzpQD628bQqRdQtm1m3lWvGscIMaD1GyL7Au
amf1ZjI0GRH+rXkpAZ4+BDE82aiFKHLnc/flEf7zwTeLWF57pcc2rCk+E5tv2uNH
FrbNietHL14Wxc/INQWeKoH78Jq3COPCNcj9y6Iyz8C8dgzsAegVoR3/F50N01MB
2BKYKcoaNNX7MfvvEtF9siD+oP8TeUvVHWsIPPkL+tMVH1uGfwRBm3tcDQpVGuYL
ELddAd90OJfPIrUf/adevrBDpmPQ4uLEITh3YWiaGs03FNXMWZ4+3E5IUjNOANOY
9ItahR2idMeoFeLrUHlbX2n3Qbe3TZJrqOIsgxuHY3E0VlU0H06ctW6Hy0um8v8R
/+rj6GVoKMS07a6p5Vybt6uIfMb8hQsQjVvWXk/gyrxdFK3fy675cCnw0mBeNMJC
YSeMyk2qHhBra8WR+d1fnTkD7XJwUu3HNVd/bUGEfGlbHRn3TQRRb9XIa0tqDSzY
KxSipQl7G5MiLLFVfH1cpOEmOiRzR7gN8l8UiM84oe/GaP14NakgiGK66HdTGiXL
haElSGFVo0pnq0CVvH8DEGw7C0X92tZ/R6TOChUX0TTfoBvy3S0poGk6gvfl32IT
ZyU6hbRR61kUqMlFPyOjvzOWaENxkboDSAIK6wxmKnrhujB23CkPHY9vkfVJCYpE
DJ/PqK03z+apCydsOe6VwlbGT8b9FRYIvPwLOSsW9TE62V2ZfhZBHw1sJm98Hx6f
H/RuEKoaKk3wNkqLLOiuKD0oRIYWTn6k6Hz4X+Urcla6/ZAqrWOiFnqYZltB5/yF
V9gFf6nY+3npDNXxeHgOE5R/edpStol2ez8fDC7bbfg4mUo6V+3HN5QD0dQYBQBC
pMUJJQ228/0F9cwG40TUhSI3X3J/FyDXwgeT22bHUGOz3AwZvw+g1Jub/Fmxtsk+
jtlY9MDYCmzDVRlflIaASgIMuXuXVWnenTR0go+bFXhedZXzxps1tTKwEbKKwGml
vqeemsVahnV3nbtot95DZTpwXWcvtd15+ZZLT+0CuAYlkJEZXTfN4iWc30Qv5BLF
yp1zkTxmAHhfEPEHZKOkXF8exeXT2FXHmk4lgJPVZ7d6r2KHjTcCUcTJ3ZYZG0T9
foIpge3Bmi1bPFpqKUjLQq7crhpVvu6IVzxAc2AbMlfXdrHqugfbXyWkI3hA+YPu
N4O6ER6ARQLks2fmxOLJOLXciLRXzBzmtwREMDxNJdoiiCPRKGvQ2ycKNKew6w+a
7tvbGP1nW/fTltC4+2OHpu4ORAelHGK+ef9omy7Fia5+OhW3fnUNbd5inJzhH7c1
IJx29dIGmQBySmHpJJosdLMXyRQsFejab/qYivnUVP/YFW+YlJtfmJPnK9dxOqce
Q9qOhCNur/HFbBya7aIBwi/sXooEEvRf67FFyDMW7mbq0vKX+YunhJtgqOmucbiS
DH0l8m8vqejW+LLaDF3cgB/rWoAyPyuQfFBvZIX57RZRCv588jsVYX74+NoGI6Lp
gsQqyf9j9abF915t7p8Hwzuy6jg/8JglQtCnVAE9b7VbYKz2te6c8+ylsx+HI3ca
SBhoYYwLepDteyohsw0mlxLLL+KMF5+9/Ao1uyZ3b93O+R/8Mx+5W7LEdjcN7ZJd
AYEjLtmBkfpE8MskvxICwXq766NVgYtOUDaj6iWJRJVA9KQhqZ84Zmxsg6KRhs2D
sW70JSx9dy89IA/8dTD3flPJjla/3w9sB7i1IQNWFk4Ukd8pLbttGz60uZfCh5BX
mW764JxfHnG+zMxw1hErICVHZAR7otTnYqO08ccODwZjSborUHnB9bjhq/L+5PZs
vOqAHeJ+YxxSB1DFGP38Lbif4NyW9HQQuo/rTnKeGdzw9wimu3MTlB+mrxtfVlPe
jS/NAsK6KF5vDOh7CcLdfle8o9SP2w1hgsYyDux/9OBfIkV5aIxSvvx/FU4d8+Oy
cA6N+Uq+RiLeU/6/cQ7xZI0hZv7gnHAulM22qfBQJenVQWkdi70KIHH3WeJgA1Fv
KIbt/+5VwpXnsxrNcJQWpc8d5plE8WDJq3ccvertXDbLcDQpgMENbYKkoch1m+Te
qhLdYkAoi0/KwA5m6PXPvi5KfX1t+Mh09AFhpVMzasShkErJo4vtNOC8R0rE3/fC
puXAL5afvbBEZhkGJAqC5EYzm6Dcy+i2uyLYehTrx9JMrowmyAYXDt61y30JGZ+6
EzR5PW8yausCKO0A6jWE6Bbt9Zvc7/vBZktvWNWnnK0a7CMZGz/14FofklRsUqGY
rv+XPAlI4uRDzIvNFhsFHANMinOLe8ykQNxqVPAqo3vcxm88neNgF+NFyw+HlbRX
7C0i/OX697MHW1JentTvN2ZVLEPVGv5xdzDTJmQBJFMFJ9I+X1vTBdev5H3GGwmW
sH4di9EAS/EbmZJNEJp5kSc6uSMhGtWZTNwleh5oj4gseRlj1gBqHxbR38jC6pXg
vEeIYZKdV9VT9WUo/id2REBh2F8GiQOREyjg6SwlHw94/t+W6Mx+HCdakpsqELoj
UU42sIjx7zQJ38QG9PDKnVxe3CNUozKOibjvANGYzBirkabGy3hC8G3upnQWN0vH
uXv3DKvPehGKEIg6Mnt2/k4ZrESyHxz/WKSUsrceKpKT29sMLiJoAc9cR9JUk+Wm
bOcfJAsMnk4cSU6DoezOW+5zQBn788CQiNGvJDQ6rw4PXaeyuWcnksmlg7HglI/D
7nQHbuO5Qa6nKof+U7Pxt+RGw584yDotz/sSjjiER2YnvSKmmDSU1FxcsZaeEzbI
RpItfdaKSUDwYtoMnK8Y7fqYAUCNpZ2pxUQ9C0+rpiUO3fAaSN8h0N0dqdxnI88I
S+0FTgF6GOUb2twIP+iOhAOtKO4F/4FWovveWJLKi68erIKCqKJoUaILklnY6Dfe
uMu6cN48PCeq2KWK3qWuSSqe4Urm/EZ/LjJu5douwyxcAQHEATK30TWVFONpd2ie
n1Y6C5BwpnCJTPU8d3sZXMY939SZxFZiMXYycV+k5qJuleYoq4/EKZpjuoJx1CdD
ED1UqxeVg/Z/fqNeZfQpYErZXZhd6BKkYSe759hCqUTzvGwfVEoPDmpzbhvJ4yQV
mjbsSyyXVOqmere5mSMt4aAWrbDgHeOIz8d+bjXOgO8QjdMkejCmoMtwszjwdzV6
06lTkQLgb6SkjBNmhmAAXePUlpxeoICFqDtL8H732pAUvz/G24KlszTOBinqhtO0
4cOX5FIetCsGbAyqGzYSzcGezivkyJunnzCGW2ka4Wkc6b8LgYmh+IcSvHgB+PWG
QHmU9Y36U3jGzzSpJzMViUlneZhSil3tTdHmE2FgeHd66GkUodn91U+M7ubrUAnK
FhKcZ5rW2GeNNRLI45jABNJwLKzqgUYjrbH6+rLxf03NQug7HCW29xIrUXjmo9wd
lKxuvKArEfBD3fOxOGEWSqFL0miiBXF06H7BYYTaPyyLk3gyAREaAxjwIvO+orPg
n9lrVqmW+SoBEjTICkbjpxPfNsJ9ZmMQSUCC5XVIQ6/8LrTSTjA/2a+VqX6E1lNv
6aiD9i8gktBqObAPPWJlhbCqb+R65enkYDsQSAtWbUP/tHBraostYK8cI3HCtdNZ
iRDfLFD+XOf961ngb+mbYDagxFJCeNbpbGy01hKF5zCsVZLUPIgf0tlhFQ2D4yqz
2Td+QHe0sS40jtbkZdR0Qdxp+ezmziKFgxSEgrcNOEVgh7JkP4jhH/kR2E838pjW
RmCwpVpGs8VGRZ7IUivvrFbZF23Jj24aGuE2/g0Y+j/3zX/fnqS9VUiGciAvX6sM
fQGmYzUB6Ulz/Q5Z35HRmJHs70oaJAUSVeZQHQg7OD+U3ILJ2xFu6p7AWOFz6F9y
ppC30IhMeH6rpI32zJ1Td9fbdXeIF6SziadPUXatWpD+HiZi2wO6S0uARHMI7DDR
ovJh4wHg5kNwZm0FYHAnK2X0Ff3RDijp3QgLwf7pbOuERv+H8EXuY+cOfL67hdRZ
wm8vFdqK/4+IlLL8OBED5WdjpyZL8TccL4RuBvZ1qgKmcaaY/gSrpjkHDAUARu4l
nTKZk1s9ehqnQNo6+wFPhdRXxLbOfPW/uyjAV5YFj5/KmGo7JkMpa3KBjGVM0uMg
WzvTSw6da4Jyzfco8/O0fnYUneBPUzjM7G1pMXCBiKOLsB/aq2Q4MHGd0mZNXZ88
KiZyGrBk1I8QCD0hlUjv2nvRlsdwFDbf4fjnAk8PIZ3UnqWyrZ9LGKPJjmOCgLoU
Eh+j/3g1bX1MerwDkUumusVCUsJctlGoeQfYZ16NStndBGymKgwLLuqupEeZA5AO
ZE3dCAQbQf7hrOrFYrFk3Fk9D80oLdYM/TEGVHIBe6hKaQL0zSJJQuYVdTlCURba
ScrrZH/gU80GNPBCUdaqIuGHll2s5xesM+VxrvNR3VUWlbHoccpwZtb3KyWRpzsJ
IqiqeIbBqWGUpL7HPImsN5vdX0AiGxKqn2S/WBHJhM35jMVBaShojs7x1G8efALN
mX6RE+dMSpCy0PrwCQMHb0WuK6r1LDEcpE1KiLoHyQxhFWJ1W9D5m5q5na5106jw
qUnVXYgA+0k8o2/OZJYlB4OzqQSzzy6q9EMeR5Xiwkjaxa3xs0n1R9QRjKMv8Ml9
cMgTdVUk23vI8A4dLFGQ4Ik8yYKrhsscgYzMlrWqiAOkCrPC9+69qAhd+MX5anQL
aTuFJs516QxC+cwqQD8vSCfGKvy4i+JO1jpBNhDRDxuawIsNwA7wDBU45laAyims
6y9g6dGVxVw5UxNeNyx/RbC9uZGkpSifVJjQW7oP5KEhRA6ryzWcHQUkioF+EZs9
kXus1v6rjaj70+sk9SgJVPhAZCOYj50Jp8eVW5yDRa25BJ+WKScoetdxhDh9KABw
daIZgwzfap3sZz/PDndnkweOecio4dACOInhUI2zgcb4z+aVofh1bp0vmzZPUYFk
LwxaverL+5rtM3sKhVuZ1UFgvDv4qZ5bBjA20x1usQ/DSwRtiriZZjrgez4kEpeE
sXPbxI73A8cycn7i5Al1+YRNvIiTBv9M0SwPzNe77pBbWA+wkYx6e3jNunIsEn3m
wQiwRxmVetfEwm5yhwEhcJOCBxWwxJLFXO5it385PsU/coOner0Fg/gJcZFRWjl1
QjQthNbHo07k25bmJ2FX08b5pm3XlQKwmCCV0azhkSi3/zv+BHpEQofCKRv8X+bu
BuiYlZeSyteSdJVj6aFQYd+6vkANzclVYZ+PQ8oY1hj1RuaS5XirYBXyJPRYCPp4
HMUmyI8RZrU4JHXarLgDvot4fV2QFYqDMHtwUJgdqvy8qFlf/KwVqXBmHG9A3tNz
EH2wF+3sh9F5OYNUf1PSq5YY2bq8KTSb5tzuyuWG8VKjXULGrvwldMEqS8mAEGRT
VFrKJOajJDhaye68KpRx9lF19iyYn2zR4j8Q5jmE6H3s3I2iHJ+4mYYpBDmhIFi1
ySwml15AIM/AgbdIuMe2BZjPEAt6GknO39G4RNB+0LvouFuNkhFKTeHBsu7hMsTY
nSMzjHt6mPGZXAQiPf3X51L8BSqtOWTKCR056SwD0ze1LDRzu6HeldiU5rMoDmrw
VNIFFHeB5e+niQBZN0EuvM0DI8dA7OKKgEFgRDLhFmWkgF4c1EX3sHwpfHXCIUMF
/VexGjK3bozslCjxRngw4JKpS8BYRuhKDd8M+t5uEBw9sSWtalmZFo82yWaQHVYE
I9/lxYzbu8h6J7jpRsBOzZsoNv0xVu5h/4AlvyuYru/UGNrKQ4uyNrPnMr971EVH
oYh7s6VI7fRyW3BAil26MV0OVwI8XmwCIBJ17bou/HmnPq3aIOz+ziZdRgUIwJcj
A0YhuhSWk7kfBAoSNXNkDje5Dc6Rp7us2XG5poAAKbCw2gIdiHrE8zOtcLSCy3U+
Xc8jRXnZvWIR8BUg+p1WJqKxsOZpglv0lD4Qy7kNMQ23KBdXWk+BLmx8j79a8KsB
OwhXrxh8hlCvcGIgwpTYMblQk7bsM4CQc0D62ly4Q7k1I3Eu5dv1aiSn7vIKmYE2
avwz6FQITdKIlI5Kl7rOdO2mZz0ySmq32V5Gq0enUwKecgcq3mcgwiocdNj80Mnq
102DQ4muscVwSJZ8PsO+3RMeHUnAvYbHCEYpdGUmYY0FUZcBGf/Q1f9Qwrs1i5ei
GGvMUKcTlV5dJfOaCbZzNey1DMpwz8jT1AprSpi5PA54JVHpuaH4ddQ61pK5GVly
RRZBf9p68nBM9YOz/JasrF+hIy3oo9k52DQEjKvc1Wv67byF7ZcqcNFtniJwEDMz
IGVlBRCRwjgChe8+8iGTPyFG7iLUZF1I+P3LXOmcNcOtZlHkaq4zXda36H9L9wz1
XPpDEB4iKX6zM+bfD0SIuOeAnC9t2cCO+Y8ras0eHFea9DVez/b32KX3MUUBGF3H
o+EKWac1+C6aFOVi6OwZtbF3r2R5lt0Lx9Cu2+XZ4qfkTSwk3PTA2e3Xly8Y0rS/
gkHomwBmkiN6/bs4pNR9+rTyMMaG2eS1rpWaf+1ERLTtbp+8h5Q7G4xdSBWmSpqG
EVuq9zfIAXkiM/z7hr1BSoZXIWAL9hwiwwkqMg2FnLLZLmdc9S98WfFOFS9hzoql
dPfnhrTkpzqEXrh1tKzn3Zbl3+H1jiZZnjpPQbe7lYu+1GiKho11SNhCP3aojyw4
taA3F32QNQHKKWdqFOlXRq250H3Ss/Q6LlSlrIlF2BhFdsgw2M8Zin/4w/qlLtzP
PpMDcpuzlF78zGjow176c0bAan9VZ7hXvZsa+qIb5GkbpWJa5lzTAIPLCUupSCyZ
rpufrr7Z1y/kC3UzncZxMoqeM2ZL9YFEpSsaUtQIRo0NUBf87lCIE7YHa2SNblUk
BTQo7pxxnQJ0h9LlVe2d0dEv+WC7WaEcrVdkhV0Xopwmc3X+9uWtq7PIE6D7S2yl
0Uza7FCLLblDfT5x/KZnbMnjO6kaODtdC0MSCmE0H0taXn/jH8K5N/e9ryhvwdFu
1AVoJ/LgwFZJ+SQVxUWnAp5ajoyO8KRDjalqTbfL1s2QXoMdafLQ0ZydrXtBcpN8
5xSm8Sj6jNEzCl9TbKt4Axmaw6U0/qgsQMq/ozPkgifS2oge11yFc7krP6fwbqNU
S2AQuUPdQCvAtSQLCD8ZC4y0809okQ9jJAZJ2F/8VG5EMrieGz/Z1Qr+JxxSFP1Q
wS6cGOhMhW7M6DWBGpBf2guG7wXwbi05n3EqHkYPVVIcjOpwT5azvUyL/NzNIowZ
E1hKdnl24INCRfCMA88twEn537qWlHhGgT6SoDdlLS1yFS1IPlzH1oxCCiWMfQfy
KA1ILwU6ArhCje92aMFnZFGHy3V09X69bfLFB/iAPqyr9zFhkcmxw6fMY34lPRQU
pQaw8DvujLCTq46runQCXqfQOohLagZO10f8BVVLVQakQyXNJXaq/rbptbpz6J9k
KxP5vMfXBsul4C0xGhyOUbQ5g6Zzr+DrvwtmeYJO3IYQ2Y9E+BivlE7QnExQMJjD
jEcYzOBtDTXYcA9/CGOg9HJPM7Lz13PNHFPhDVE/xBO9ozmo5ZORemlJNNIRiDMZ
8h5m0KzcA0IwFLpWdIlMQEqfCGpxZsQku0/ZFSsBo6U4ZGK69rFgLEWKnqYVo0gS
aGnn/QOXf4M6+4sM8DWWRjGXx+BSxsBN1MppeNKz48okoeNV3Y85x/ErLi8iK2XV
1sSlxNnibm23gkzEBrk5CUhTPB82Zh3VLkmronVx7jYj7QHXzQUQ5TRrqf8Nk3fP
0M4xDWUTsnggQwinGnSR3at9hsUEkWO5ppYYBaoLRf01O0bzEbvt/2g2KmJxPlDZ
k9QUlNckiM09gyHEvFxylPoh1Eip7S4zp34STPGhTg68uwP35PUjrSMLhwoRgmgr
2C6V/rZE5AIys2jl4usuvBVZ6GKQqExeaKzUfyopF91LOLFvmxRRAlYGAH+tLvvX
mewkj/7xB2BbqprjmFo5sIhk4NqUlF3e0yA+XQDN40QQEjpedkPl3BqBM63ud3ou
C9FGNTkp9lHvuiJn2Y7P2562ugtBX6RjkxeOmIYARhm91egoD0O9myj+bwkzpV7J
HHKuybkEihtn5QYJ1i8e1I4ev4zXx3+rKYIXwgsucEQiXBrOlPMoeKxGC+8KGPF1
hSTGSsc27BoFFcQFiMdx4xQ4G5cAToR9BIPVuXaqLjcox8vdUHGvOwHJXdKW7XG6
50eGyg3Ltd67DrX8Zcit13FDM51ppG6i0IBS31Lr8P2YELMir6Jomh+luYVecjXp
wCzN7Ac9bTbfwqtaXyejLXoFygGuKvK5H5JtIBPy9/no8EMMEPG3mtxfhg3Zm4Lu
EmlohRE3uinMp9y3cgnsb4l/1cyS/D5/2661oL139RUIdJfNiHtFOz1mS29yN6Je
qS9ezFMf/NmbPGNm2rSK+/jeirE8WRbZVHY3bBnHbTxcGjNSs81+wzJVjFTsv6Ny
fAJXrnBPim+SG6icWD9oMTcxyM75vQQk/wygb+D6LjR8rAoEljI3PDF/S1EgmIel
qr0nNMS9bkafSWz4N2k8/laA+B5gNZU3puBTJIkq/0DgyN5DRDTEzdckbpsWy5YP
UllGbCF7X7oamYt9DJ2aVm40hLz2tr3+r/jhmunlSTF9JDmWSzY4/vFNJr+lubzw
G3Hdih+49+LNU8M5GhhUnIpoa5CABCJbO08JFuJXB7KC6bDQ5vqlFDwNbEXyaPAA
acvarQeVWYOzVpXe3oqePTw1aMXDx2nUkCl5LdoxD79DyzFOdSxd60a0Ew95JpwV
rD7fOTCiRkcrjRvx2+WlXA0+kX0pTB1ZUUbx0TobeqrFiXGgn40uRETuotlzKg+V
YgadfRXgWPZoeg6T2MPeXEC9i0YZs8RBqAp8QdzJKot29/c+eaFNn3jgHpRasKUA
vRLGJCCIr7huZJ2AW5N1V4aXkSQBStNME6EdsYUe1kQ3o61qLT83I5F1/dvTdEAJ
y4nW3xaTdlS7eGOPQEVV7ZjLv6RY9FPmU7d7yw4J3QmAFmdn98kVvjzQ3Dd6LgoE
t7PpjdgtzwKXZfHQ+XKyU+zOvjVC75EHXWpVlBryUh1nZ4JsdGb56nbKfNFEVFHG
MkK+J/6Y5rf++UB1sxT9kl3JAB5LFkNzLAFJwmrj5pq+NFikgxPKhegGWgfm2IzD
GlHoUVn93tU2SeHS8Ul5rLbqkj/vl79M2ZY8XS+MlzI8FDcgGfSkjOKLjjc5dih6
MInd9Ky26UIvgAV5HIloaHFFBFY058mi5VUyuUQbU2sUC9eAaANTsj7WmFdZuL6O
AGUKm1zDyGt6vADve7ZxVh+rS1TGJXnL4oSx1TAA6J7YSkYvC/qp+iDp8Qdw92xO
xXIrdmFdnF2UA6rw2/3UimtTEUCq/KQKtPuPI1FcrLVVh3cZG/Q0+Ao+6yJpVPjl
Fv0MqGFSgLLdnsi7RRzloBd+FMkJHcEQ28yzqPpIKOZdbmNPJxKD1AFt80SbyVv3
RoAqrvuFvVVhPNfsUtNH2yQmUayY754oH0CjZUrSPEavOub2qkkCAZDQ0lJfbENC
U0536f0lG63tETJAa4xTfORx/6mdlZBRoIc9tzD+QAS6IKaszjlsx8/cUXknbwq6
fMZCkczJ2ofwjBFxCSwVECAppxEnUZs3h1a9bAMmN1NnwTjlPRTsPWpT7kKurgot
xru0p0peo6sQMLTOFxaOU/UFlbAgovmGOBmEtek41sllqpqtL+0cYDhMYzZZWtqf
iaRET7MQmA2F8CA655pr0RObr0ApFZInICMGgizem4iHj7gS6xA7ud5WR3VJgfPU
78bD5XGNWKxtDGQsCiY8HKVtWBTh04lub9K7gjz1j2ZGGbAfd/rE0yJESy5Xdck3
IWAFqlyGKjzWtqKRcGIMiHHAlUsHtqcA2+qK0L2W36GsM6xgznEAoK9myUYMyMwS
S+GqhvcSO5fOLru3qd+8hOf1wHwij/MKokqWXrYnthD0OZiqmFS//wwVJWjXEiMr
mI8eapVWvC5AKyN3ob+9K1UPeqB41sdmu61VwFOA0LkTXNT1i5q1g91yy1xikdBA
HSy8+jMP11wMvB46U/1jstyMXNMiPgwVbxq0CL041wHO2dR6JewxJya4SlyF1sDY
cJlAX/i5nmWXxU7yZQO19rKbn+dNLuiccJGgGklBjrX+ZlPV7In8MnugZyXKPwy+
LgHHRe7GTZRhmln7lR2zEQ844dGvxvtikkYzZvS7lVbCCHy3yr3dBE8o240BeutG
MC3jJSavbHuG1VSp2NCWMIKOn0CSoEGBcUO90FJgH3s32UVyKVePXbjcLqx6TWFr
INaEHJkCWpwG738UtiDolOJDS4sIXeD4zNS7M6O5kOlUzkemg1r+y6IH81Z+nRil
FXt4bsiKMAZNcdR3s8qxYpw9CjIi5wRJ5Yc9lOnpkzGuTIZ8KMVayawFrRyzCec9
hPTieaSCzbgiepbYB7JiWXiTwtupbRp0+/EXBhBkMlT8eLmP6VSbyPF1GNGH97a4
Gc1Xr/SF/2tN2Hnz4HOa9DnIeWe7GNZv1DHcp7LSE9YAoiEKPtkq9o+8AJefUv5V
z9+r9dU1PubIMfvew827r9S+tj2C+iiN41zYbRvwlyjHSYrFZaSpvYqPEy+ry9ld
2d+fuR9MxbslZMVwawcZL6eQNnCTJrFFTOAKWX7j7Egzt3JA02BaqDazcEXqSv+m
t781qP7/s7JDbz1OIKcWYNoF1/zmekYvCbL1L2v6FK9kKTQh7MDLqkyc3R1u21DY
/wnqCo+Bf4yUSYwcVb+sCHU0wXM+gBmPhRq0ASTwMiL/05jSvcl5ZlDPIKxs4KaI
mT6NCv3NqfyjOj6nGlVJTwL9fIPSC24ZgsRhDm1bCJX/3IIsVNBJUvZyskwEOYCf
N6uzaauaYHaiPv4n6Vrz6fcWYuMUoaQTw2JT4vW7uyfWtt+PlyNOG4hltrxGwGFK
g7o4yiq3/wyP5RXMWJWt4yUMBH6Ar8YZzbDqqMvDAZIR1BKbfJtHPbv24vOQ49hQ
PV16vu7lo3qw271sF+HeXkLFXIE64eG7w0IbEXxO4Th1fFLzwYPc6Q9NoxyN54TI
1pxAUQ2F6xrcAZlRZdbM+h8tkZmcE07L6X2quWyIla7Zp7nLfw+oCx8aaZkpKASf
m/5Uv7cagMhyojing0M7ZYLE/KuIqEq57yK2JyfFVBH9k4ln9RcTLx6qPYForWL/
Ymt7PbTbltWurqG26epsLsSntpdPjmV0tKUwoRNdrAmVW/7ez/eWa5r/Mlkq7nbq
O8wP8MP6wODXa23rTfmAc+heXUYyHmQx3WfHN7jIS2eCAm0UnpDWqUQYBJ3vopQJ
eEWwB1XflZXTZG2sE0vENP4W6eNaIcSi1n94W4s/+07k/G3SI67Xbmx0pSRZfi2q
EoPVlbPuqtuaS8t1f6dy23zTByTJRNNiwAMpubE0Ec1JmRa4lhQ87u1OCGLOO/vu
QDzzxh/kvRYdZRpSDNCQGMONo9oHmNNmMwMixmuoSB/0AmOng2yBy3nxc3JzitIK
tDEwR1GO3C3xpKiIxuGrG/bx59j4uwCgNrti+ED6Mw4YFQhcyuP/gvqjdrVbX4eY
Ndksp7k7+QtT9eGDysdLzRRnxqH3r8PJJ+8WCf+3C7fUkH4TWzWsZ/+aAe7QpFTu
P0ayE/HhOs9KON12oSxRTahrsZ5lRXlALX8R4Uhzwqu3w7JmtUl2JfZXopJT2rKc
0jw74Wm1yNbhPCghWOINXtxULisowh4PMN17RXpTKLG9OjOe/Im26lDLagHQ7/Fk
PjhQadMHVXQPJBkaz/9PtQoZzmMrazFAphEb0ezjxSY1hVHghhX482iq7xD3wJKX
FSEY1azjfg4WsHglF11LWhgA5/u0XYq3R4lyb2XdmlBejcS9uBSNWBQOXzALIOgG
N914g2jS5nIORmFji3pY1Qy28vgQHfE3F/oUvQiGF0WUymvdbVzD2Ov62g7/ZcXr
fUH6a21M0rqRbiuLpyLDSfO02bShsgL7a4whEL3HIn2wYrnyXkBbBubl/nAR0O4Y
rDzhJRf67n9d1RUJJ3zF4ruOaSGeDJyly+kfsLnQjqCmbqdRpe69EeIg2Vv6CBmT
P2S21B5xybwiWAiowZN2kDcPw5VnqXP50p/OsqwRfX+NCo4uK9hWtg25ngjLfrzS
skto5TYOPbtKPBTnEHHHtfHJbA0+umOwhRSRA6fRHTKZ/Q1OmdwNYAV7qI0WiCHY
kWHrJTmF5Y1X3QT4hKCAQ/+QxSghGuBGlRp0amvR3AKXG+Sb4Cg5KwVU13aYHFj2
ypeD8OFlNnTJ0SVAP14gocXkIN13KFYEfIqJdICBaynPVGVyoO34oApoPmpd0KWd
nxaldc96o48X9UcLRzidEclMw4PfxPx1vwJa6LR/GelpVLfxjgpcF7/EpFahyUJx
zJCCCFiq9xnMhrK8I5myLBuY1fNzXMZJaK+JkQHkeEHcnKM4ENQ0+h1i/Aaml4qA
wJVY1mxgUVFVBPhv2miyo9BA3Cf/CYQntDPawRhqSEw7Dojwl9LLskGbGIVCwwrB
QenR5rQIbABwiQjuYce6hmRMcth2PqrZ1Fsf9iMCPrv1/r48LXWLJj+FpKEgMRkC
bAL/duYTJUZDeST8A/WGao6AO+/hPvXJdk/Zz01r2X9/aTmRWw/h+A8rL/+Yu4aQ
7DapGuDQsK6DO1Auk3UI0mNE7AIgT6khbw3ShR3bUb+OWwwdW5b8ayEvAybRyhEB
P2iMpwwaARX8UrtNBM+CDMHSFIzylDSPRJ9eNyNQZwa/y9GSBe1uq/CiH2uVvMzk
Z6eEPPzrytSVGcs7O8EYySnJL2pTHP63kXyoXWZxt1evi7oMM3SM/5Un4W6cnjfy
68n4W1wyqTeI6/DcGugPfal6Xw7vtP5zJjiOtjf4Lx1EPID93MW1twCP0GnQGrcA
BbwOiCUIEtMqjraVUVkkZnddwKUKqekv1jo2kAq9Nc6i2Zy9JtG/yqf1/NzFVpme
XbwaEwMsY1NhWgvF7tTMrDB9H300JVtJS0QBpnooJMGA3fSXTwEJIFtxlpM/VCrF
P0P0Ua7Qh+fok87R2jr1drPsxLmaBWj06bi9AcwcQRrsvxKuQ87uQ2XXZNENnqU3
we+YA4hi20QiFPi0W3HQOU75lLz/ArTLg3CKfEEcnl/xtIHKOvHqiGFJinxyfxJi
u85cuNLHFgved70a6bEDDfQ5kyrOjonsJUB8wxAW1kT+3Yt81bR03qbqdlRfxZSB
SnDItUoADdZThWZNRBk58sj9z0+1UzTRwahUOZBirkjBRoCPxmn+RwSpzsnV3Sbe
CzoSVdbw7kB9Oeoa6VHaEbSBeK1GuryXTpFzPtlnjBRVMLeh8KPMUSDDqCtGUZ+z
AMB3OasTCz2WJwz2MYIF+1w8K/lDcbFGm/64MgZWSybUXkLrXowL1BCnKdvmFicq
OCNSm4UGAIoQziHy90mxvVCaN10CZJ6YZxDLUN+MLJ3WgxoXVQ+D0z5ej69Hr3GH
P2w6u5qAernSA2sltb1GEd0NgpE00W7YKda1hbIZL3Xgk1za7pWvDRdkXDHoA8Y7
e5uKjAAj42dZ/3WvfLRd/fTCaqdlSmHNZUbFU7s2eqb7KhWOXIy1FywpOZAUN5j7
wD7aO2kWTCy4/L9va3EWBvjfen83J7JkEi/1lAi1kgBLfissQVKYf+d8cQNqEpiT
GdIn8JEeVvwobtzpGyfv7q+vCh8oqR6fU2+H2gbhECuDEhumzuo5hfYFH5F4CF4P
7zuxPFLEKsvSMAMdvOfFyyHUPOfgePo3rvjHXd7Fq+y/nEaLB0LV5XrB9kbv4KOZ
RMCfF3xW8RfVDVm7XY/IFG6lKueFG5rOktWu80ZvuxGhYqZ+TQnMMbh990zG/aC8
X57MV/N+mfza5cq8R9r16IVGEKVKYDVmAbot0v5T0qCdwEYzCQrXbFI/wyPuU0t4
M09TZRbfHIEfLNcLhsE7V82SB1QEnORSdZR4CaoeQORC7/KA1+hyiuMx/SYcHvQu
DSl5NoSHJir2dojjpU+kXOTe/FUpvuTJ+iw3N/otNMralINfccyNJ+/84d5/bA3C
AmjHK3Aydy6AYTVXZbkcQLAf2RRjrefXTydcDy27ebq6vWA2wHql/7G7C6S/ZHuJ
18gsi5treIyedLsxbz4uG6Vb19bXb93+I7GdnLRtjpWohOXuH7xfnHuSuRZJ2qFI
XdRGy6dHPPS1f+SWAY7zHR/mN1WD0ksZ7Jgqn0gmhRXuPOpnJyC9iacDBPEIJP5M
F6hp+cvyoH23PEXaPLrEueMlT7XddOmtRREVSop3sSJ6P7UnFrwEr74zGMsMFqol
U5lcWlV6Iy+cwSRLNFyai1UlbCd0fWbEeUI2RcQDNRB3UTaA6pBCAIIep3t2S9fl
0a7RE92NorjePdUj4m1UhGq/tB6xRUjQsD50Zx2tWRifxPatiRjfwqLounM5dzf0
v8BFIiGQIYxqunzJXEB0DLwf+NmSbRR966z/yBTKiYhnRccIQy6DA0/R6A7najJJ
Uh8aQATLmXl0dauLkA49OLKjXOAdIflI4XkJckhAoaqr9g5/PEcIQ13FrYlkR5Wv
FAOZaGjbqBoZuGet/FaiucDDC56LpNQdeLArWnVDv+nn39NHMOZgnUtkviNxc3G2
0/EmhRSAJW7M6uKFNp+KQdtZ5/RSUz1bqpCKAlEUWU9bcwpwk87HUtJkHZZdDwoE
P9yYD6+qByC9Co/hEm6c5OIGgaYGkaaKif0egDW2Mx24VZNDjOPLvQlwkKaS7Iw5
iktQikFVtbzXG0nMEVA2J9iIErJ0Sk1Nh+2YJ7k9e/4rTqQ2yv55Pv0tMA1NJXTb
he7OAt2z23CcHcZLxLHulW6QvFuDuQryhrvGx+hCtQem1FRM03zwaWmp1YqEPGx4
LJddKbP32g38XogwefsAAa93GJXarJ2y2BNallgP04/ma0iSFmQOaT+QGKAWcWI1
q8rgfAHlXEUXorV8kgo+CZkML8vpRKPwww8vPkzs+X+lsVt9TpCLGw1cE7PM1DDM
1Sw+26elJ3iJZsLTc+W3LIn7gf3jDppXD8W0Fi8XnLyWebif98FI1I/lnQJK6WEp
E72J2dw4Fse84re/PFG7XsRXcZAM4O6umOHo9nH3ZAosw3asnrf7TVCWfNPjEW2i
SCYpc9iQbinGTtsHSUQ22UhWRE/H+yDPIRIrjM+f5b1O3/m3vxuzJfp3LVDUAvmS
2iTxU6nAUX11Y2BowCjwQGoU4MFUw3RP7bPmrUvz5Y/dJBKqWh+KcXNLy7k4Vrjk
CA8QMZe/bOCopMTfZ46adGWQdkqlXQ9JDEqWMUTmaNJGzrbL8g1uG029XdlieZnh
IS9QOnpghtPBCp+nkT3Yw126Tu6lyXPLYReO/quWWPNLzABnmKJOAP/XOenPvz52
YZjpcIMXsR8+H/Ha88mlXrM22tVPbsZaNFcpUF2uVa6Abr1z/ct9bFkwnagWEpn0
DwbptoQWCd3bKokoV8OgytAcRpCM7xVTcXZHFjih4ouB8JlXuBlcDsmZi44QxqCZ
NklZ+yXv3iQL6/hljgYJzia5q+PDCvKvHR0YfOtSC7QW4rFUuwNjfgrjxb6txqig
h9t3OhdWxLpg5c5D8zt/8R0fJJ5XVxRy73I3+45SQL48zTe/Z+ofZqX6yUYm7Rnl
vVvzwpC+nZo4jddyKhapeoUWFEGxbmXbWNi0czxx0hVtylC1B4/tIdOvEnuhUYcd
YR04tJl0DrBRkZBn2EBlgYHdhAaz5UDd9D6nUiPRc6pXLjrgMojhy4kGmtXw3Pp0
EUZ4oafXmQaVPF1OSeyyTKkfcfVFQfa8+Dxwi5YbyGGXxOpoH02c+be/ULVGz0pu
BQ2V9zJkV7NgRarqFdVYYUcTDtR2ux9NIoGBP/y//h6aqr0vcdXO7ShXwI3NbMkM
lxtQdq9LsjRuNuKil3TRZ/ObDLwXhxQBFW1CX9EeyIM6bocGq3/pgzMVMYJQH4J3
+tyeQH1FGY+TeVb0+OknX3BoYYEqIrj2G6i0NE+/+GQCEkcCWmaamU+Fg2oddnOm
IxGWtU0ASmwPCHRu+eH8MRHSbZOKyN4UxxOa2zLc62UIwPnoQSx9JzBeZbV83hnA
gcnztwZ03PzQJpMLgObkzUSrW/y9m5EpzJlga3Kt40Ix3h7Fmk8tVZ3n6xGc2gTr
SLV5fTROooAYwTbqpUZuQpF3U8u+BXTj6vO2vxtB/VPT8Ia73NGQzxy5WAxIamtC
yFsWTrtzuGx3zcR2HsaqjO3QPkkhE35om6UIu+Yjx2zKbWQpSgqVs5g/KZDlU0Lq
mxCYqV6XnuBqb25AwygLNly2llISEPES69twLfzblxhYOB8wtuGAsfS2WRGYF86V
rxCU9r7kxRvJIcjS+/0679UaBF5Ur8pXG3s2+ckczX0wQF+TU5v3eVyrtU8bTxbK
546JUt6rTfGj1bVx/sEViQUnoLQ8c/6jvhNrgeHMdAAiL/ac2+yCDQ+m4Axnf1ds
zEVpQR/4bTRnZfvqJRTOwmViuM4XoUlMoI4BGYBQfAN0/yVFMqbQomcwaJuO8MYz
oJKaSkrYKrIRd3wAPj7USIRvhTfFGu/lS471m7UnPUplq0eSm4chswaCIiXN2OT6
IrEcijoeQVSslju+BETn07bvHWutH1qKSxclIHIi9GOydDv2SuehTIguOSLIJ6vR
QlKZFXGRS6lWPxbEF4V+W7b3875Iux3UYM1K6nqTFnXpBPn07+CERIh3PoulXerL
RmMzb+ADQ63eEGn+hsdu2MdqRcPitPcfzW6q0STaOpCRMtGGc4sRbG5cQB2h+2Wm
E0t3h7NYgZ8FpbT66deZYJZINGB7ZaBmQGNGH6Wwxp2LMjIN6TZlIFB9V0/sb//P
kwx5zgLqjSR4GRWBwnYVZW1ODIIqbmoKopu94CT3+FTSCwcSIosLslp8+xYGnQix
5HDjrKkCQ0UQK7+oclnBJWs2vzgl5lKxeX48NPzV9hq8zkLtQd0B7Cz8yxQhZCA2
0EuvsRNAdowqVSr9lwsJS8P4LNHXr97G5awCt7mTz9tmG37eKHEWZtLQLBQbbGJI
VCa0zkWTTtR/PNlHfMlE99e/GVC/sTwLxdGB8NRemfzk9aGcdALBk5nzpEhCJHDf
SVPWnKYXURnWmO0lgxXPByDdO5GMbuRIlIeOCHrtTQxTcl8OtXiKYD0qSqwuPTTb
7kjXA1n7rYFVCMciSGGDe+EnjzkQy1JJaULUKlxWtsc5rp5sO3B7HwRDRvz9pGi0
8AdFNELCOTz6m2xeBDyy5WPSSepBBDdriln1fDIdFsGd8KA3jfXTPrh7Bqdqr7nq
FJO8+VhT+ejTmV7WNhHMzv5xxMR4zFBOov9wkWYB3k58emAxFjEqOBh0PlKdIVoF
xDlKd6vaadHoSrBZavYO8sJwvQexHWgSE651phyW+LdfA+A5WBByMU/yxgfwL6Nr
AV9wLm7vYtlbirR4IJNtVhhdtDrb6ellIX2Odcz5icxVTqAUOZ8/soOG9JOSzNXb
5BE5XDUSIWm00qu3rwgkTbg4lv7fngH+aNtsIaeFhZI+nPaofG4VUO04kHxGdDDc
wMcmS4SslZe2F+OR1zxUDuoWmih91AbjR4L1NxOgaQNVCm6OaN+WvsuQda7ORo/2
8r6AcAJ/NulXfz0F1oxuOPfIHT7X1kImMuh5gny9lUj0BJmQ4WUy0j0q7glSaDsp
V8MvS9fmuDHgW1HHcePbncbQxz/pzK1YRdLIBy9UDR/dnuaK87nF/zZ9cUGKb/LR
ied8rcxWWicqgWz7OdDXcm6lWGqnmsamGi3n4v+njTUs8eYgeGCVeMSiimztzLeV
Q/AVMx3TjCKni/SII38Yizk9G7UExCV7LpqJYEweS65MjaxsAp/pbplcXQIEnvJC
PjnZboNOa5UAI5gESz/EB+L68itgU3PN9Cboj4cRwpX0oWu6Ktexp0ioi9s5Lb8p
0dED1pPEfy2NHYNJJ7q+C50+KsqnMJpO1eeU6BiNiYz+dcVrKddVNLJ8e31cfvY9
A6UEsNX7Ps92veHYITxIVQFlf9sa58mksbrbAGPojOLkWuqjwKkUEzbJWB1Mvb+U
CkxHvSnQrqdtDENj9q03HRJNVGH9oNpgClCJDj886knwGt9FeG33qh8Dby5VDyQI
hfO+p/4KZbVfEPh8fJ40p/f3khPjXq+MSdlY40tFyQKahZAOJHyjJDfmdJJAiN25
LlbAW/LsYCLLscDLnn+q90b9SQd8lCe3SUQvf3p7VJ4MSQWUH0oClx8ZVJQ+n60J
omnJ/Z1BfWdpK6kQue8aF+11ptzBvHcyKKUuEBQsGFnXgCtjxj7f2AallC87k/kZ
KjYS4gWoQViobPvZpSLFRDOE0tb5D99unEe01SgXgG3/jwNv1b8S9pgPGKEHGktO
ZP3fvLaMH3HLwjU3R67PO4HE+24xuIzfjowSZFEx8bqRu5HYePR0LJOatjFOvNF3
T8s8jKW1Fp6lzb4pRMTLNg/XmWGMGWR6gn+DOU40LP3WmkC4bHxo2akbEy2ZYmCN
L0IirGzlTptfopk1eWBQNSr28wLSxQZluo2jHRiKcQd0fboWEk8aUccgKgSAz4xT
jMCa406xMhiHmxGkUaR/QyneKolbYMisxIab4fwHmr/vDhDIKOuk2lVyOnKyrdf/
FVJR1UvHmY5OkS7HHu7X0kfr6EFr0RIO2U5c5LkhGC+Op/8ZFhcJx9pLEmNqlAj+
kjQRJtDnPFJtESmFjGycleGNfNpAZ5wsYaRIUn0ik4eEGyx7MLPeOeXNnM0bT+aK
E6DGG+/henJf4EOOjR0B68DF05rzHB5BhSMU/LWjv5/gdXlq5c3Ly7Vl8YyC2ieP
VirNLB5bks6lqyQsr+LGWPDkV8CF3vT7ZQKgzjrMyNPqXKzQvo11tfwbft47hk3O
elsC/vsaAz8AekMCL1SgRb8qsW5gj7dLh1gXbw3bQbRDlK+uL5ihTnuiVM89vGnd
U/33VYZsGuCExOsVVP6eCWYLrhHpZ2xMqnubINCaU3LgxYRBEcm5ycRsjlehC4+S
U0MZnE0VXbtJQ0QfAzCjuDOEm+IXQZWrIZVBoUduCJO0CoXsi7CFloCQlZ0iKnQ2
eKeG8K2g7nQIJvq7PQ97ao6LWMUj/SWNg2fHnDSBdWTVHYpHx53oc6cUF4gGswab
HsQ4aWxhUSCRi/yOI7I4LuFLUIIiBRRgWC7M5og9GaURgXfHt4MsQmLz9sIXMzAQ
Vk/C04zXUD7XJ4FsPxBfF+M9Jmqyufrzirc2Hrhwxq9UIl6QM8GMRtP9KA21ZOu2
VH335oVT6IItf4nwGaVbDjmcYFpOXinft/RFMl3AyOE64Bt5B0mZQT55V9ZqhQZF
vmIYExqreSiFQ6NXQJuDYsTenAd6X3QpFBmh6LGiSUy9RM+pvcSe9HAgQq0671R6
iYY7m7G8iF6yToqwAF9UqJMSC6GCFWRz6tb/3X0HZmTg5eTgk0JDM2MYAnkVpfZZ
F0MiPx+T8RCMkNMQCmZ8i3J7FvuATGfu7RKrQL4eNEnvChccc+X11SuU3Kj5jYFS
S1o6yqcllOegaIkECSYDhhaCkT7aKgAJqNPvOFYsxvTeV3B51tKvz4QSiYTVRvS1
2JHaHqF1y6nC1odj4EsM2P0duB8sOH7qnHGdvCQmluhfFimOFIagWcoRrLy/CGxL
DaiYF+7dXOP6zodeltwR27IhX3BaX+zoqWLD+G1jS4Guw1KdXB3cjYXvXnkzI8ps
+jQK0+Gc91koftuYout4IC+hb4YLw4i35W0DylFSsQeofhaUjrQNsw1PEeldSh/p
aY9X5sCkHG6wyWADH3buhZrhy+N/hbWxXBYes/jkN/q8rqWlX6poENHvxjVSEsNA
pQZBpgumaNXJniOKydGm/ch87NecEk4v/Sp2Hs9QYf7exC2N3VQ8a4AxXqJb5exb
g+f1biQC2fdiLWsbGCVI1giMCxC8b6//tO2pWqFDvObSlY+Ku9THsiaVIfm+GXFu
FWg0uyapv1rgGqYp925FPMFVTzXh1NV1RjIEZF/kgI2zV1o6sGmKs5+HmRw56+Lw
AjgEIuDSZdug0jeRTg71QXVxpHEtnwqv1qqoHAW8okRGnllQfJjc9ezvm8u0bes+
W0oNhgfiaLqiqiZ+K2GB4UIFzNQzPspGZBDEMaeMGQmuFGDwcdva7C99xQSxNm8d
BMIMa2x0E1xq5NYluHAG3v8fKgsWiChtH5BoxR13yo0pt+P9ZLl74AgMmXtpKIvz
UgvYogeOre/8DuR9nK7SvOlamChmcVrqtKSj4esgm9C8iQqR31sOeE9PRRjTIF6x
B/PqiapjPUPI173mt5gn5LAv/N5ixpfVfv7O7d1oKR197oamADIvtYlZ6mxG0qTg
CHXE6t2U2in+VJ42FHDksMMMvI90Zq3uJROlQIAmCqA+32NQA/xn9jqcenwaJVuN
Y0MMW3E3frhfkZWhJylp+TcYk2NIhVI33IHvZ5ZcQHhH3zdvIxBcbgE50tEVs5Ab
KL1i070I1WwdTm9Zcb3vqptHBgeToDgqZAZIWMhLU8DTa97MRFEIrMPxBmonJMU9
JyzI9wlfo/x3nKRMZhptofbum8H6UL7bgPraE3+IPmaonJv46IacdCs3jfVZXhA0
0FyrRJoTnl4qMkV/vGyan4vEkNhxU439Z06tp+fuf7QhwKROkMEvYq676J5/plZ5
RXAkB+iL7xoMiz915a+P6+HYM/B59VW3TYhEQ2oX1H7kYMLQbSiUofHov4/OtsWr
Eia4Wo7Esw9Wgzxs1MoFg/9b0na1fORey9ik7Pwu3aHOIUunbgfSM8q9MNPHFQrB
y7NRPxLMtN68hCYh+eyR8bBezL9h7MIUiUE0O8bRpkfp/WowP7jL8adaDRvXD2/y
ApRxq9ZFpM72lztDBnsbEHArPNRJm6OZ6t9ciKX0FC+6194WAhyOzjAUIv16grWD
YfVGkRcsjMv4t25U82UlYCMxgN03AH//5pZ2FXMA2oD4jr87Oq7BM9NMyI5/MqVJ
zbid4dlfjnl6+QbqAQ9Wj0X5910jeyeFxuwwNIDQZZfEEcbi/0lzYVDURRDg/dkp
nIcWmJiyfrun8lXwEFg7hw4QH/yYg3OxU5zyC1gD2dZslDa3Dq9rwWtcqzsegV8a
muc0yX/ygT0mi3eUaZIiy2uKxEA9Z+3J1+Dqd8F2vPoVL0ht0abs+QKsGet/c4wv
UGFE2PNOWTW3e2B/lRwV+GIPkf1f6xu7sdKZKI/sTMdHrDcctO3OygUmo7akWmvz
DmqBnVghVLMrFr+8P011zqTaRtBOwDqjAKw/dkANbTpxl+S/lBc92GMyzGnhVXgC
n4MJyrdaSiOUZRDlbJsk0dSFikhAtuLYsPW/2tszMy8JarNQj/x2+kZ4NDxg0+08
91k4UbHa/J6w/KY/WoYQoVKLEIVR/gqbW9wweAbbpn0dhxf3A9M1Ks0Pmau/NRqA
Mo6HKLydZ/InViwu2R99rfeUW+5bYV53YutBqyDi0NmCICanXbQhDYrIXAq/rrSV
L/Wgvgn9EJqQW/dlKNyzpEnmuturjFYwgCSRvCRQOMSrleMQXyTWWdYaC9SWZI0Q
lnUY1eaCK+aybVEofqnLuUm/IwFpfu4KTT5KUloTe8MW9IKYzp094Hr5WgzP1MvC
gVYt/3GV5EkzJWLyrrDNmbJqEJyBSDkomi17qrquk2tmOU2xGc48PkTJ92E5ut0y
ziJJTaxiJQg61tNqV8CiOfG3X4YlH4SVjVvB894gKeieQHeARbn2fsegDOK/L7zy
Lad4144eYVEXzUzI2YlCO55bfUNbaRZYBt1zhjx/rQ7ac0mtOT15DQTvHiD8NTGj
efxJGimlP/syAuJfF97NUQYaa7vWoHSux+WL3dUf7ziSHww5AW5PqVit00FYOD7q
ADdsUNRd8A7c/mx14JVtx2pG4xHxG6EzoMbHtlfyTb9YEch0cvxtN2hrfegzdhAi
gsaaaA526FMLTL8DSboioNKXLO6R+PXS05x0B3s6WeQHqao++kYu22gg9Q3ZKIi8
Y5WxkUgK7w9DgSpPxfGMogkauyC8V2weCwBMm8uKbKnyBwL6cOJ55l79y/oa/rEe
69rEfGEESK+RmvT/26GF/jDD3JiiIW9D53XFpeIiOiJbTwWEnSVngE+MHxcoADe3
z874dQImI5wgGgg4fu0JG5QQQ4iG0aM75UYheyiUrniORjLL9+/ZkLjCDL6n9D1q
/+Sc1URa9OjGYNr21S4C2UhwZMPJP1/RPyfwar+eTotdN1fD3wVawOGcFuUVJbo2
wcmGFLI8wNJIrSYQcq29rTGB4X3ZTMLkAhp4LN8z8vdttYIfJyeqvP6XXxn4EVsv
gcl7JxbrwgPCujydb7RqJnV+ZZNUBUwqU9Qzc6RUdE1XBESPG8rvgWD1YYQx4KXR
gsQFB7aJXz4w6uI2jm/HM38MXlA4M6+o3hNX/LtMTKQoWMZOGRK6waddTCDKI1md
757SwQ4YUoKTHv9viYWApEL87M7AbgLhk4pWE08WUBHwTKYQBX1za5tNFojMb0DO
WfNYnMybQfxa0ZYGDIbl2xVQZMuetkWrL3MBnoDM4g1TKoANYplSqSSOfy1L6wgo
5f6fgP9HADdQDt0pGy6+pvBsDCqhyxLgubGS56MeXSSnzROsYJxREWuaZI2Nbvp0
kBjw1P0tf3UN2vxXXJKT+gmg+51k0CXQ7OLzUSXzt8tETIAKmXk5C+H2nLJ1GSCP
zXfPpEyVtHaTsBWxASlFgcyjFoYa7VwdHC7/LtIdGZ36F73y2acp3lRkSogaNY+x
reTCTpoZHbMVr+1G5ywOOSM4zQNzFfZnBjic3jwyrbk218ADkIVdd/35vdvCKLry
Ux5d8Es/NjeGKKm8fT2q2U30oNXgq0KSWgmsOI3Dxv50tFSftvnpiPwb6tPWyAwY
GKn5Trz4wfV0u/JkV2uPGWe/odrDJWMs1Lj+dYYmeMRzlX50f3S9QrJAETfjHVHK
VeUMRvNG6tOvdwsq5NTjOaOWlD2z+kdJ6NERTPFYWbuvaBmWX9PLKwFMSS4eFu/Q
7jiSkO0tNII3SZKMzFTx8zJus7cjqhlGtNgdMb+FZoKxcGapg1ovQgNAdUf6uW96
Q6RZ4kXoDNr4ljdXpVOcTKfWn+GM4BjeaaOOYA3f/5xvpJP6KZymN1vZOT6m2Q3J
nyT4BKh7HwsA4ZhJlRvGMsW48AtgNIsjBJ7G3cnmiy+xp+iL8YKeKbnf+MHcS2Jz
0rjc/MI9PVHtf4d6wOzq05e73qkYOpY8ZK6WFACUV3DC5uwYaYAigs8Z2P3yoasN
gmPJ8jA1xDfYWLC2O70vxWPPPUZnZV6NVRikSdWlymzun6kOZjsoLUeIdtcUw8sc
QgzF3cKuLHrBdobfvRLIfnJ3NcARrvKcIjcesYGkl+X4I1gf9SfLDMe4/vKXiYPM
YfjIZyRrdtc3Mur3xUWXG9kbASZojt/xW+JBS46i5/oBsqzpRTH2y3oLhJaCmVYa
Ro5AnJiF9uGG99CFgtfauAndZTUuafQJbXCVsmcK/mcvk8sf9+YG+FDMMeoAJhXd
FCc/Qt9T+yaDxuWmxuHZUtM1lZlkhiRB3ajZ8AuUbMsZ2JakHBMgMNhAwfeFK1lz
uFT/4YaICNoZoewoeMQYk5aQA86AlQPzMZjIkcJa1Azvn3FHZPq6vtN4STVdcSDe
Ua7D7QdOSTWmOI2kTK9rLq5nT0QpFytsh7kSuPky7loYcTokuFurtWdhGjUIChZ9
cQOU9emhXlsi58lTtZGcksBIYIQ2UineTA1D6FH5OvzSwV+DaH8dAk2XYvYCcRFX
fxf75is7D/z7UsDH5o/HA7bftAvOJNhwT/WAzvuzQoqBDq6kBJ2Oxp7bqZIllEn9
r3lLxu+A9xRGVgXZ2sfr/NJWzIkS2PX/EWT/1fyGpySnopJP7dASYTI+B6Xo1BXA
rUG3qjzRgzyY9yLhBvUuW4myg7lw1bUHMqqeNDYjUGcw3PHubOCa1GbIwNWwWxDc
W6js+oYHpKoyK/U9XitOXdg3J9WHSjILtg4MaR8XQLJjc7xyX4K/dFLY/TRFw/NL
g+PEpsMOldZRH2Cb423k81OMJ8oDG4kULRaPjggOd1G54yOIzKuS6lJPfo3PjRVO
50iQpYIx88VfVmtRApNFA5zWWqGTkjAuzAZGu2AX2gmdZdVhPX8B5zu7FhRI2QYN
PPTxCbwzYDFA/ADcbiU9v8VQXcx/dTy4A7mKZDQ/K3BXqsEEptTNUFSVtYtgIv2v
3VDRLA9UuMzyaLP6lDhhqqBA/4UUlALTdfLjxOo+0i2GVKRNBLtQ6XUFGdCJ1GNt
CQR+MiCGujSeCd+kdbHr45/mIvz5VCqMwHefzSQsuJwWzdepcljPaBpNjYDtCTny
0pKIjXSj91WFTVPuTqUpR3R4A1hIsnXPIMGrNUiHW6ywT78R2m9UDrQ73mIJb0T1
hZrbsg9KkASWE8OCdIp7L4Dbn++1MOZAO3WHMfyL1e6gtcll9r+B3d9Uh9l6KVgo
5Ws/YySDHWHO5h1CBnHB7o3QzS2SJUIBmPR3mIe0qnMzzztuQeBdyWuVl/oV+Vy/
ymTTAYsVzDhpubzv/iVzF7T2bzX0Lxa7HslsbwYZJ3uXyBfRjT8p89kT2ZUbQbfg
MfHyMb1gQRtNtyZIYD3DNvQA/hVw258r+u95Qy5v/6iBMqSaBinc0m1QAFxBjRpI
/cv3miJD/h6ntjVytcJekhh4ux2tYveM7LCRXf8/IIPrh4Ul8ZFqFn5+n3HZmsyh
KguKgnY1+2257oyX5GTgiPf+Asl6I/ikedtfLQYarkCWDd6upxuGcDMMvymZED5Y
10b3M+cWC9y+uTI6F4K3YrMgrWAEsRm+BhMoWeDElIexRhELhJWy9Uua3Xg5NiyT
s6fMGxAqih+M6fTNkfd2pLeTXiuzfyYohLLyHCQhs9cqnOfjr7Gqv6FlxdpNrM7R
mSDhkbz5zVIpC3d4pbQC4xHf+D6Y5nx3SS6X84LKcQNqgbSCdWhqeFi1gZQxTxXO
PTqeSmwL4YrtjnbXwxLfeCR6TfYPFZ/MviEinEh1DCv41Fo19wb1/ierUl6pj1/a
RTKbeEriOWoNNnWS4UigawFQ3Qp452a8OzAr0c2YPvSq1X8BivQ3NlJhSxIDdpMt
rrDyYc24E/khmxejwIlPbTRnHF/IetVenUBG5IfUDhAXN9bxv7Miuc1gyrFUmwwO
0kBhFMG0TfblJGK1wEkPrU1mv9yNUESlOB+0fw20noIMkHOXjkaQu9/67x/a1ZLq
VQjFi4rhVhJZTh4ETr8Xav2LpHTeaaU0L6e64rJPYUmkeutUdux8nfBeXSxYLFur
j8NXbBz+nbb86u2bTt0PbQm4IiPWSKSdZQn+sojgBiQoM2EgpMLa5QhDBLdux+BI
Hb/ujs25PtRZFuJwyA5yDoRJCK/1IaWrMz6kHHy+IN2vdRjR93/XntHQL3E1emBH
c986ZaDdfylZuioYVBhCMQ5uYxiRwaUnueSSl7+WYIRY1zr6L5MGoYsHyMObfaOx
jr+jh+1fN6Yvkp8rlrpsZWKr5iQVQ7vXAUUFnqGCiRh1OTTqdggEZFS60FBokEka
20RX7eNBUhCBfwU5+wAjYDlQhoT+o6SbMQ90PlKsPJdMCtreNfR/ZBAEt0L7j9d7
buVSLxgix/XpRWcMDBMyQ8C805JqSbWmMruBVFKnIJ/NaXEmBqeS+0THkvo2Tls7
LZRxGzjgHerRgvLtVAzoizSmtzIt3M9OyJinuvAsu5faAf6fzxPQWuNv2PUsiELI
vt5kTjDNQjNGfacUN3FWvVxA7FQqsNT8yDqzKqDjq0I2y0ggRXN6OKDYBiqus7ZS
szE0sMpy7OHVh24i9tSoV3cAn1hDEGqchfl//XFYz5ZzyRSBVSM/7DK6wVaWyqf9
mGH8AFq/WJfpTqAVNFTkk2fq7cqPZYfP4xy1va0obMyzD1hDG5WIr8XpQGkPCWjp
Tj8uX/vz5Yc1z7AlDbYpZwgaqddd07j+SxtUiByqX/GM1LKG+dl/1+VbEm7f5rpx
i3I0L8puJRvDdKQ71neI7PWAxFEFnoxJX8hBbeSCOPdOpaLjiUGlk41eIqHGYvk+
NgN2URGdD2phcAI3p8M16gP1elo5Bk57cxTsjwpAbvJJgTPMrcN+AGCOg7Ssj14F
Ohr0yt/YAxoTC6nKb4JJc+dUnzMclMTQ7sirHQ8vg/lLKlc1AdzzDP6uzBZB6i7z
ujBx3ODrKmAFmuAYpqtC7/LD8X/uIcN6W7uHe8R1/uG2MSCcn9/7qdLBGqM8njmh
tFxcR6iV7SCsEYGFgMdTZiHFeXKixvJPpBXzcDtMugMZNk3s6vnx1fh1wcz+Pctr
kALfbQbfoO4gMSCQGP3/wfln7+smtMCcpOtWisfNjLOuoqOm2O48fr/NmaTOtKmC
nU8vOTMGEIrG3aFkbzKHGQv7Zr3WHhkAmyeitBOJkoVqsH95e7nx+o8oa9mWa6p2
QzzWJ0VsJEOAndzf/fPZ+nK5swPnFhx5szIk0HXUP6amESH7y7fRmTrXRHojYr7V
bj+6ci6nSX5wN1tTPJuz0AyDt9/ek3Uq/FwKrOEq3vqR9pVrkeHYmwv3u+IOy4HF
kuuuDF7vj8ZfYaZDOqmwWI5murX/awY0zJWviCAj3bTFEhJVpD/BajgNnFstzh4+
46bcHPdIMbiAV051dN96SR4JkL2WoXkyHKxH09oCm/xdIMskjRNGr8oJbD+rCRo5
hcoCJ3vEwMy1WS75IRpIvENFtJ6GSC1J/uVETmw6l4UEbwN6I1BkwmcP3WOHStMj
jfEgsop08Im2HEw8znd7e1lad/KCxwy51oUdO5ABFZI8YrPLDIPfDzr64k2tzC26
edQHoIbjK6RFsGC5YPdzzEVUSwFBz1ptL3cxjBGCvEUssSXX75P5hGFDxygYcMme
dF/pCgctmPuS4rdhCA/d/LjHoihi3i2GmSLT4i9gMiZXYG9Zw2gnOSrgXdlIqmYH
yfaMqc/6vK1sbx1BOyOk+M5khOmroZMLyJ/q9kHbGhkM7C6/Ru/7VfAg2UOfyyRL
yJLXi5345/f6wvV8aWQ8c+vMToG1RQbn2r8asfRnOESofx3D01Bvp7SGZGcNZ4Vw
B7TElA61Byu9qUEixYPomOLAmGpRn37JovgQ2ftlcZ1ap/oJi26V5YndRvE1z2SE
iQaET4LBZhXfsL1BvTBlFa1ADJP5uSWxrzKSt1QxGkS70K0BAU0H5UXHjFZ1duXQ
7o8xyWL412O8M6jdiY1Prlm51BDS7WbYtxGkfkABu3epj0ESenGdNk/j5ChFekju
/CEUZajNJX4NgTJ0dU5iqC5SVIZZnMzwUMvft/C2aLSelzaKtSmxlPafWnDqK4p/
tAG/dCsfmqInTPkOu1GJe66xGpBIavkPfwn72NJzW2w4TX+ieSiZLUV2n3iARQC6
ZqdFntiDH2fY3rYLI1LFXsUnkK+1UJBbA0Q48rb2cdFBVASqBs23FOifTMCAQ+0G
azDTPScqp1IekZTqV6ziIhMMK46t661oU3nMNgZnkLtitnJsACnFckv1unRye/L7
rTzlAWGRbUwSQXY4UNOoyX8WLoZlBTJi1IGymgFgEtAnou6gEwqBCV1M3m6Q0Qn6
M6T1sRSQtHWAE0fMZBp+X+v9IQHrLFvoh/gWYt759komdXAvV82WO7IWB1tAHU+V
E2+9qIcsj9HFS/e69x6BZXyJYaKAnoBPDILZKkfhH3wP/c7AnmZhsF2otkc/Ku0W
OhIOoBGB+Sv2kAkcBfJ7bxrqVe40pfCRXyHPgfzQyCimlTz+OT8aTTHfWNDPsonH
2eorl8jwBDyb4DEZCqkQ4RtZmLXa+pHYXAkgoSHWs3VzxRrPoDX2nPWvNdGKBsHQ
iH/1p4RLGRhpTa3Y4RAYYXLnVIoe0qrU2+zx2WrZKcJcaA/6tu5n91gKyerQOaK7
ECrK+6gE1ADnGNIOOXPDKo0HU6bYoyZmVS/GQOlWMkfDfwl1Ov1ZjvxaUha/MTMu
wTbInx3Bxvhix4OS0lOCTUmzf8qH2YI3UjivI5oNPF3y6lNmJ3syrm8NQVfDzkhv
vtk0gBsG8/BhWYSGvbLYl9/yOValVRafkcCYtuoLKtH3CfYMTlTvlNQa669HLnKb
KcVlWNJrMbvf/DD+/+qyYD5Fn6cO5Vtd1y3G9y7FXiBqQELQwtma1r07G9A+RMin
J+4R0hMXCLYnWSLWYHS6MDnAUilR4G8YEtdunlM2n1w/bTjvXJgXLMwtU8E9rsqh
Hb6G4SCqIbX33GBr3FKgjSHCVmQ2FnpyDKLxpjszcv12oFONN7hGSBTQ182dq8WU
q2kT7EZP7A89iHYJsJ81n+oz1/yM4lbg3cmTdP/cuuOKctBIVSU3Smhfg9cB5zCB
+dkqSp1pg4BaseWaqSlfpBtLhYSWYixyY36HSamXtajEEV9i/pryNkh+J2o4N36f
rWD+jdqdqhYV1gm9buPUVW8vbdWYjSxiuffbSjwp+wyaFzsuMEyA2Zer/VqK/ght
ZInTTUCZHd2KsLkIqMPyqWThGouuBjyxkFBN5cmCa5W45VakCTZygO5i+c8a5/mw
MZnZ5iszGFsAM2mVk23IS+ovN6jJIRkumiF3QUfOWT8XwnnFNq4iVs8V0GnuiTba
WJEKSvoVWNo6BoAr0Bu4cFHW8OBqf28aFZpyN/fTzILRNfjMu0TuFWoSuMrPKAgz
Qd+ZhAJ3bpf5HfIiONxstYg8zF+LkU0eCrYmcPJTDh0TYWB8DzscqCbvXTcNk+fJ
uL2UKcWOVL5+bxQbIBmHhIASA3fqhcxiIQZk4+xntBjxk/+dP17QEJETh97+GP3x
QwCVsZxgef5bhqc4CjxDqskefn3vwmw0slFBMI7LL1KEzFwj2pR2BRS2iGNFMJaf
txxtoCbknz2LedCs8fTBRfX4ynWgACOnFYNGx3BGsayBI7BLcBmYKREq6VaQWowJ
d4rCGKiOfD56sO0bERURUrkj59fIwL2H7jnBL7Rk8+NagqJNT4eMlV1Fh3EkOkmM
nCrqQk01YWXJovxEkEvXbJy9eqOzIA71hnJHXhq7TLU7ci83N3x9Zw1DhzuChOkH
I10CVCguJ0ctMGL1oOw5mumvbnI+RMKocfG3wwK8+K6XzGUGy75+5WxosQ68Ohu1
+LCak1ArgaVOrtRdg1LloReGCtGdQ5ek+DOFbBYMMYVMDrih8fddF6Mduow+1ETy
BzLhnW2KOc+iTngTWHZYlDfHBKtV5P9A1DwWXnj+cV2MPvFnOHfFpIyTrbp2Msct
88BALmpxUHFhe/xV1ez1s751+JAZjhxCV0dWbfsovvYq8REvarbj2ozbA0rFlL1p
C/XZXx9Lu3sAEbkfNEdy4n7oowpD0uqUT3jErjrHA5pbwpNIgi64Fh7LVNdp1a+z
s7+QoznCMOXdPvg8nqqAo3V4hP/5x/Njrdd8bp+Y2D1Iw3WO2R2GB2u0rV/Bvyxp
mO2jPkI39vr9QWgZuqHQ8FwbvnRGIwDJ5Gv+lY6KAckWWDlpJO9kIWMsWK+ym8xm
3t64LhzbDt/L/OYhg1sd3wHiIRzDHVkUFDJgmkCiyDgePtB3sXqbiCdpSe1TI+rO
nAXk7p2yBINwIzkt4IKZWb5frdvMQyhs0KfTiZTTRwEbYvpSQR455ghVLXbvy60B
Xs7pJTyFHWq4cbJv6s2KBOu8j2L9p5BTLLriBnBwV7nCXohEEz5eenvR4pLtN3Gd
skZo8KViZQyeLjySaksUl2nVzRVSaD93ycugwKqtraN579uiJu/dIs8B/nLbkqGi
Sfe/CH0MVJHDmh6Hv5qWPnW95AcRJk5lPBQVpq00qaEualyO0ONds1UcngwedgWt
WWv5s0JORlJ7aJLYR1u6LuuTgOI7vk1WTqW/KFJR20Tl/BVC/bCKDHsjotPcCo9f
aa2oTwu5JZHk/vHl/+NRgRsSH8OWeaNbh/0twOX+kM7dRwHVfxcX71lXQjyMa9BY
il1Ap3d57HY+AslP+maqVhvpw19/IE89+iNFJ5Myc1dJEV/2G4/Khh1B73tVN5mn
FJ8v5L+A3XSoJ/bdewkbsp3F6P99IL6FJJD1HB/XEk+ENWMZh5KLD3H4WH/s6Njw
2E5AJ1qImguhQ+X0WkBhgFs37xiw2c5RCb5f2dhkwYFvEUV3/AJxDHdnY9tB4a2Q
ermEeYwpc5jnmgjW/CZWZV/zo4rNgb1v5dJtx4PzpOZooGovJpovymZN6kz4lRlC
9AlclZBbFOe4EtlaJ/KInXbSqcDEx31+MfMzhcJSDkWVuj/r5ZY5253OHd23NJpI
PZ6q6YJW3LHTcxgp11iBJ0dAOS2WhUjys0jdYcmL1LXCGsNqRYsPQZZZr0lSLOS2
1nYrqjlHcIj11GMHwQLURfTSIuB8dH+7s7ZaW2Ww2fglyGfxR2ja86AxWjMde/x/
p2MWiG+pTzecEAnkgQAcMDhbPc7hFqulzP3tjm/qWEAd3fRh/Quo6Xmoxs6lw4mC
TCPS7+YUHgj7QQsvYuHupGGEVXn5cjVSdBxCZA8V/HZLBfQIEOuES02mmiyOIATi
q3gCx8KuaNROdjA6pd0Ccb+Fg5QBpbLYl5Z0c028nG2LjU9BKOlZU/WLvsvGJrQR
gtiQ5npVH1QZ1rbaovoDsGHee9wr1HW0cWmJbmQKCRVx5fT+OTKPniIodP81Qv2j
1OIM0DKTX6+A1wycndRGwWhXE/QmtL0aV1SU0LtCXNIfNtTr2MWwmNAUiyg1lgBp
pM3F8+aLZFvqWNfCc4MrGoPujupWcpim61IScSPEnsCJUPixA4ZjkOfVrOEQl7vg
5WKmqy/Ct8F0eC0YeCYyP0KUB0i4WbUM87EdgI+gmrJyaonnOYp27fIHFRR/6cjU
70GzqelcRjNyjz+w3o3Hf0HAO6yHgzlXsdUEEzN1vlgnD2Kij40I6T+wGIoqsJ9m
EPpNB9VbN7T9YggsgHbMO+MABDhYjltThOM5hhyC6mdYnj3tcIOrCI3m5pt4mqfv
mA5fit97eTxNsF3Xe+952WVGS+48gcjuoi2nR6b0ltKOZQ40sDAIK2yFNv+dPjQR
FJF/oQPTL0heKk2EdRTDdx8gUOlhKhbttfBRXFY9e0H/lUIro6MPdJYQQLt/Fn3L
H2L/8HHQtoqMsUC9ipveiLmjeYVzHLVuSL1zqr2GArwpJMXmSvRaeJE9mBueZOEb
IxBSgOfNHE5lQds1lPpJiQdMoVoA7sXIOc7WB/k3Erp86HPaendgUCNdSuVBjQtz
tlho3ZFPuLB5PG0RdM938QVwKqc1CI3qx1SHGuXVluSWIqZNg90vQEd7K7UhI63u
z+zkC1uDPTvKeVf3qqbu1O7UL9Af8Hc84k58/DRZDFVah41IuETS7e0Yd+FRlY7X
/DW8xOrIyA8dm/ZCN7D1LriChpSZl1+Tf0oyzELIq9QMVhJZ81wjtEzQL+pc5GHA
aeP74BEhRKDjh+d3udKG3Cy0sVDih7eKJwKh8O0k8NE4XL3eIQ80N/w4gancFhW+
/Ch6YwOERpxBK0rwva/vF12Q69Mwgpjv8OdmkibK7MpwZEdalTjwQJlg5iomeeaN
eK1iHTDNzVqTmvw5smtlZLGkCGasOyN6FAJ8MGjMkSM2EngCfcCiMToN55tG7fSw
AMV23GywIwDAuQMumlG79iYx0wFZrfDxBSPjxw0ZmuvKj1L3reNiQzHJnquQ/KO3
3dIcYV+J9euz2qoIx0thBkl4inlv+7pKV6SML/Xb1m/4iUow3ljxpVhE215jFtLL
gCyOPv5ABnPbMzyTEPmZjU8hrWzfdNCAWBVNyJM6xbtEKklfylyreVJk3HgiM4v3
Y50EaikdF4HvLzI6xTjBRPlQ2X5r8BXb+0PRPa0cCz+1LIie/uyROw8GHIIc9cax
Iy1Tnve3qROvx0baKwBhd9rG+dSBBNKWiGXXqAGykqulNR5gmUgkpi7ExC917uFq
CNJwJi9FMifgFz4IVVggZOOFPAOZc+vn8HQbI5/E81Hew/bSGXBgbddjS7Yv0Udx
bVM5SPDGZxc6FTGMf7kpI4P9OBox5aB93a5g4Zw9nxtKD7VHRFdV+uzpZSdyWyX0
DhajvEV+/Vp1TP6HSyVGHQeWeO7pGBXArZUbUX/QlG6NPQs/mquscU8nauSINcMH
CdVOj7y0hvRUxAqvvOv/zLkAMXSyt1xTCSM1k5wbgE83hj5bhd/NNtbaXzcgMgS4
vkujfW6uePAvmqHzh87Lipd8AwzMCI2gikam1FZuMrd8HXpt3so/Y2dcSKk2Wufc
53h5g2sI1wtjWZAeK+Y+RN7GG+2A7fY/B1+K2w8EvglWuRjytqgkQV2OJQilmfYB
6UJPOjBoQ1WWavXlEoUyEswyqEFdqTmEQFhvt38x75GojNvYdiIxRYKYP8VqcAJU
CfOLjUJ8saHL6QNA2wZPRJHhk/xYR29HWF30MrWr4VHDKc/c0EI1MPNFg7SCtpib
L4GJMohROn3blXDZV9emz5wDR21cVFIj397f82Tl+de1BTeJ2TBEbCKSgO7EXkSj
CovpGms/DVRu8/7a0lCtwTMr3v6xARqEI6YDgCVi3ZFfFmb/oD+3Jd04d7kwvcKy
slIAI/+UyJlosif4y0+dnCL3vIsS3Uc3rcKuVjg4a9S18+QE3dHjaHM/g+8IwCFC
9Jim+C2a/gbc5dHgADMI2gcbtfV2Gg/jUZytk/9OkJnwQwNfiexr1OgFbUetnrln
iJIhNVs8GQq3mE1Cpd5Kdvj2C1u5tqVys5L1aFfhRcylQvSgvv+/lbZe3E5StR46
J1b9L3WQL0VCZtCO/IdFkbomRVeo1uwkAW5tOY4GW+My1aAJP1rv/F+T0wqdbXbP
riwQrfgnxwWMjaKRsyy8bgvGMUzNZJkyXRNYSDj/WyeD9sWKsCtk5/2hbrVsM7Fr
C2e6evqJ1h8+KNZZXTggVpf247I0ijpeoo+1CDYe86Jix6oNqpHeFFe8vO4SJsXC
FFLmYFTfhjASInAcAI8mgwQopmHBx2wqq/KYrlg4J5UqWkm+Wm5KFUhVoTtYH+zo
79cZnAm14LfesrJ6RVbvzZlARDLVe7ABvN1qLUfM0LV74pOsQJ9HtKmCo0FglYYi
EZrvcZ39PrTj/yckOvxLt8L2dTb0PfVBOFiXstn62yE5uLyp0ZUO1fd6cZqDnNfA
3pfs/CsnzV3gjEHF6dNWYu2d9eSU7GkFEFEGm9HrHpAxlVZXoeSzfZDaOluFJE+V
dunnD99ZOteOjIwm/V6JH8PZZ9fNlDLSAzJgMlCkQ0n9StdbHqpc1MWlJeD0hQmG
7+QTZJ/Iaz1qMCRoDnI6NDjaKVaAUjL7AqIJ5jG7hcXtuaHkGDBKC/fXYQyJXFnD
TDjpzB+zQIphaJVxRcPjx6MicQiLQhysAyhkYV4By2KRJmppFb0kgelMDla3MgWy
w4CWYDQ2t3Pw/lWOdA0WvuJLzzwxw0qXRhmEHHiQ1y5u6qCsehhIuXBYEUgihsra
4DCdI7OX2Qy+pBXr9MGw+ZLOWDjlLUXqn67r2uDYBzEiqqO97PhL/RxNCHIErCtF
1e3LVpgJffgFD4OzSBKnGu5ybmFhxIJGHL9caPq03hgq8KyqaGBWJolVToVTnm4U
GEPtVUsJfd+ezzZu7IkclCyaVil51blbVzj2ukoLwh81FzzQlgUVxJbPwtKUWiRa
GNtEajg1T895kc7u7aLtoFqoYOQom0hsyyiBBEGd17Wfsd0V57h3w8jPfPQiZ/kC
zMTaVQ1a8qWJ3OOxjwwrdN5XMFv6DtfdWMT79JLNElpwoPLvIRJuy2FZNxdrjzhh
CYqg69P2UzO1+NRUBCkCr1FrsHng7h68Hvx6YXXY6FmqLGT98yYbKyT3RE7wAebi
KhdnJTEG1r3akytzfuQ+WJKRtl2EsZOUzfP5FVQwqdc41RSLyf2+5bnNVnE12/HF
ungwHK1NAYs+2Sb1L/GAHIO8z8K/JkQTtDc6fZ8HyLAg1RVHDYt9MVZcR0clzosW
qrwaqmXSEvEWkW4ygy77nufQneZFAr4TqtEM+FO4Q49CKOxte93jTGhyAhs4WSgV
AxWuc01heQuqsspaZfSJ6P3TTQ0GGB/1ZNEuzERm56E5XMzdWtPesHnRbf9LXUHB
J1m0Q4aEe71jykcYB/nRFshgNeFys7vk26mCtCV8y4k8pCX/e+ikSq/NI/GTsxSm
MFCRQ49SNEpOXVf4YngT4TEF0TAoK6ew+QaWpkoS/LGY2qKjLGHH9T/AMRWEy1ZW
Lc9F9FMnYzAz5rgA+hcWwFVOpKrU/xwC2hOpPkdEmhXlS4EpvyqiN5qkocYCfRrs
0ZrZgyoMv+VAI1CfPIEu1ZGETj1buL6Py9vK1ALioNC2hO7AJe/azsn3JWvpcGWU
Hu669dyFYtSu28yBEkHpNKjJEf1Qx1gqYxed2e8iRSf7rLqK+nP6FI84kuf7dm3G
GXv42j+BxnlPuuVIPeI0z5QUKniKAdeDVk6DvrNDFyBJf2Z6+V7Wc+WWqg+s5+Of
mwRQrywdMHR8HCeqwFEUdd3cccdTz3nKqF0h4+g3B+9vSvBT/62DyqSt8H3OdvZL
iONfGBGqWIZfFU4MYCNXZJyhAUOwe/xDJmkq2KBLag7KKMFDMt/CfcBuveBYrVWS
EJljE6UAU3HJIh/ecYLChGFpVW2MJqLZgqTKaKk5bgUF2xEs37ZWFGBNTXSLFRFh
1meI1j1C8r6ddAF9+BQdea/5480aW63q35g32yLmiwAophCWA5vpt2NsbxUB3Vic
F5jdYxbgC5uGLjaoGYHqAPaNk7oj//EUJee3irSmHwzX8nt80U7pXQiUXI22TQrn
duUslpkjrw+DYvr0LoBhcUUugjQZF00Bjp3EEAxBMUtUhdmeGjeu0fJxF58Arzy3
P4rxZ3LxJDo+HaYBZpvko/CMFAz0oi8T94BOHUUWKU4huo6yfaTmq3qpZZ8vp/u2
BGAdz6JgbeUnIib82Mjyt5tMCYpd0M+xs0RXLWJ/kDymTdrPG1iI9m2lACcNRB8P
mPbvwre1XKv9EBdw23xNdYBi+w9xTy81fAwfRv94MoqCHcPCKKcZrEIEJJsIOqZA
lFf1HLVQXG+eOfKWdSngCMhcoKVGV+VgmCJMK6Wfcb8=
`protect END_PROTECTED
