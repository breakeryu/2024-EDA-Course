`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+kmzqOh4F+qXQC9Xp+nwe+Je+OikMKpDc4EL67LQAlkE0IHK1PY4inQm0+QCLcbb
ezV6gnxnIjoXjsCJLpYMxLY6p5qPARjhaobDlN1WijUDkCfzxUWR97BwklfAUSGY
6e7x2K2/E4FTnrXrws61+ru9dqLX/npJ0ixPF8BFSDmoGpCwcNtTQTqSLjwCfuxV
CBnRX2ZBgJmk9F/j3t7bPgWbZTZlvMzKyYDrHwwa3QvrKGPt2oWp7xT84q1kLDzt
gAf9lcp8MwgKS1xm6oKpLeXGlIxVEU8ICawmjISTghVskuQb11f24ahAt+5a8vKh
Ul3SJKMvSeOlhABVnhZry4+7WcWzOs9LRd54T+hdfrZzhLdk0QERxjuM/6yMlmtg
DaLmXMcyS0Lv/Oc4KAH6gnntq2q/TYjArsH/MTOCYbQbOpCV7+SEXxQpmBMqxrbh
yS5XZkYf33cecY/nqoWWjMtCDAvzxp0sVGMjhlaS8UM6xLasbdbD0PF6IYWrdP/4
R2pze5lV1pWQb4ZbGaifIFncp80UzdPcDEUEnz7YEbeftl+1Mi+NPzYpzffCqSBu
BP/8fFwaGU2eMhj5aXaBWXCM0kXJtsEnhcvxWTP9M5vYFTR0mK7j4jRfJzVz1mpe
fmLviALF2b47+CE6Ydlom++JZMMksYEfKbVjHL7N43v+mp8l+itjgazsjxGxkaEj
EXEJXEDCRY2U+O9029C4Gg54JE26qtBtVgO3aFdqcr6xANctKFBb+QmnkPUk0xk/
4HeDRqRFbeTO2RdyYCo4BsFKqMFN8uU2l7dGy30MOnMsA5cRLI9UNMi0CIfl+jFF
Fj8xNbOODakyeoYJGEaJJt2kHIXdyUsTYCv3X+OyuFREDhkz3M6YSuyTVMUslMEj
nSi9VfIjXf6H6Q9AmbCZYKkXQf8/lDxqP02jxqMrexmPzgKErwCcU17R4GMoxKF0
z/LE6rUze8BX+8rlWZYUPqzYple5Ua3PTW8/XRhtakfyWPk3GLeGyAAWV2sXwWHL
v+H2qogPbfjqix3l8ZEiPK54GjLbjhUd/KKqV+G5nQmyg0/3evbiVZczqcVpSUDb
c8QiyzxHw7CYQg4Yvhp9QcyAPzhaOXDuwLdRLRBZCRRp/zbC65Tkrk62vcPM2ZA9
FGPPDgppDgIMCE8ut2RijLzyILnAJK2qkTH5yVan+eJ7Pea20aGnsF1BsTcdYwtO
l0zQ0WrHSrTJC1oXurCrjSvV7WRbk64pPPb2ZX1T5u9JVyjPLuHfMaMuggWuRAPk
7cyUl3KFEB0IHdVeePmpS8WLTigBP1dvtymAq7jKW8jYtglG3HdSk6NbnCVF6kXW
maLWo3XZRUzEJYwXsGC8hN9ycZfpx+6GJGzgYrs/bDXXhM+wfCN+g1OfPMGJ61G/
X52M2IF1FO/wNu3ZL125ONwfjqHbEDBL4xv2MHYtogJb7gM8TYsmdU7ddZQL98GV
50kRhhuisRwlAFs3MXnf7SI2rTfj/IeUDCesuyP2mROrwIKAfgaaY5aEdPO3GwDb
dQsvBZH+9187PJPult+WpYwDbbnJyvV3cEl1NzgHt57uSkWpl7tRnlT6adHeEl1/
HGKz3r/0lIfzvbxHN5zq7m11qfcG60zlvaMCsrwdMe1R363nYPvfECrKYSOcFa2H
9dO9JfWvRKUrd+D9c951SSQP4wi9OgeO/tNdqToKs4SKRv5X4h5cw7NZme+KZdvr
CbaeVWNY1OcE/u9Aj6TOn87ri+PIxC8OqG7Wgrk+RqIbIlVRfnx5508JvsGBTgFM
i4c6trrJarTUD7nz5P8bcPDXyXOU/PnKDztjaf8Cri/YiPZU8Pgja4xqr501GYi8
dFPJnOQZrLLjpVSW6Tlr+XeA5WgFnbmZt2ShPyXB6aEUAbfHaf0QghVvLDzLoe7t
rocTAjK2YfG48r0s74HUUrtAq7vntvc4rP7bZT62TNbY6LlmWEBaMfBxqrw5yILo
SydQyZj4uZgREhl0iT7wHZJ3ThEKQar2lRr8fubSvfu9XpAQkw6RmPBQw0m5Hdwn
SFl9vztYMaru1G5/YEhpwIreKOHcA+6NSLAqjBWlJJpZKSbJItGVYT4mO4l3DueN
6y5ukEQdw6sxNVXisBj5k39A8/gYWl2o5osu/q/q77fQezXWnY7f1hHxbP5cwx1B
H2d1TCrpKEl72nRDjPztFBRdrg7pKEsRdmJbDYoG1TsjVwgCvNoPg691B1QYXGH0
8JIBS+SPQKa5l/v3Uy4Ck1xeDEqbaHQyJaVSeqqfiIKaOafkJ3XcpawycX6nXtxF
wps+4YRjgv59JJLMKzF4ppnyQS2qDxtPvnz1nuNOkDYEsr7hU9Y8/MhylRE9UOw8
IF08fgcwCGAGsRGkHcWO9yegmfceoJBVNVBAdHlH6GtxmhWItC+gxOQYtzFGdAXr
l4wis/01vPx+UtHf9ICKn3Dq5qrspNk28cy4ocyJt+LpdIr6h1zsNxTm1+N+HNbL
YQNCG3gjnIzUFK3C4wjnezBvvermFAI6LoJWGjgYUROGkS8hBB0H5P4i8o4UoUd1
EnmOrVaKfK9mMTZ4MNTp8OI0oJYN3Rn/ndXnQkr92rzOI60kgntgsIsX/QII4yds
IlogsMPGd04SG2kpWsaLEHkBIsF3XWxFHuVVgeRzZVvfGRKAJGqPr66b77JzpnLr
ASpIYAg07fBTzZ9FJ/cexscRRp0w1MvZLFNXV6Gjs90LdecVV4h7gWawciBOQRv7
RbXakrjNYd04Flh9nsVt9JADk6WGUUsb9bkLDaYXW7oRP8W0+Jj7AOGY0nZiFi7s
cPaLUdxfVE24zlAGM5FfYigLt/vTQ2y8U8gOSbrHHo8lG+E559gbG//Y+WqANVTO
wAZGP0WCT0BdrqITzNbEQU0oPxl6KsCnP9zy75mjat5YSaJkEOgED8t903HjZ8Xm
NtVO/3mk3SzC3z+W216uG75QSxlwXHJsrYy+KVoCxvNhnJmOP4EYKqYr8wsG+9LZ
Sv0EkEG5lZH6fwX2fYGcPqFkVpP4e1llDaezkHNOagXnGaQg6WsvUrh8Otjp8UIl
uk3qHD5XNXYgoF6LLii58s42Ng0Oi16pc0+2I+UnAcyem22qPGDtCL/BSowX0R0i
MyWHSr7bxbNSr/+6lK5/9HIrE5tph5GpNavwdv2kpZLrq6MzVybKa6Cg61lSdj+b
ugi+6MkIM4PXk8Dp/OS7xzxPdJoCD8bUd6o5dL+n2XAUJ7SaNTlvodgtVALlqsXM
MzUhYLZQhyRGgCzG5A9+FA7FplzL07euM7Kq0swpFdTUDuutfdZ18PxpfU0ra8oz
H5Ao70wVFcBwKcNBezW64IFedjuaoAOPtTQWdqA7yC+sXpZsYSfs9CmnzK/dbvlr
MrP27mU4pDtqrT2UBZXPitGm3pbedTcn3F9GuzNtfdzS1AXlYPeAvDewNcJ2NEJp
77P7QEbGQzVovsMGug+ICBrbDgF3TmLPovdZP1oYnK+jlWGnrufYCyhXSdWU0i5D
YsIr10WiKYzznTvKzcC7a4ONsw2JnpIUhjA7rSO9zI+99dYN0KswXtLbrasnOImd
7IpjeJ8jqJPu9ZRwX9XOSs7M7kHnTP+GDwsgHxBHREsNxpFNvqJhWfE4ntu7z9Ak
htyrRjCPxYmAeCc6xqgPnjjaQze5S1396RcdVlaqlzx9fIf9DYdx4EJAo1UJhSb4
Co44PxoZ2Rhzl3xz/oGRM/wvxD2v95WN2AT0hr5bB9sXJr5uHkLCOeY+2jBFEGBc
OuVg6rV2Kuodjl/AaRdQEA9qwMZpspmtC57o8WTjQr8jjY27ue1DceNWFXelZ2P5
GWpNkVj2bfRYLVcjZeR61GMyc+yG8Lr8vzE+/vmf83mbOqqmiLhy3R6Uwt+xPgGV
/o1f/lzCqtuJfOiM7YBYuf6fEf04+nKI/KTSB0XQZ70fzCokcDBxwThkABZt75ex
2ggk/aHow57XlzXgZEx7DAOdU9Rvfvl1WHNnY0VDdaM7rp+0seTZ6xTTL2tO17ob
wx0pc0Sj6YHXn2XvjRBtVVF/6Y8ncXaqsmA3Uo2x2l1xmkz/yWXf+2xbfMv0epHM
f3eQgqqBoxd1RqtUAJtK78IZwpBfA3OKTOFZLo+fAZyfWwYPwgFphvIrQHQJ4vCG
4fPBtVuoQllgQmF/YxRTggQ84CQclaWBEr18lfcP3c+UUlsxQ3KtysWQi1F/q1jl
nCgJznMbCwJ3m8lt5RWBS601ZwN+6KUrkUOIWJHnxhS0SneGSbzquWYW8TZVeOm7
vxCcoKNWqi+9O3gceHhAGw0fj5oXlvnMfMqG5jQ9wCv8Uitx6aVT3I/0c7TzQGyx
0DgEdEWbw4G/aUur09kahZ4RQ8w/i84fxAwdAqPX9GC1TcrFtvE61BqScXOgeTVd
rznBLiwrJZ4RtfZX4lRPmikrsXQHY7G/WgbQwMzmydRNaw34fXKr7iCp9RUfK/aN
PPuiet9WNotRuX3GzfSyOrjjm93YbFQuS/Yp6EWNSqdXu+xHUIg6JuFPXOkzkPkj
Yn62iw9J2DoVIUYc5jqS3Wnw6kaktkaPF+uve/fQO3HUwx7CneLLYUryJxkyDBkn
JEYg4+d7th1nR+pP958IRnLwmr0g+j7cSHlEwBO0xW9rHUfqy1hTldumwAle9Zkp
Sfqb4bppxecHypIXNe55QWCyT8dL1rNgcZa8JShYUMYbdQJ+Qk/MwssLYDgLkDUW
r5uDU+epKXGe/zbowjHVTOhP19ikQchLqS8MrqePmBEmDpQU/3PZaGNvTEr6miNU
XzyKWO0jH5ctQvSztXHGFbw5cxwoUvAp3MdC2ysjtGMD6jczT6vsgcOa6b4SfvID
cNs3DPwkZk4L+95ZZaIPglJWdvNbbc7Bx85s0qznqhNpf5sDVb1ZZdyrmTrIfgCC
HCtD5kNTxurlLNHuaAOZ86L0Di/td2TkfCCBimPpii78Z9UQZQQHc7Rk8aVaZFIR
CEuJkS5HKkl7hnZ1tKs1B6OsEAwgGEuTJgE14L8y3ow9ApJwUX7U0p/2mA+oSzPD
iaAee5oB6dUKcMVRl5pXcUHrjjqnXVNxlJujVWnoQutLNrxgGaGJJW1qGapQHrIN
iGM8ZHjG8FQ0zR7TY0ijE/+QnjcyeyCYtU+7vIT1YA5ZTeKh3/SYrfcCZVSh4nFD
BE4z9A+0YIYqC1ZOa9sqBwcmFTVft7ivDkmVNeskm8jYR7tefYzdn7OyIBPxSnit
tlrcjFhXbrr5L+VsdrIR/g==
`protect END_PROTECTED
