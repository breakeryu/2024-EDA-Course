`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UXN45k0u/47pX5WizNYrneiIZx1vasvf/4fQMyuHNPnfVU6iMD+CfLNl5uXqkekz
NxUpE8TWdQCi9LnBT04kQYtv9CYmqDI89Cdz2dNyJQwUZaq5wu5wpTCmrnhLu1mJ
ZtmaZghMai1oCXEmPsEwkQ6FSBNPJEzTak7zYhYgdf13n/LJidXuGWW7qDx5X1/U
Vp6NpylDB2dHW26irObZ6378GH4Pai/jaWxP8J8WWs1ZaIWYQf3CuHqJIHWCOKiW
x9vJI54AwRafbP0JTFBM0/4hO5QpjgJXHscBEBKiAmtwbHMCBf8zqwADdFVqDFqt
kjn28mHST1Nt0yNmcvRmDRptyOhEKxPWyU5g4RPBEBqGlGRsblaurnGly/RKUZW1
`protect END_PROTECTED
