`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7rMqvVxoqzgMN8BbZ598Qry+608+hwnPBU3j3R5ZHtBfYtGKCSXnXLtN57hMdZ/8
CUWy4GfBU9GjF27OGMQESn0Vs7P0zlFmYhHWxO2t1ZNBJQM21rxhEFq3z6qQoxE2
bqnLz+yTsb7QJ+R/Bq2TFC9RNeqNlNVPu59lCCf5TRhxPlrPmaL4OsZOEHd2tNbJ
geU/A2nZpu35vpUCRD3PjIw61Y3dNhFn8ppoWj0Y1cV8LjPXZlXMJxzHzSg0jW2A
pWYkEg73YorOAXMT6xiyeDt0Xun331u3m0IcG3CizAkXiwOrHEVFf6qrEibd/PZE
I8LE31Ziw9qSexQ7ESLxIXaz4XRADfNqqwALPloPmqXLULU8fEyG85WH7KvGN/IP
iKvEPv6cxrAOlglQ2PydYXOGEtrNXDw+zdyhYy3ZnEEz8L7gNoCKQz6x8HpTLSEU
1jzgEYt/T6VtuEI/GrooKINujXtqpxdJZ1zVPw6H8uXpws5aj5BY104ld+n6cs3b
REyHHax8GoKrlYXquNl9rd3o1RUkK7GJu84gdU0jv5HmkjO9uxNX4Fwf9qIMfrnR
fBbgDEcrsvuZp+bkrX98lwE7RgjFBQmyYVgyEZQTBhYXeDs9/+Ij6cnksdsCOnzt
TmCCq9U4AsMfKFXQ1Z62f4q8NQ/4UxI4MCKTU4zQv+LXlvf2CkZQn99PdhODD+tg
43XHPwp8G76xLnDx3aCiY3VK2HcE1eLz7WiZxJ2FpVhuVjq4lg3Lf2kJNym6Rq8F
oJnJ1je0KIARV0GDrQTVZqz4jSw7VsAU+KxnIzqJiiYgp++fne7g7icQ5/NKD3Sg
OarEWG9iHUyEArYh6OlMUidP9q2WBQ/2LvjRz02L3BpLhN8h/GG/gpKQPQlGk5R8
rQcpW8Ejh4Cc1Ejwz6OqACihqVWantRuGA1EKvTz1GcDMmMfF0eTjHgRTzpHgoWZ
zSz/7DHNWtd20TDEKXWwpeUdYB7R5wQxNSo1KNF7vhWtyNs77cyfxk7OckN2assb
wTXkmWTQni5C4C09CiLvpusO1qaUWyrv8G93dRlz5DyO9oCZ0X+43hVNGm6jmpt3
0ASSzk8ah/aTgWoD30AqL+Grf+rY8n7pyzOPYZ+A2Zx4TlfxntO0xj/VCuAXcSw6
gWmWpmA/HewTpoZcIffmDkmChKYiTD9YWvGEimFe+Z7qyaK4o8+gqQktecSFZMXp
jI683PYFQvcjvSI8nD1s7bNSYf6MbyYY5gfe0/RU8+KHlB/6dbXqzOLnoWVskQTu
pPPOG+esPr+6y+rLl1ZG4b4fCkTkhnH3FPu3cwc2xl50fE8kCD8Kk/5nlvg+mAev
UsaXjqB7nwW13fXlzonsmnx7azyYKSmehCEpUwRZodPOc6ka5s2tkLME6Hs/2w/Z
3xkcwFcBkkNd9EwaIm5NFT5HLejMFHObrFXlwDmqeL6Bn0JZqRW7ba8lUMJsTtqQ
CKYkefP97ixZEotDl8e/IJYqso9P0qZcLx6n7ISOcVYbMX3izsMbC8GfsVDoAaaA
8EEUAbTlusF/0XSHHRmWaECvhA0IerAjo4o4C1f9VyE5+Md4ZIKfqdSgOgIAtghi
RzjUyGTic4kLGq7VnvNS2FjiMGvzD73PA5gpy9l0dBDK2o5CuSFG7DluuYajMTBH
mXxINiQqdnr8sG09GlKEh+LyWRZ0dSkvki5UGjTXB4EfuCZIQ5g0G0R5TSiQhlC/
asger7HFBrFbRr2wK7PgTeyvECW7jsg70kXnme7nZDnIP1vjnMpo3DCsOVYHLNLu
tuM5Pnp505I3wUoDCm3BtTkEEmdCui8+Tagi3YDDymC9oVd7OIk8ljBOQ7N3MqRj
WslHgUSfhSute+oibkp77oRC1wJXewlsQcVrpyL6IGaTNkkWBE+67mMb9NjYuWXC
QVZwbtobbA8b1qM/JXIZyEhpjZ3Tr4+aRSfIBE2nc2nwT26/SB8mzTMrA+ZrrHC1
ufos53YbzaZtczMBL7+x6yGtUuPWue8HpuC5TRfYMBN5/Sg7xtmnja0W+xb3xkEd
mG2wklBBg7J7e/Pl0s/dyGXXt9T30x9qa8fdFRPY+SbusSmVVg7Q2RZfHdfY0HjK
QExe0BNLLfaA+IeEh+JDU4YRtfmyGyRACbAClRAdWB8afWLtyE79gh1Yo+UiM+HW
87JjY2neEw8HjP9IFKSi1w5yQMJCJmYvBtW+mwVlFtz86vuh7sFAz29CdZA9+p8f
jfaQkzH6BmxpYLYnQbxPd95pJym3RWJwgY6EXXnU/JA4ry8pJC4xmhJ++vwhW27s
gW1HB5vcjh/xgsuWDdvAlbnJ486vhPmYfp94a/Ukj8sBHWzoHFWMaWdlgrgzEPJX
V89BwC7UE90Ot1wjaSjWtBQ0trhMMzmdl4pZUwMSi0/ZvR3n81Uhg/YgG0jDgjsk
oX5MPb+1U8wZzA7eSruxgq46e7IIbacJ6tOHPXeIXu20GgaHBzrTDTV89DA10gKt
kBf3BQXe46PRlmM5n9nm+cL35eGTxwhGVkD6Rh2AFs6ATYbeF3MCs7aRRXgqH/uj
rbyFfPtj12Qunatk4WBQbokLthaKJtILg6vDqpY8fZ6rkeLhLV+tDeyqsfHVIB3z
TSVpUVqHDPBVWmOR7TWGutf4l+rHdg9dkMsU0KFF0UsCRqARgMtRmD7NcjUTlv0X
paSP2bn5ooCnx/+aC4EZb+Tf0O3270ycebnm4K9T4yes4JuymsFGf/edTFaMsoyV
AkWdK/1yoYVeboEQOKr8G5TM3Qi7dWPzDrH4p/+65CBqgzSOUJBZ677DCjDTH2dk
ePByRhA6KRKwABsmLMz6/R0yRT3MFAVt3NUcsZ6Y7ZWGbZr9cJEyJ+P3/0xjiBKY
oKJknyhoz7e8N5yu/xF3ICYeSMvPRlkNUuy62TvkycOc6lJ1FDuJu0sejGFeOpla
Apxb8d8OGnkfnW1nP3HcwKH41eiDNnyaO0wCxY36bTZPRaUmRlA82TOnIcjVfdLT
oh16w7PyDDLZHRQwPLHS8WF6lg4CO+b/jOGwqfV1fTPSonK9nAPH9LYas4xNfPZn
foleQIT1s8dYFHBcM748YICh4HQHx3R7ZfnZbpSifwtw/LULZiK/kegfp8OgxSHO
UUMvV4TL7eEhNu3fS7jdP2NDehdsbylUc2xhUmNgRkBE1hOHdtCBu9Tgsz8jLy+9
TBfCEZo99uiVqFCYEQmM2HOoiWSuXALkCnHSjTVXuXnIz99MojvC4vFUhKU8N6VW
4p/ENWgVj4WceUqM4pEZaV/bDNqW1IRhGgGud73U0kpAuCxyzfvZd/BV4mJkxJmV
v/uJddMUfkhAsT8EkjdQwPnO/lgcocgMdHDLg2vjssu2eYu+jX6ArsxZnPGBgb4R
IAWnkKOyHfhiyGmx+UP3H43dv/E8O8G1UwAab3AhYNlsZ66yrhl4brT2LYAqNBvC
UTOkxcP87iqomwznFytomDk+ze5PS2IgZnerxou0Cu7+WIV2q9dosPxjsVsfnJKT
2Y6jy8trJExXnYCUj+n9cjTvhbdToIZ5gJ9duMbT87BadPp9i+y5nZL2RwuO3IO+
ZaHO0DQEXvzNWtMo3wGgUKQfCKGNEkWkvPPEU13ifpoUvy2zqXLu3+QSSdC4cRl1
NcWtE3MHtLpllOC3n15Y4RdZwDib4qQYMo+nE6yQ3ApWN1qRm4BlhJB1xQFIV1L0
/6WU42fugYHu8f8VE3uPpAmHxaLZ7q+7KfH4WKVoj1I6CwgGF/XlK+KvJ8iOHzYf
sFWofGa4Tlch1A8bsk/r2E8bHHw0jEobbi07QuOSG1AFL5z2HhTeh1VqX6cs0gGq
bmmDARFXsgSVugv310czalYoczhp9bKbZSeCGJD7fc2bhfJEAPPu8hXChphlwUz6
gMXzPgSwF81D13nY+6CLlYSmRbaGf+kDL4uEG+ehpfL7sgv0bUz/mTut0CeU3hVO
B1PSK/vjDP8Pf6TOdhb5BAYC0tw8MqJX3meHz7iPY28WrG9GaqfquxQ6zuOPCQQn
5Am/pdZDLU1T8EzfRNaujmQY+D+a9pM55SLShnMAFW/Y7whnUwROnp1QMAKEymOY
guAOkkjUUsfyI4KxFv0FxDEraK7QCnC6XfT4jigNrKEdVLakVpZGEuBOtHOSMxka
zX6HIr14SYOfc/Xdx/NTzTFfB9U7Xp5hN+vtzsZICwuiFQ6j19ohYX2cNS9Wot4o
pX0pWAfB/JGVVhKMywGj5OSYQdasdLsyPQHVTzbCLM0ypBsvnLAMIhM3BDbIHldl
5jjHeNLZxBNs628jf+1dpFsWMq1w+Qh66Fs4lQcKU4YCRbw2RqamrZpj62BX3Zaq
jmE/wE2ekVdvlYTA301ovHYLN6ZjELC1cXkwIUGn/CjLaRtjR8lI6ylkn3EGvG2H
Z//HpaS6kPRrvZrSApax95GRj2M9mYlKtlkt1Ixj6BU0zEjE7w175Cl7nK8b0TM4
f4yQCOXijB4XWVxO5bxEE4Yrk/3HTxyzR2xcbhUGDjLWKp+FBzsIxxVm7NXXXvmo
7qPyp7z2lO4bAlhIIZFa7IC/ilEN9WFeB/K/JAt/+ReyoY3j31IIHQx0oUO6yjpa
+i+5jXmFJmICMrL+Lcx61DF5F+ecNMJ9OFZbZ/Px5qLOGiXlLmLUvy1QQKgU06JT
zGhdOZe1XtatpU/4/dswSv/H9hU2sOVRlDZl4I4JHXyZ29b2IgKvvhixnb9BTsiZ
sdUgqFZKeDRjDNyNbUQO9Lzn6XqM3IXJjzjF5hVtSnFL3B3HgnfOV3m4HBh/iP08
GZcBX9qtTkJeYSyGNLwjo74I0e7W78MgK3LiKsIf0kKDConNM0laDjRWq4g8nTKT
v0Hyd3UZ4yJriim1zNMswS2N4/cUZKZxduyFBOxiwobeItIcou7xos946ZkwVMjg
XLAZU3qzyzbM0DVjbetYKIA4ufFziDRPxt8mexAVG2c0+/iFkMZJlko5MSk+I3LA
vczdIdpSEocE5ofQOJsBrfzRBPRT0vX7q9aBVupIE/F6il4X6Ma8OSsoVu/IDfFj
VD3vWOkfnoaz0ZLdlmJmfoHLzqHu+Kc8a1hx/XXbiU+MqHPt5FwLFypg92GsZuKi
t7NtFz45IwnR/z0VxywEMdSm/J/yXP4MX0GSFq/ND94S42xNibisGCFZoX0dVUIr
kHodhAYS6oQbwpsH/9bW+bQQB3YxnsbmEfTs2c2Nr73IVUEots+4Nlocg8Hzo0f2
7bL9D0cDGKiHtC1lUClqq3auLn1NhfHFiA+510s4gQHnT7AXDsj6JBWXkGUiUrYQ
74la1iEghUyIjXWNXbPCaBbePz7XijSj57U6d4S+dqZUgWMNnm4uCpbN0pmF4VUC
8qFLWjlJ2mTk5+qCZL2xO9XjkmAbN3sgkhliZ6YZ1DyVC05r9wMEgkKnKbMwqGwp
Jd986WZMvvTw4x2uJUZ0u2Mh6ncN4oz+EgVDyGNoDVQ+L5RvuUMN2T5qXIFMF/LR
qptt1ajOA9sj7IUv++Z5A5l+lxgKu6Sp6Z08pdRifmwhZPVnT/Nee9z8Nig/fY7H
mMCFD5jVL5RkjxGYZpPzrnWhoNFVl3odi3936W31kaMqBJuofTnd0mDha5KPb6KS
CqOq6mge/KpSGbSGPTm2k2iN6QJt/oOTgWvZUJeaziejBBY1Z9JlfbwbUd2oxnP2
Mss8618++xkARKH2enYPFo3xcNd3NSQ1r8w/74Mhb2gsk4DlB+1ymGYtMdBbzZlq
x1RpQaP5VwLwW8AoJuUGJU5cc4fedhHdJ2rcnYCSp+WYNCAsUlapTh2sgrmgXba0
RjcA5mgP2Meh5490n6NG/CkYJG/x5M2+HpWe5rMl/oZDxawIvWwPPy/k9LWI9+hi
+4KOtXeI0efwOi6ucOoRc0ppB5y/hQe7lwoy8wZxXdjh+9BuYYUHFmHSvv5dED2R
rO9WqNWwLEbaZNgJZV4vMia7P9YwzMFkCQtFPmUdA3GmI4x1tpwOxaEFUC8uqfCh
MxLo/mCst+eIeHqPMEphOXFihLroVDqYHyAf0Ve4dwE1fzb7asbnI4xF15GKhl6Z
HyMUEVxV65NM1GFutHFelzSWb7KHTHP/SS8CBQhqqr4gbmpzNKHCAvz6r1UmHKvA
UtyplMynp6I5exYUAxDa8NBl6aA/Yp+vCZ0HwOela26PjaEUulGTfm6T/pOw+hmq
G+qE2iquyhcEFqyLqicFRFe7wYmtY55cr1toFgPZ9esBcoUA9UexGOVCVsMqoYwD
xxPdHEQQcr5AIHB4P01JsrDXc1m9MgI43O3XIs3LMv1RRY4T94D22dI1WZvGmXfe
lpanTX3jkXXgXy4aS2wGUiiCHsNrGBj0SPZyfHzEueX2+pSRb2UmLOHRP0rPJ2cZ
02ZaXUSVPvTJH1m8euzRzKDdn5hsIzyhhGO1kWOuYESXWpdERHLpT2rq0yKLPjCM
AYy4Sobmw7FpASZOMh5HQPiq0gV62RBFHIWh7nYAzeaMcBBe6oYI67BmPbqfsUi4
gdW7F1GDiYnPYnEaozTO45OdJpFHIYXaniUlBusc9M57aDK31X/RqNICZDJ6YcG5
kJKFYQlsmcem3BHowLy4pL1mNdEQmdmYVp1PUSeHDbKQ30DuXpTFnyUI9OFWZ3ES
NO8b0YJ29zfSkbQ8GL7Fu2VyV9pKFaeOQhSofGyD2NfJFki5kQkC1l4em91Z5TAd
WPBAKV5+VBMA8oeTrnkPAij0SH0MI5O0iBs5lHhZrFzNjS31emGKKt/yhWAKPLOe
mkoPobsgl6OwnCleQ1BjSH70s7aPW9bUMWyxxUH5DtBKgoF60DzBTvCTL2/2fBzU
ycUECQc3RvhjPEI1O3im6YFj5ovb0k1I/AFg/jDKeAoFDSkx7xmLQ89Uvn7gU25d
aUJyv0CLnQFEKFdISnqJuF9Y86XOxNUveBgGijQpSwOijPLRjGUFZeIhWhEiqNM8
COTXb90bsR0leUfkXebmFxzBco7MUPmNmg4PUdt38Sades41BwzW5X1CGcKN/jN/
/+ioL54MgAkR7iP0xxhqAx72JSJ+epSM3+oLmvlxOPCG1PvJH0Cx4iCehdYNJaGB
AZc0Yjnd+NNQAhCDFEV8PLxcg1jpZid6nzEfIZrF7uxQFOC913m+Fp4tgu3qwyi3
eV7JdZE0diyJIbO/xQpz3g3uPHf39wIn3esm4JJj3zRl9pvLjrQBfFXSaiH2bvcE
PhHFBh7H0gs4N6Wfm9hwAhuT8MD9WOjI+TdcLSkXpKC8aQolTs4GwXjkO3RHVNLw
6seDgqNr5HRBN2zZT3x/nOjDtqtcGPw9NZxbROk4hm0DG+BAVulaNFxRe7MlA1PG
gwaXBRQXRZHWFjIDYFWWtR4ON623h31TryOR7xAgrnzsuTs1sTFXQSB2o9vO5+c/
A+aZ6UYCN44d6cSR6Tcx0cG5K94wVy+VFVPWHQAlBjiRg1XeFgpA4aLtIx3cO4xc
nBxe3vUSlLMQ2Ojt5SXwUidY5iOlAaGum1ftosnyX5lczThCVApU3VYKeLC2KA6+
disGAOAwz0S15VjA4HOn7rBNaflT1lA9TcZtUerUy+xn9qDZWDkYZ+XZT7P+Z7dr
Kn06wFx9Y8VKJj7W50OqoQgAozPYh79pp3nlf1nt9beGCzlQEKC06mMQ3fOjVNUs
ziUttFuUrmC60+7j+bv2YTuM1yHO75X0hJIZKr5dql1EbjpTDbzsGselGB72KRcZ
E5lp1AYz2OHpknMPo2PWudzi1wbzvTcY7mbRRDlEcfbVbSIew82C2ORzc63sAOzc
yBYiHv4bkbbdLsN5EhF4z7GFWuHiI7ffuJvQOTQk/hlvlmLaU/gOwEPMPZLacFxB
SrI4ALJkGXtlqtM70n8fABbOteYPJGI2sQkcnN+QXtSfQBtIXx5GoKHCPqJfOR/f
PUSJz0kCl0DladGuZkfw67B50NUrdWDVVvrMlFUY+3Z66JuxzL1CtNVIpxwakYZ2
ckBewiHvPQC1/jb1QigtVb/cSRAdBCJGWP9MK/mLtNI6MRrclokm3hOQulbRtgc2
97Ify6JsldPT7L7N+VR8IXGkd6PJWtwBtbh7+gutZeQLDC8ZhdgVoTDd2Aez9L3A
G///b2EAFjFO/xnsD/60xeEqGu8r7q4kW3hLDS5zQtGPNsTbjP3utfnWkLqJU1ql
IQfLiR66YBUytdSsvxtCzVdClli1aOmOpxRBK1fgVy6SUo4bHvkRHtLyIu/wzx6b
nx2Cpe6uf77FfxKi4jUc2jKdSXYwn+cmOMwIGO5DeG8/A1T4JFPElUhguPaRtRQN
jcaWGNo0t34yT4Xdxsb4MImd42UDsQeyApNctjKy0R/39g0x4Ouu2UUlKLyL3Ibz
1HzNTNnz/mOIqEJWtR0TE9cQ3Ac2n94WtMfuTwxRnkeVLJgnbpbBq3N6qGcyL4v8
z1NRWU5Um6yC6KKvH7eFwSJ6nvlcOvGIuc3km5ZOUmdmxlwsWpRufno34Siz7B1s
u1B6nzSRcGmse1kvDP1lwefIODNJrCMb+RUkGEfxKkG5dD9Mj5hSMwtIyvlcoah9
t/YEzxI+f5HzXaGYsXJI8nuxRIqOKGgFOaSwo/kTXj15v4ZTKnPRqlmR4AEbzMdt
uQ5UgGtz6B4U/Q6ma5UCwf0JkyQuwoMrNvd1R3j9BAEuC1czSLnmvU066RQtx9eV
E43kKr3jslms5Ua9w66rz8opRprjRUW6UkKiT/4Lf1Oe92Dxd0G8imnHR4qy2+to
LFNDpgBbxgOVSQ72zL6PQuMqc0IB8lf1BssW3OFuW+rzTm6ik/2uwvLP2jZuAYpN
SlaJLX7TAI/YmHoX53qKF6aR5x2wNjYO2VAntOMBjyA7Ww0JXbHZxBKFFV6XQkbg
yDb2eLKEDqsgi9eqs0PRpCMDyLO2cut/UnGLM7Pr9Mf2EvS0CZ3u84ZpJ0KNqF/W
XMfe0aamTWXSRDJ5w+3cy4QqJj7DVZ9xJ0piUmGu2lvPYLtg9o3eq3BWHhLWrJmn
KzWPVh23ng8RP/jCZzoDALE4f3aufjJkEEwyOhkrNefIkkkNBnEJLvWuIfZe93LC
AL7CwKH7HQaNy29lfSfG2BVkEAi7lfYlnYQIfyyH5gBiCFh4AsoNYwh0nnPvjkaY
CAwtCRw0NCQZ8eEGSQjNO6kzW9kPfR5j42mrQ4imf4ZYXVN9FLjytGfi0lCjSO/7
NUjhIxU7ItQwe7a/T6ccUgBKI6Dvs/12+J9w7q3ugHE+WcWNwGwGYP+T9cKDG/ni
nHGgBi+UzG4+iiyBvNTDDuleFFYGjU4S18TivF8kMHdMq5oNmaZZk4cbukoECk5s
hkTHX5G/2QZtikEc/TY+d5tB4ZX4MrAXpyDDUWHpjLdSo/riblp/jx1UZjh2jHOY
N2UPgyPSEMD9fUumY7Oqj4jIM/GKeISGM7lODE5yMsrJGFslW07XNKFj8ziJ9uXy
GRhehPYr4mc4XpJE5uv0HjCEm2H5rBhWC60W0rM6jJmUzoozqQ1o9wX6qxvwM2ex
YQcmtkxeAIzCMbmbv3LBTdWoQ98d9ZjLHyuwLjujQLKlSkuYYP0rXSiuUTeiTTwI
AP9igNk7x6OTgUjIVGyGN+FBl1msJsG0WDLJW9PdMxUoh5W6z1hjNaHYWZiBpein
UFuEGO7Bu0WQhu78Jvy1jO5c7ZtkC68VY1PwOnUoXZE0XlBojAtjiuDQZ/WavviM
b+NuTo0VtqhSH8xMgdoHeeBRv8g3YCfgJmC/ufmKI5Fyk/4xzDKWaJVc6c9Yywji
QVHNa48IOw3Blcyo6yfuy8sVFT1I1jGkugZEOBU6Ju3kww4AcrLIEr+oOvpoPl2I
o3uHL3GJ20Zrg9scwoq6/pWfMnHhiKLru5Mdc2VhYeB4VXcUd/62cJBgpIzd5yvU
iyPxpnhCYvAlAKTQ1gNZZJlb08UOSAekhGenF9Q2NEyi78ctVD/Hnuirq1rcmsq8
8ti9yCGglE9ZFV/dyAPfdIpbyNSWYToosxukhyIzOjg/ddZW2ECBtaxwcDd8vR/4
bv8S1ieYOz9UMJr4PnSCirlfvHUeeMjl9BpvNfmzx/6Fy7F2viHr+R0gI3bZS0vn
10w9cHupFOKZEb5yS+WLMp6elnM7lvDnW2a4WsJcXwUFfIdMe9n0tFfgYuj13ygz
a//IVqGsR6a4Z866AnC4EDW+SNYxy5jNjaTLlrUSrtldywVSHhXJD0QcJ+hO92a/
z4UiLeRBld/bL0p+z7Oxi6QZW7mqSNe3fxOizWS8PeafSDLCwdH3fc/98hzBBhoa
O7nf/TaIodr3+rV+kuRT6x9nYiSmRUry9YxK2IL3UdUC63RzoHs6/m1OSEh4Ov2E
smXf+oJQU7uA79KExPI5Le+bHHAajwb/a8+DiZGAB7r/kFEcD5SnUTzoTrUEkKoQ
izBYoEC26/BUIsuIQbYg1a5MmWeX5E47NqNszsSut+Fpsf5DyPbmBzA7uGyOwskW
T8oWh1vTrL2beX8nRBFuUXWvqXqhsDyOxj6vEW3lsut38ptjqiY7JdIdMW8MjkAc
yRL0KLYb/bwlyyiHn7BqRXT2HtR5lp7VqQAqaa8u2MlEuTB3HtcY016aadnlwMDy
NIjrbxCLatEYDwidFlPTRNKZGKswrwPNAfq0YEc/xVgPK0F1uPXCIzram1lReMdq
kRQcOOBP8SgDAw+xNvup6B33gkHRxmO2mjUnSgug9mwBRuarvhpMPWumBwKyG0zg
Oiku7iN6ysBbPtTxcl1QjnRC7podsfnhFJlia3iocsx8raSiFi2WpKZ9+hI7dYXD
jgB/richDz0RcjxAfDb1XBNSAcnjijv5vTxtidn+37LcSGwJmOv9XALAAr5wWlqW
uR2jbCQd5OBbeJ01AHUuHuH1jOQPBPliHyTncGSXLX6nyiQ3Ayfpf2DC/ebByncQ
gjthj1SIXpr1jxQyh7CBiplkYt2WHkyvfOSNAC6GE3ujzAyl/bHSrMJFGv8CEXyc
4WAftP9bnDh4QPXu8iozZvTHXScyqB10JYz1/2h5xTUtrGnKF/4jprau/GWBFIon
ON48tSRTRmcg7mdYiVRzB98/53zKqADYcxT7KQR3uYApz7CxM1GVEqkyd35k+VAM
6xzg8FlUWKkLkwTAdxw8UZdwTNrXavki/SOTm4JG5p9F7WnJnB9YzRL03CR3Rtqm
QYezokkzRvGObrE70SOrpF9ovdDmG1HdymxsEMmsOwSq/hofZnAfsosX50ao+Wve
CUuDl1MWs4jDA8SJvhxjPzLEW29MyNt+15L/7gNkv74tRvCyXVNy5M9NzSpyWf0z
sr1IoUs2E2G3f52+YSF8PdYGEEzOe0AILw3b09fruOzuvJRcRq4mu88XBOf9Kkle
ipbGQTe2r+bcq2/JaX5o+tB+6kaStuRG5A6hWZBEzpgP1ajEnRqq1Dz9os8xywyn
tD8EPoCbPmRYukp8aKB237PFfUZzEdqJKwcKKHTYus9T+bjJB4wOslJsBfSqFO0U
f2V7PYVUfak0H2Stm/kAM/NHIPD8nBtTFjzmUtZ/VoaTn/xUZgl+CZGODvqWUTAn
qfoN3M8jJkDFD1K3CQesIOGZul7F69OfJ6B0tnTTpoVzj1nHOB69nglaBqVsm8tI
KeSkMeaTmGT0XippELVAyFyyjusrmUoavHnQFdJq+9+qr27oSXFDo+kMS5ihczKX
0VgCPAnCCYqjCi2+WlTjQDAu2M4CtGS0NgN/n7gKd3Bv1totGW3juFMhj6xjx0Z1
q1FUxRbJ+JQh/ecvhLYxpa5ocMYZXE5X8zAP3wuzWhD6Ll2B2MNP5ErLQn9c1GFH
qo7r3pO4Xi3xnGMjHCiUnnL+cz2Kon+0iHBzFmMug0Dp3AtGGTwfnPD+FTcNUTuQ
eubVXbgB3ElRyb0FkqyEecJwMyR6BMCYuW87KAst45t+nT0wCWUABPZsh14EU4W7
5TEV7mp3QP5EfgLq6cbW0G0zH0xZ+6r9BZVcrnW70Njp+mvURwE79mm3SZxZAjLn
PO6JV9n8fcXN+UUoXYO7CyatEWGK9nUMRhGtI7OEXQtIa2pi8tvDdKq5jR7xpcyI
TaURqg3Vfkea9XimcwFfp/ZcnMl/VwZ4bndqBowI2kkhOouruAJzKO0qyMmS4iYJ
WhQjwc9Af1SHPeTcDNogSwVOe+IFy7htU04jZp66ucqBC6GoJ1dioKwSdImrysIj
73uQW1ueFBZ34969bPikcmFouLbyyFFos+KNAwR6D8nCiMv99B9N9oP8c/k6hzz8
s+SsKIXpoPV9ZehvEEEo0nzOedAR222CDij3+p/kz3cp/YqTc3RpAL7wd0+EjDA/
VwCmYiA2WuYxcMv45fOf+cfZrkApO2Lirj7paHsZpVjk8QpnOjS1DsMjjRwuxIiv
Gy1V8Cs2vgjpqORjq1HyR8Tw0YDGvgqDe8sRx/bZIfA8fpIeQis0LcmAlY1SJFkJ
/XOHL8rP5YA469T5hakZ2AO50vXfqTeT39eGCLTrJQYZ8ph1wGwptakDNaGVvzrr
iVDPrPZjdikygI+ybj5J2ZuXEypRAEyNlfO8I1WGIbJWmiblB+SlHoMTKfvl8QGE
EvGMIcstdg4LfaVrNEDkmM3r5hFLzPFpFrNlV0pLYatUZHdFVqSvrmwQUNWZGY8e
FcIK2WdXSAQq3gsiswa1iImoTi4pMzlTuKzkaXhdhlLFAZWk57REPy/wv6XSV80a
9zJsDhrZUGWDRDvbs1W3cPBAd6MqPlfo0WV836O3vpE0MbJkCb/0hhtQFAudMkXd
TIln5UY0dUskS8Tj872/FN+mmuNg9BNZFxes9VFc7cjyvzn1W44xh+bJQtvc3bhx
whymW8rGN1Ks/FHgtA1QMyHxZFHmqNxoLd+s7UkK7O4TGYBdN6qJBDKHCao2QsmP
kOBgfqjR57bTiJC2NKn/WUEjNdUSPGAzRy8wsD06OtFO9E20WYXWpz/PCWaQ622C
sGxtbkWpQkMOq6tmayBlZa1x5uh2lskACIoYcQhRKMa96DcDg0gqbYhBNFykJl90
3pQ3kRZxaGhzcg7bWzTJQSPTjj3hlbxqTtf0VPL5paulfztTpK1I1R34GsHioKFc
BHvR++91IZa8qGjlCPKflcsnBiToTdT4Tk+TTrSQDdR9Vxwe9AheDVQF6bQlCpYN
H7sOYreXoF/r6MpPv7J7KDja4gC3eJma+OH7bQd549Y851Je09JwjK0faGq6gC9q
Oqb7FNcz9C8N/ka9l4Om2go3LZafQ/QyCXoiSrMF/cu9Ide0inRdbZsfdQ0c1kcX
fuzMBtKoD67MgJuBHnOzVNNWPAWjEhHgT+ym9sWAL/myRhvqiQrreJSLQFSL0odf
VMERAhSzzYtUYKr3jdz6x7rQDU1IcOSd3ROEfrz9DfQJGC0QSWl3esHSZoO9nq7w
5q4K1G2RGiTuJ3nKBaIfaYOpDWw9GmrncpVro5Bl6Ex+GGZYafgMC+WjLcz4b1d9
D68esXNd0xaurYI5NbmYacLm7pXPDlqAsC4EYcRbhgOXJkNb2iwNLA0/P/dneGXV
/oJxmSmIr3mq3VcSZK1v8SOWu0JpK2cQ+wY9gAx7ImcDsZPv6KIgHY8L+Czph31G
0yk6/2WLuqQifYsgYsZy+RGSRvOiDj/3vVnhopEQ8Db5ts2ss1BHA6famae/VFff
uSuyFmOGAvhpINrhTI/zp78IZ53yubDLO0FFoYTsNRZPlxFAQ/Azh2ZkFVBf28G2
mwVoZ/Cf1NhfhMxHTI3ODayDqDcy5yKXRenJBIBNigO/l9he44UU2I3Cv9JmyAKq
GJmZL2Tv0oQvRtX/v72DljO4XU6PcKX3aT5lfApeihkCrXEIOgjC03KmJYmLZ1wW
kCAbEb5/7kvJPZdiH8YM6UiHQfdTQc8WwrQwofVr2G0PoFKWgPNedkFR5BckyUZ2
OyHzTFsV6J8Kj6FjG/1/DE3TvltuYYm046+1IeZgmj9plQej7mHuXGLp9qIXPfrf
4pINWedlU4cXXSqhoEcwwk1vT4+L4rJfSoD2Yxl82bIjhpk1fRta3xN4al2YkXYO
hzeD6sFubWFn2QtPYqXDzj5pS9DGeJT254haZYV43e7zvYqaEzFyFoFnqWmNSgTl
KzAxJdhE2PBhBLHlEOxKUo4W0HcAa6DQEecUVXUYcblDTOX4tprpepyIDuK+A4Hb
UZIHvXeTh1w69hr7uSmi3lnIUgICcPPr8P34ocPEk92AzdQC0L/SiWa2z+nczyrz
Shqvn7ZuOwjClie9NP9FxW4Octhf9xR+HMwRmTvNp4UNKvgpzYLNGfG6nRKLgfcq
uvzUvgPBfRoKMX/TkRGjPdf1AOr0oxWaIn7xCfZ5V4ZBOdymUf0YS8GXsdipgL9T
ejljfrkKG5bpKixDEMExiFd+C8Qw2Ca46bydlpjQulaFFHW8X59L2qpUtKPSsqpy
oG2zeV7uiRyhxt8AAxMSbkooqW9lt2hqGFlTh0H9Hd8Q5txqxzHzvPLxJOK5sWXU
De6n6mR6GUXSCE4JOBA0bqnFe/oaQiQ8JBH+1EtGMAy4GoDSqk9ooKnBTe3Jq5t8
RsbZ/g2XuLBAD50Qsgwr7PdmvEiE2sz1uuVya36EGBUaH5q6dFLZ0TlpwkMqlOro
qTLa6/xbMe0InBZNOkBqUx9QAIOFcbiX5V7gVM04LTudrOtdKuguu9LqyO4sA6Ui
D7EzxMwbb7egmDnflkHasawXBypuIjbo7JeY1Kz6PdnxddmI92aXHV4ZjMI456wc
3XpKxxNLTgUMA4ytH32Xw/86QVfz5Z0lTFejxf+sebCX8e54LXN2W24vJQ9P+4+O
IAT9J7xd/nY+UnNq8qj43nbFp6sb01lNBKAwvg2ngX7J7iXXCfY7Dw0nY3lnJTMG
0b3UFDiZVNSbmybAzGqL6X3HT6Z6xQunSL2LW1/68iaVGqzud6OS3MeMovgrOtK6
cmy+HvwjtlDLI2dUp55P0xnrQE7HSlvzaPulVm93JJRrhpulDCa5XpqSRskvNcAR
8dDPZyeEeYbz4rO1LEZH20mfUfuAWmGE9+3OFKVan/pPgmXtXIZFd3Pzcg/gpIvE
zuMJSFLij5NWgO++e96K2aFwoTcc1S89BRA7yliGmK8gUWdO5UJ+JwKfRjFcIJe0
BxfjDayed2+D1q6iUW2s/jvP2E2hb6rIifUjom6W7zevCo64nHBv2MEUKUqBYWLh
BN0ZN3Mh82h9S0kPDgjpgkBAOyhYxziLIz83KA56mYCeIuF2wqjsIWq5NUP1n4vs
vgj1+HH8M0WforjXvcuum5QXPOAVFd8mQ/mUVFeURVLCY7+4O7hwDp47jdfb1bLP
5qtNRgjP2gbQSvWXD0Y1XCH00Lzs7Nrz8acPaNjj6AQDQaAa8UqW4lxKqTJCNwh3
F9HdSVmE6NuXc55SCEhvMWGRdhYJkj6dSSn9azltwvQSdna6Maksd8YBwHR9eTjo
WT+yU6wfqce3a0KD2S0cL9xM9TIAqHTq8cuWiTdOETWO9kjoaqY2eVurwCWcPTn7
JeCPmqWnQqXBuHY0zgCpnTo8LxTjut78vTpEXMRjVQm+6RceOvSO8jqhWGHmusxs
v8EN0JrtI/a4iBAMLS2OGMRs2iwcZPHArBP4WWlhDbwkWlSCYSxyBlZQ+1FsCdLU
OA9qdliZkGoEdt57w+D+3lIK16veZTVeI4RgU0yy05+CzoB2v0+kJfKUae3L7QHt
21Q+GY34RVjxNxuDqISVh1LKzJ+g7oPdfD3D6zKm+jgvuRxbVfdU+CuNTk6sZ9ZH
CP6JOediK8pocfu4RgPXbrOSWsGOmOiZeEsluxB2R4BiDscOHFAPf357ijJ4Fmo2
mFC+TA8Y9DjQTTXH24K5P+v3DDaL10weg+RcfXvfmtuvWvXhKo+9rI5iFUzsmRlu
LBrfxQJAyhAcPh4F2P+86z/btqe6quWDO8hyGaxZXLY8O779SHtKIauMh7VX0ngD
09K8bpR5ocU2MX1Unxv0ErcdHKbRkGxlv24+WKu2WZ19uUol4r6inbQYDOsjdDX3
2ETZlfXxdU6KfuojjQTrNI0Cn1XVvQtsQj70QZ1XY4Yu6fxqYfu48IPticAgopG6
VKgX4egbYLLZm3mrVpjugECGP6lFMPT/R4uic+L6EVB4Rg6rM8ApoLlIj3OtIpDp
QNFmZJdSGp+uT8iUjTJB+MlfIQh6Os4LlxVhQVmZ5XctFFfWhxb5LWseZkbsBLrX
726Ru4Fm7q/x4wa2unAmIDovxNOjUf49La8lIyobk2ohDZNioikKFJcFr+haOKTT
m1h7jBUugDZ9tZ7/qD2Vqg/UaScQXCZHOi9Q6K0P3bs6PxlciNWwqmyuEMKFTWkQ
LOHLovmXpqoCS4QJM2reAVlNwyoyZxES85rPZH4bKgjzsad1j4HEWBU+xLqpgfOp
4FJTiUDYGSSNjLZGtq97aTrxKBjDN3xlUBOTOoSS/Q7adZYAwGmz3N4pRNu/nYe7
QBTabuMUOzGEqVUD9vLs9P1LOeGWPwU34KoDtIlornGVjIxsUOpvjZ8OILMbaZn+
P/yqJfsCEVg7sD/UOxMq+GhClDX4UeK8AOefv1YluzuA07jhh+SLNiEXCF1LHoI+
4Nc0e7xV5Jh9/7d6iUOEb3QpF60dhObn3GA9CzWimn4uw4J2MzqhsjgPJ807bmv+
GkNgZwLCMthAAA3ipf+33E3JRngII+aDarA53MmU3SgYFcMCZGL9V8qFsPmAhb6W
tgvh9uxGkVPLy6JP1h63r6vbg+rCz5f1RmRNFkipZA8KQS1ORIFrl2tTzjK32Pjc
9xkKAKtjjjZGLHVLy7ofUPKmrtkdCj+/E2lTLSTqBlt3tBrio60+8c38k14GGO/j
WFsNO+K3EIp2nV5iU5bolPaiBX5WIMW6sBU/7KFwWf8JcK7ww9KuUR5e4LaJomp0
8rzsiljN6CnabUk4dNJWA+K2fgL88A0Tcc43v+lPeSevMWWMzRcIK0tCf7EC+5T7
5/ZfunE9/Kyn57SfJ2cmLgIjDbQuCNj9u9L0uKEW7/idRJSFXWu0YUqeKz4olPHM
85IC6EEHM769nBSzk9kX7N+EJjBU5zH/30X0wvOp6lwBIdkI591TI1jUDWAGnQrZ
nD34YAnawEulPNl7haSxUxBMLPPaJ5wD+Kyst8DHfO+G0P6p74uqPx9rGvsMt1BV
zMCz2CPHaEjiERXSQlMdnv+xVnuGvex7HUQ1jMHMo3nZdzxVAqEvxcwAkmuB9pxw
GJnJrvliGXw2tWub0+3l7wvuIgQhxQgEwrnyksf6G7+utZdK4JgV+DsySAuSMByH
PCQoxTrGXOwXbj33abKY7T4ZhOWDwaVFlN56fLTXo/4zHwNVkrzC32+FBlrjguBe
yulF5J1tf72oVWc0EcY2zNVFX6CXk5IfvRjuSgz2sOXiyxDq3Cy1u57GqpTS2cVW
Skg7ENGhYL0VB8Du5C9N3+T3+librkMG+piRqOiyuRo8WHpGi+Rn54rtSTty9BS2
9sc+ELW7DqMhXNf/RFZVBMhrDPSriKUQV2gl/zMPBzIZyL2dWb9o0GxRsVEiJh3+
vmfPthDcBT95FHXdIf1aMg4LWQ0+vyVgAAXBksisRo2bJqSb4gd97z18DAzM5bsm
qNHx6nxTFzl1debxcs+pM6LInmpQTkzdfbt3vM0OThECqkvONE3vTZdwoq7yW4zM
OKQFVRfVtha+GTTAsUnFrsFvz8XGBHsv+rQgUa7B+TBlcsW1iCN8XGVJ25WFJ9l+
lzeaR1wrdiqsvOoFoFwMM6HDUjkLlCrVVokUumzWC2pUrHYA/bPfbijBQrLLkwJO
4R3B2u+sEJWNE1+MqZzIHlRnsFFuQhhOVRv5fYpXx3UICWxcSgwpvzhgjkE0lyZO
Hk8X9K9xjp3Q4Rp3bchEkGXqBcEw8w5t1PP4jVOoqZqsIfyOj1BRZQ4t1kr9JBFa
UmzHMWxJOhWKHrHiv/mobusFMb9bq7WT6xxIDpRu1MS6283mwbfWZyq/8Jnt4oLL
z09x8ZXYo4UwLwBlOQuFxOWOqE1Zq+OhbSGEekTJIpcAwMhyufubnKSkSkGWDIRz
W7KZJ5XfWacLe+7YQYLGlyRfYXjO4730Kc/YhtLeRclG5Qg2hqaWnBBru7/r1xw2
El4By/xjQ+kSxSZVy0gJfOrePYvsduHC/Ovieu5r/jpSV/MGaARGMgZFODkajwJM
IV23scjM3DT82P1BPb2GzNz3S7VtCc9jXEtj824IRaDgKxdm2EID/Lgj6XThT1x+
ceFuN0gzrc7HOo+9rVD3puuSsv1XzNuM9aLmh1wQOpFbmm1QOsRW+JipqDg8Fu5N
BaPXR+Woqf2Sh6pjLnjUyc44493WzMgtPEZibo/h9KpoqrJ1A3nsrF69+mAZ1xzx
84GikKE+7gbWkVbCGJDAxwqccOLh1DagG5QjJ/3wUQW5pBXPIhFwFA6b4Tk2A5x4
ODESnSFjoKi83fdAdcauTFXnI5XgieAezEGtpyGl4gSMdgEjKp+VVM1ie8ysxKcM
lLn6SJc/4jhUc5fKNxIaxHh6HLiwuuHz9SDOiplG0SQ47Xd47azmPnh7afATVUGA
+QSuuW5Gc/ZxZKmG2pakVhu7yS2AnRYN+h7m+bHQlCsTzWWYHTG6muIy9XMeue8L
7dfNUnh2OSv4yf3qe8x8V+FwD22RoCHOM0UOAfKnGqUBgg6gN/w9ji8ZY1ybf2Xz
Tg6N6yaBe99raijCZ951iOikSjuXQg5mT00Eo6M8oVXfNGU215vfXxDQkI+jKrPP
C1MsnQZU4LRwIaJtTSC5f1wNurYMo7eBlbEVk2UyjOhmN1wxqf2ulkuCGWqYlFDZ
B1TDW8RRjhLdEpYuDLFQ8rncgZFL4y5ETAIOe5zhdt2gN3NxA9l0U+iAOAj+YFO7
C9ZnTZaLE1GXIpBegBNEyO3YdNnZ5sVgkqypL7P6hEiK4GI1o+gccXBE+Bor4197
BSclcHxI37vVM89KIShYW1/h8iNbVMwVZn80wDw3Ot7nK0AbiJVs/xNtg7VVm0y6
LHd/CQobhCKqMBdS0LBlT0NLmnFTIMbR+mZgleWYnlEcSDg2arxawjClZXnHd7v3
CC9nJeS+GIGUmJ/M6+rqfZxpOZEHyMcPiZeqoSI0eT/OuC9IHe/pOQW6Wc1OzWcp
zU4t5FYRkmM7tH1J7Wd8QGcB0VPoWMJBaefyTob1jW119I/Qmo0kYmslwpXC0On5
vW1rQN5sWetwwWucCPgjZlxc6qSISwhsdWM/O6e6be5CWKqUJ2jpAKRmx1mZ2LkB
75ZoFMI4iBKk5vf4Xia+3SQ9mhbGbMhb1m3ZAq42EzoX2oGxvNuoLXc6ICnr45xf
nkYlO9kS/sG393Zvd+k8eCWvduEUUVwIo/ITWjbyhGheicMNffuu6Zk3u05FieZD
j/bTvQYdGgqA2Kp147Jik3fK5m8Ne/bHlU9q5m2o9zGoP5XdvECoFtiQRQCfXqrY
1FNiI2wCNmAwLHeYyDIWuKfQk6NQuCY56owHzmNyOjdItqc4m9vYaoQ77OShb43U
xnwsR31Wg6fqXjTr+hqwIhCCNWQAgX9+BnyaghuzpaGGBk1YYjzrPsQP1+P5mb3O
BIYFFNx2u1KIVmnIyE2aZsQLSjdle9asaFOpZsw8CKiJht+5kSqwZEW7jQeh6bJs
8cLTYP4qYRpPj/Swhwp/bdDN+x1ygNvf8Z/Jo5M8X52esdTnnFZwgpKjtQWhpQSz
jWLrD/berp/exUiqqZo4inTf75j/VzK0IoDahygmKjRkrcVgoh2fowVMcjh63roy
8oG2yL9Xq03ZpZEW2L36DaIY30ZRJHr+BWvA7zKq9+q2FMDl+Dp0V4kB5Vsbt1Ba
HF2CqeCD4gIiCiSqxSB4GH8tMobBtwCi93ZPop3Dglm/4bf1uTQqhT5dpa0N+bH9
3xOLjVzHU5GPIVDlqqPTgqQLZP7ZtuaW4wmPEBiw7C8VW4e8PtkS+OEhh7jlUC+z
HsK1bWVTHqbvvXsFGjnIJENbAQ0/UV/kaVC5y6nV19ZXeEHYq3BRjRzqTZ8E6NLQ
6vR/W82gx7/c5YRnvk1oEeuv7VDft8k7pWeLBob4gd48V4p6k+wuoWuCK3klE/Zu
vl3ogYPOXMuGtKI6fKMwpf5lXIfDca7YQW37e1zT0muHuTdfwbgDxVuHaHPoQUgI
GOn58+cOZM5uvsOqDpdxfeIBi+BR6A1o+GlkyHjGpnApnSqAA9XxEeV1aFFIqnfC
ojgmhQ275evKqfkHT4I64hpWrwCa34rv7uAf1LNhjPNjAsnMxO8Vc+l1LnlB2BB+
BnJttw4An101klF7I2jJc43HDEtXio7qALHD9PVsymiKC/LO405BWGD3nLZgwXgj
iw/+dEm8n8PTjP8rkGIAVBpVMS7ZXWHXHP+CszerJj+Sp9up8gz9OFjCwEENQ88Z
EE3r9udDv+q2gAsh92Xe5gt/f8bVgQZVQHq+mUK+CYHtB5guQtt4zwLzsR0WusFi
Zh7MvAp2/nB8cUXN4zjOD6Tw9UsAjoBkZIAF+/6I22/vBRkNtZC4CpWUzC9UIcw9
//DECvjQwdquriRNvFFk7k82UWtrQNjH6OSBfk2zlbPRkfAG3nbCePNotH30HeF2
J9YvlF6C+o0IV0/zjrE2A4q4wNdmPFNn13gGcrCulZlTN0znroo1eOKdwBU4GOzh
BcLRZJRtVJ31J3qIUwD0vvZazQWPs2hI3JNzpVefIkc+MnWwtyhnJ8D5uv0VCP8R
jN+YILuxQd1s8ZN8K0jev+E/SQdsjv6DwM9QpHy659/aFO0oBivMWwzl0rcwocnL
TRQzANsOxiT7TuR3vHuoQBIeKW4UiIiKKJly726Tix7qLsxX7ewnBTq8byETKp9K
uiIV6pdUHY4klXaEA9K9yLuWDl7f97hMpygEIbxsLimAj/WPcHNu9tQhMEy2H/gR
UGXGORP+FlJOizojr4qS1YfJOCUJ3j1cVCAmRIh9wMum3KLbSD2XsA6/82qH0Cz9
KxJUAOT1MuwNjYLKdX/dO9ani26AW2vReDYQmb9/ZWqMlzM2OS0NYx3xxan4vKqT
PJoXxPs6nKvVWCFgk+Ye1syA42IENfzXFET0i/MWKbd4ktaOsp/2+j71jK/23+nZ
uh1qMCVFUpyAyYlCurSq4/yC0tvb8uUrJUwZKm+zlm1ABhy1tjjTdTCJ2yjPYqrq
/duCQHz9YYpHcjrRnCVdKuGJl7lmB2Vo6tSIQFQzSZaBzhrnQeaovKSLHm+LG+V+
t+RoL6Fi58+lelVVQxiCJjhjZc3I4YjwhY3X74FuRVPRyT+1NRDlfhaIExxjYClQ
KLAH74+SRWa6m+vEnf/EiPDHEUwJFiE4HE1V6JHq/XH7T2mjAf4lnZTWu8SbOevT
NCiNRR8mBXdqwk5px0DyNeDpHSWpoZsJne8xKvUuXX9DlU3Ji0XQFuJ1gdxHVjS+
8k3QVKkVjjEYCTmFJMLqTrs6VCwHKhEsBbreTn7qJig3W+VTDQvEOQMUxEwYAAFH
u1VysyHB4WdOt7O5Rl/L+4qUZp4O8nDBh0ZQ2dk4+VlUo0TLjKKLKQLsC78CVcAs
w7qfc71tCzx6FJwqoWRziEijV92/cjMPxO3KnV0YhHWjgivSQu9WCK8ToSy7kbsN
xRJfvGAJkbEfXdrLxauYPgFWDwyYJuxBN44bQAxEC9utwrLdoRX2FxoY7a2XkQ5I
Br3MCWKwQIUCa1Zz2c6FsDfyufDwdmRJuH7UXI0Z/rqTcy74WB29NNhkJz4Oh1KD
tmbaeZeKGFDIh/S6dEg/6xpIuPk+WUuoe18hYRc63BDRui5yzrzoNiz7ZNGEpwAJ
ee67Zo+K7waSyakBUsXFn9y3JjDfuPgRtLZhac0r2TY9dXclhm16Wiimlb5cM5u7
KUGmZYhfEHVIhyxXi4etjGgrQDfzioqBupQOEaz2H6Jsfv9GzQ3Wtp3LYT7jPpPP
2xF+9lB2lciO+nsseEWZTMOqtSrpqg9aupLoUDxy+M5mbc05/wuciCzq+R1P0Io+
l9SMQyDpDZQh0hPn+oucQBKoRqtaGkCtIUVNs0TG6zMpbAWildardxRZfzrPs4Ht
7pv1g7zgG3e3whG5SJsGfOhk5WafqVg20UAiwqDl2AYjcPcih7mnZp4O/Rpde4K2
rcPqTOW/VDSZWbMSeAGppTPUjMbiqeFYZdBHTtugckSh32jW0QDf3ZgVpjUGsmzB
XSptnsKl60/2/ayQl3IXVtMoJdRXBcfhREf7WEklzfyAHvqkY8wjWA8ijafT9fRh
vfaTUx+xBITQK3VwDDstwF+HoxfWddbemOMRNLiVQY6UMD+DdDlwG0mpece95wxa
vnSLVxxt68gyKJdznOjsIrjjTiA2sWxk3PeodrNlKp7hBUWAzQrfu0kf2iVTfVOJ
YLBRrUpmir/vJP9k61wVpWrWiVTzvMTxShpkwpBhIVRjoptarxekKCe2fHQMxhEY
YAGCtC3wmMPrNL/e6NjzKqI8JFRrfOEy2eUtlP+TeZFWLkmv2MACOACqaCTl+Hm6
mgq0OxlBRFLAXMQx6Dy/GTHZCVf0hRJ/LGxlt4gCFuMJBQXyJGrE/WfydB9HmdUr
RuA/HyyBG5PfVzgxtUon3yhQ+//SCdMg/XM/yKgdE99XnO1nQijWoJI6h1nNTurw
G92yalPGNhi9FsyvcDPQrEuopVGPxzKEUvmrFbUmaZNZ/31mnCVuks25mULTcr+5
8PYlkKEbA8dukUfXu2887YWrpyZ8u85Kvaj6rwT5mxRt1fLO70T+591H4SvdQRed
6a3w/oY3Rq+fOAe4UNEKuuUdxGRH/me+FxXdQhg2TRWoHuQwZOXd4ZS2+XXJkFWl
2vjeicB/vxwXWg9WCQ6/TfMGe2hNnPbz8N0cbKz+ij1mxDpNrVkNQ21hkU3YrEdH
aCheDtULa62rW5sR1Ilis/Xc0P+WA0at/TckVbdn7m4mY+ojfKBA3Uv08ZDrGzVl
KIsC8kjn+shLSqxemYAJ4yuroc3oUrkIgsfJBzk34/Kx7k1fMho9NEYg7XKdX+Aa
zofdnR7naJu+d7JLP2bQ1kyIeGHjIqtrkdyei4tgOMptCBAldiFsr6zi335mHLJk
TCw6hXU3jwyRoJVRMsPZQDPG4YZgAQMR6jpsDCKK+wFWx0IEzscTgm08a7E/Eu0L
NaohUar84r1r/R/nHHR/7R+0Q4PIDVJ874ZObrZ0ZDBrhANbkPbT7V9t05Y7OhR+
ZDSCq3C098OdoEjTl0ul8RuqBpZ3Arpp+r8COm11oXx3lU/f1+/F9iZq+905Rw/m
3MuB+S6pY786OauQqDYYP6cw0ERXMlnCDmJJvrLEHnT1bbIjYCbGR4//mbV9QgJr
aHq5kh9EljvGj/bUI/06ELr4NXlbS3nMgOnjJyo/1SEeraRkCpRHnwihvYNen30l
bkp/7ad7wyo7uGKo5yIx+Fg/iZUWbD190xdgFBei1s/lr8j2yLc2a8Em1q2nevZZ
Fy/DC/iTW6PY92KaT6lZoCDUz3SwqcFMam1NdWuQYw3a20ZZfwB3h0ZU3zPO5V2R
8oBlqPRbo2gQFJr6xA6Sug6nqL27FfxhjRotl/KnlMjF0z9otG3j3RYWjW8EFoHC
jhWJDSZQq24/kLn/BjazG7FI86oZD/QEUcypMWSeo9C7AZlZiSYV+RYRlJU3Mi3H
pJYxcTMY/IHIkWZmF2DOyBofNm0Xv/bkf0fUfYzxs1DNw/u3FiQrtBhA1eaAAhKM
LBZaXD7dFB4MKmp795rlYzFIaiG1X9gQTo/N0Q8COP2Dp/NOZ8ylxYpktiMaKZ5C
sZ2mYd0DcmgfvsQAGz4xKEawwo820ZTstVjcUaebrUvuoSNdu7YqFXym08Hm8KNj
NFQaugvkegwdB4qRS0XGM+rpdD4B2FUrji3jMMBDD3B3dldeOkPoeEY0ueSg+RH7
4eJyK6lB+8n6tH29ZxwXXvqIjaXEb8oJuMKV82IqNVBcGzAw19UABCluwLY3ySv3
j9JDG4XLlw1Iqo6UDgg+lgiTc65AdOnJacMx9goXkNAbY8zNXh6/oujv51Y9CRmA
JbIjtm8x+UR8TSsOI9o3o0bgE38fw5wq1a8RC+ScCMGGYNeA4owHqkl/SWBE2zqt
MsPvQJaUMhW0Ck3RHcZ89NBwFkCZvHxeNpQSKcUF/zT1+gvfiXer/lUpCVd6uYUy
3qZqRFUFy97pq2afp4cfI/MMKzFQyAqBzjrT0lAUdGo3RZjudmuUOBopTOmb7SS8
XZJH9ubxh3dX53Nvr7KnUgzj7RuXYmSpD0vHkCfK12jjfv/8IddL/ew/SyQlGn9z
xvqc3NH7RCy22Rd+7Fv5OK7rHxJlL4KAqpKn67Zq7aSUHBVXOchsNWSfFUiom4NZ
C8GG8U/lsadM4GLOAUmBDTqvo+jDCi9eczcub7GIQCUbPoTtVtGlbaeM7rUe2emK
MUD17p1Mto7siVB/UheKuH4pHKkqtI9953Un7mXEQzS1IRwnj6m3l1cl5gT2t0+x
pyoLzB1q73Kw5/1XpGgO0r6lFmboj1nbith+NIVwGUZJe+L7ZIbcU1CwUuOQV+0O
lBXfXgbWhaZO03M/elST0+gDYD8mJ235QyzGs3vF9mTviNq+Nmic9hA2N0gtIHgI
CimJnFLdlF3cAKAOO/o/mdpAUdE8zc4fMubR7TFQtW6v83RRYDzDRsy4KSfnLT3S
142yBVJShc4NjcJ2jJDzA4RdjFpIiWHjSVgVH1e/bxLRZdnHpth5a0gsTIRqIvfr
xNmIlAFRSrUNnYkXuzVqSXAj1VIytlPFvA2ubEQmpGH05Dd4lNRzpiC7R559wydY
C/s5Pf7tgoWLWRQxwHfJwRRtKu08fKhA2Dk2tX5kYZ5tELsBcbeOOy5BNVBsppXg
fBjLGnOC+7rdsgdncrwEM8Sji1+mLrSOzvO1vsnAMLAgWmOG9I37Y9l4lVVwIUyX
qeFgaJuTmvGGpRKReSKYdFOXQwRLiW6XpszRpmQJiXaeF4rEGFOTAaralbk+nEJy
9AhDzupMeHn1R+/36qdCwVyM0VnfZwdwQ90rMCYhPFs76cTtTSYb8i9xasB7C7pp
uUxSYPUZElF3Gm6tY81XlYTTrslKGTigKp038jI1AIL5n4vwpEmhi3jptUza5Cpm
xCWaqbxeWn+vfyOa3kOBV2IwCmbTGt6GEd0XioQwCyeoW5N/ARBQwqlvMiAT/6nv
T51ZetmhdMRmqHlqtyw7E+KKFQKMq6wUGHymXl25krcRusoz/NL2pAgw581f8XvU
rwJQEz8ml0gpTbpxs1Zj3t6eBoDr378xgxAg/w2OnUP5FTreRUdyn//xFXx189yJ
Ti8tcH8qhwM8qdOefGZzhLdN18wrRofDd879OKNPbJLpXzi65RqEVVHT0rKHX5X+
tmsIV+RA7nlvwXumjNobPVvLzd86dRWjKIxzeblu6Eagp3S10229sCw7coEOA9oC
uvxslLl0dlhTooexQhWHNr016UNAHhHpQXJKtnzVk84MCeKEN6cAxaEeD+cpUQ/a
vqp11bzFcwpT020fPPcERReLeEMZY+ONO+7BoY6/IffHsme07tRNIuGRigjXW93R
J/2eceQRX5ZzLs7tdisQBvKLE+snXqh04WkFtE4bchAG6td8HrJwuUWaKkx2FgEF
rxR+ZPRVKcx5DKwwUHwViq7dkgdX0dIHvv1DLQrgPRbpMfLA1Z1QxCDwqKZ5ajEF
vjkGHi2uXWFmatqO4SA2A8g35gcAS2SAtupLMqV5kDA3KZnQG6LePBcqv0wWntNu
wlPHNA5bbHpbxjbnvktwqrtlsG88O3w01twP5GoDDfwoaGAJFXsMvcBU+RIYm8Lt
IwIzC8vtcSqjEBNxx9EZGEVyj9iGZmdgj/ev/Zm1IrYOaC91xNf4m/IlLTAMrY16
2lGNWReL1IIYirVHI3ionAaq1TPMTtGRPAEdwXk9WIfQwNVkjhoVbkUPgc6UQtak
49lGP6F/zpcloKmEvVFlMEGPuqDDW8wyB6M1jZ7xVeraRXqnaYJSTox3EbFjjqoF
Q7RYK/pzfTHatKMUHCB+LbwhWiA8+utb0Dox4/xYDJYvGWPgMwNx4NNQRTGTzXZr
Jox9WlcbSI3lo9rkHAS6bK/OBwnp/IWHMSXXetYhU5FBeEMwusV+qoFpGqG1ehHn
dxPCuH7cdeDVRrFbQM7HL7iYTbUb2z5fGVg6tnbRzDlt5Yckdy/1KG2CLBlRCSIG
S4LCxmsXJcYw3A2OgNgoaL8kxeVEwyo2bVomaQyO2Suc8Wht59DwpLgZNf+LxA+0
s6HgLKB8BdBI1Yff789SCb7tLm4B1O+J/yVnE0DKcoCfmF+BbQIeNRurOr/LCgL8
ZNTb8+dM09O0ta3Q7ojWMIgv1kBg+ZDlCRhDCzc4+4FSVYQEvhd8i5F/xeLvL1yc
ip6mpUnXJ5xXrbLlzCUnqAdIb4MVu3LWz/QT9ay9/j/d9aUOYSPZrzPQ1zio9rN6
Q8J+hxge7281NVkmSEtxUPzXzLWk5+tZnwXgGSawov67tO2juJoAFvww7pSmhDjQ
h5g00gj2mBMjop0awY7+PdgSv0z+M+hxX8md+bOv14WDKnDwM9keu6n2x++4q+Yz
qU4vXp//pXfeahzTWbYLs0qji380OjD3fZ95YCQDArzIfLLj1Evlyi3+9Q0OjXdV
xqHjW4oGgC2PkSuBwjk3tFZpi34/XksA5Nft2jAXaOgMUelmwGFfpwG/EN9nc8PQ
G/NUWNvJeUnMiuMJ1u2KKOfGlRDJjn+zoFdpvsHOaM54tbNaExZqEGdvtFH+RSoR
aQLtHiSv3V8YESlYYrwrWurXqNd3Oei7gnLscRGbtwHlwx826yOht0nAChtt+XV1
0eP9ivbvUoQ+2ZpYyfpL/elAaJh/bCAPIsrCwD0T5p0JZZBxX14KeWV0C0q5LANw
ifB4iHP1Uq2okSMz6SjmLGeHX9KLnaEWcyCeouzzVt2soM2y3rprwNjRHAdDvRSp
4MQu5wwNpdAuP6fPW0E/m7G3vihcJx4xrqvRQyOqE7tpz0HxYY5uuyPKTAvbsyeM
b4qsYM+tGvOIGh/6ANLEcSkikkVzDM6+3LkxHh1YDWO5AsS513GzK7jxDi9cCpoB
+uRipWQlPEIhRkl8xdjK8LtjQQZqorKbvja/PWME/0AZ2ODuOGFKpxbqN2C5auua
zRyUMlG1kAc0/YZxg6TF2JSIZNwsIY9czZ+hL5I5GuhKFeWVgswZz3o1gTobBtKb
R6cwmG99tGBFzhDWeOa/iZtA+etMUlRX7lxW2VNWqM9Stk+CySrrDE2pZpuMnzfh
Bb2dyKn40bb7ZHnWAwn452Mfq3lxiNwD+lu+1fKHGnBR+I5pTHYmagbE4V0rh8Rn
f30Vb1N3YAMS3WpPL7hbfb1C8HLtsBOBlw4LT1ycwiS4qZ1CKHgYc51vJQ4fO9Lh
gCaEr+v7dQlzwWuPMq8t5WNnT1ZPsO07TIqrmLEnm21ZnT3uhsEpj2Uf5yYMeGVF
nLu06qE4X0g4kKO3HTQZo2sEQA0RyTMePXnPuB22ADPBGGPtfvmKY/B9elyBJ44O
4rKfmcHbDJbk23wgjSKMpwALdjSqb3uXu1aRizI/prGlnUlcMFPx/FEwvuf4QgDu
r2VK4VU/eioVfN/rVt29K1kXCjjripQGADXD84OLA2gJsMnFYe2JktbsSfYBhhM5
X4JpZVxRCMgkWMK0F889tuwlIOs3MvGhQHdlel7qfYXkkP6IK2qH9FvV0hxmFIph
eX8UdUNbzEt15LLmV35pqqg00Qfi4hRruyaftNwzR7FPnwHH80evdC/6NvnbseOT
uB72gp51d8EOW/eaqqULsGLX6CV+tA0nXfbmgOC685lA76TR79d+jXxXc1Y/J4Ft
jsHVy/cKnak/UUxr6qUAmVnFAWm6d+XEU+iuNTl6cTghaA3RXMEbDO6iObBaZG6R
D5ae1tPFasGhW3DhB+n/kOVtWHtS26O6vlCtG5/gRqjJLz4I4ya3R10knPTCG6vi
EBr+F2QAik4neQ9/9rAsW0ZEnaSBEucZYU4g/frAtiGzI0WrgnO0gFpbcTqEN61+
GWGjaxnL2KFnR/nxhpTznf3/jbzfiuSke3xoQHyy4OguKRIK72KFy135RwlmCruV
daKsQHHbCsyG9IPuGqmPpx4VBIs7a4q94eTBhmQ5b1ncnLnJHfF3AM+W0OSMTJn4
klfl2wsXm0y4toSx+agz3FE4j9TWfWO5IBEKKqHESkL4ycDoX3BPYAYV0+O2Hz+k
2XbRR4iFzSgkrdzoqi+6M69pFk3QkWVXs8gUWdOsSMx2RlvtLhF9hE9WSDqmsRH2
0w4gGRGxKDlDkR7GczxMlTMI2Zx4bnaP3qwbhjka3W7OjZhcyPY0fYDU7Xphd7G6
mw9TRB9DZEMKosYVyq8C4OWlhs4wZXaIINdLZnwNgfQ5bFiT5jVKEAXY8+NlSIkx
F5zVBZvits2I0xAhw52rqF4By8X+qwuJbAousE2RfvMzAD7Yh4ebEh9qj+rvkag/
/jumcFNALMmuPtB6uhXQc6Jjc5ubAf1HW6HivdkoiRS7DtzED8z2lRVYQZmjMOn/
GdJCyB2EazWT/Pu7PkP8bjPZppXs2YOrvmV8wZm6xCuWrf8XUG2BhRq6iS7L+UdO
MrgoBeC4cNe0jPpsQ7l6hyiICdZGLDuS9wOT9dFtngBL0vWJQ6rtoWGK431jTK3f
NkA2B5QkcfhrCOU9ZMyZnKs2Asva68EOJ7J9Ut6cmJ9GFeyznZaA0INO1TxL1AT0
GcnuM9V9eff5nOGtNa5ZeN+sVqQcR0aQThBru3nDYEO4BKdKjrdvAaN/OOlnA7vC
rWU8tlWBadGNUZO/v0qbDg7+nPJYUEoavWKBG6IcD2xBamIwHIZuaLhtw5vGvMwP
4hJp0XUuDzvvCZjvNpyzR1lf0ZnM3wL7vMFmwWuhtdQD0hnRxx9olMVwQB8ssla+
bPuYOvBdba0GdIzNkMVlqy9YWyx/vqTZEpI6Kv2Yk4AkS8T9nZZh7lGVbkICyAZX
KKJ8rWXzd6oipc8J4YDWny+b7YYZKQdcGueALUj7aUo9G57gfPHNHCxpPORjE0/N
9AahBri72Zi+kAZ2HfyjE6fespTq4q6nXmFJR7iSuxymE5bkcNnzyUTNcBfaCgUf
1pMVTwtnq5UJLFb9Spz1M+Qy9vbjIoCLX6y9Pc0Yli9pm3HuGgZQ2KnTh2hVLi3S
j8nrv+BLpQDzlGDVQ1OmfOOhkjtb1U1onehwlaFw6TjpE4OHqypwv4OE9oGJdVSW
060bNaCkEemLJMTqpb+dDLwPfUFtxPd8RMIgoyTNmQdSN0x1vWfmK+5TU15UTTCh
nd6hDDQow2Leub95wInDq+t4GHn4M4JTU+4bKmLyHAMAJExp7yaV0lSYG6ImeFDL
eOEtdWXI6S+WI616XwVu7uxLr8ftNrchfKjuirydRIJ2N99Qk8HH10myoO2uA7hA
a1CLnHi4rT8QCk1iMpixkrrnLamcRDDFqJHmZLnRrnD6AmGa0v+h+2NwWiuxy5Tg
a+Idjcvu1+BZq9mzg5SVhnkHw21m9Dtsu2vdWfBh5b8zfON3k6brQTfhvSBthaOm
I7yTza+gLxc4AZCoh2Fs5sqzqUU0PwSXXvcnnMuEPlK+5mzrBRp1vDJQAoM6jaE8
oRVmJyOPxYULOUaIWQyZoTCeHqIHqP4Xx9pdd9TYOTtYpr4Tu2IsBcyEv2PQJbzi
nU0zNbZrd0CWkXM3EF/9IOvObyzE/bpkBeCqc8AAg5ZWVcGuPsDxsEobeJhTJ1Zh
WAAAzyFK+PQ9LDvXbo7YVTgZk5lQSjVT57tYWEPLx0gd5dK7ErcNiOeNBvYPjF7i
POcD+kMZtCqoymkQUbJZLp24vodGs1+Ywl6QX2zi9ppfN5m29V/0pC6Lt+RbMn7f
cyODQjA8mL4bgQPkuSjHEs8ojAT7H5BhpWEqQSbpVknouw4eNZgzIoa/wLelHatC
SuJLoYY0vhZEI91tFElHeSXdRIerXKzvOcHskkt/KWXDtz2k516b46lb5z49nzM+
0rWnvg3qS4GcdvaXxyrLqZcwW3kG/7IPOAiWt9pdiQk647KQaSX4PNeTdXl/LxYB
rpTmLTWIAtlU0lxQwEDL+axHzXit1SqXhHUr0S9jyeo/tujZtMARmEH1Z2iryUik
UCdSg9JVL/BCmczgwlutiVNNQuzU+VKIPBosEIJ2JcTJ6XPOLnwZLJWnxPLy6FQD
V1io4B37VM2Y4c2Ymh1TW31MI25aGFYXCoI+Z7Pq434vd38Bmt91eFl14sZ+vkFk
5exTQ8BxJ5KelIyAAtf4OhleF/CLFGD4DJyh+Bpe/sQn5x89iJH/JgllPI4Axzcr
UiFZlXgkWMEAzppjBnhGFmmGTJBJPFSX/lji+dnoJvEC+V1PxnraPNJEGte8uIDe
ulNylm7vb2bbEpoaib6JtPDc5CissW8FAF3FzA/+zH3vnmMwBAI1llsO7ljuPLQS
+gbvGEmp3+vLaB74PlQp8ou+nqi+GiWTsXWOYhb1jHxFzVXTFzRo+/t3lEWzCK/N
ne07ZwP9IgQYuWd6SM5Q7vGugt71Aie5yRgc01N6A8QESxpdfALkKGCFPae8bM5s
yL8AC9z3jyDJEwHbAUS9SOAeJsoCr97Cj1E/LVcXU93AydAmECaWDyTsu20KnP5h
OO9ibgOR2BgD/9DOpRUneeWl7W8+fY6qp6kNQN2mQrGYFYTE08X4ShShPavw5L4U
/dgluemgOBv+x1Dvz07ggcrZuekvUAXNb7g635FeCl3b7MKn0Q50BvqJmkS8OnMl
5E3gUcUjfeKYhA5Hqky2Djt4LXHRSNUGRvUmrdLRvFo/ZU1v2pIXtdJe2AertOVC
OsQWFJDFyJQo+TYXnBP86EdwOx+SCWReUi7NAvKoJ4W1jo+fctIlMEiVUQwvCP/R
Dfl3yit0d3dhPc6o7W57VpWlmCG8BF7waVIdRLC8263nntRDgOLA3o86CUc8VA/M
n5Ja4CIXmuBeltCjpd5z8gkUXnuMbg1LatWLL8Kx+Wa1Y3ulHsK1x/ZaiMY0SMTO
7Z7V/F39aMKtpSgjnQk1ABXd7Z6ABzPb9PxacIDgVyS/wXWKShVzzi1yrWKvJpeg
6i4WF8nXjpOkDoc1Pv1e+VSAZoVZytUk9yU+CrmgjqmfPMwWLTlgugLlb8Xz1jTe
pNkSbxpgHSkzieE73tkiWbAXcI7OCHg572+XcsIZYfjeJ5mYJB1bzAw+YtG5OQh6
Old/zM55LhyK0/WsHkOInxGcp+jLt5B+OCfucZSHulR7k+xZysB9FACaHcw+INTg
i+JZf0eqkB8S33DdlpOZTI5pl/hcGc2+ET0qlfLAyqaYUg31GR6fLPk498N06VT0
AZDJrfzeD26NGNh0Ywd/9xqkx57Li2PZ1vs1coEtftPoVOZmBjl5rLduHPjcP4pT
DfH8WJQndq+gI1OZzmdUrm97gvXb+W8mZOu3lwCc9BKVloyoZ+gp1CB2pt9aZbG5
CTFEMDJau52qCci4PsRq8wh6Qt+Q67d0SiV3ppWoXuTL1SK6VbDAId+/XMpMbGvV
GE7A7YPxkaViDldhACmoZYuGlLJKNchm878hUSvdOs9Wjih69vYykb9Xp5X0stni
8yRLorOCeej6jVu44o5ICdqB8BotAJTFcxyprIL0WKc4PUeVmW0mjgoegKgP7hbK
x6kiJGZTOOVwBILVP6SAhKDBJVeTxg0Qc3uR/FCvorr32Ba6FXatuQ4IslU7kVSb
jOmQD4Sm6PUgu8z0VMNR6UN+Dwi4vh6md9aJ182bhMWv2UvrPZjnCj0bLH1IN67+
QaMUhRi5/d3cz1Jt3kWY+M+H1+I3zAMVrhGquwYAJP5gHbcIV/SPxOz7jqhLShwE
yykFQfdvbdZdqd6kcUJarC+YlUR3TAKSFvE+WNy7C0jNFPTlbcgqKyyz8lw1bA1y
o3KvlujESpdOJxb2kaM+7R7OCPObfjMZ7Ya7wzhk6bzIni/CCqlPZ8NKNzcSCPlZ
mAWLGWvwXE/ormkskqc4dNaIvd9llu7eEdhV6HsV0qvIx2JlNpFlP9ZD5TXiGvOE
3p4a3C6CpIXaTupyzoKdgk4BCHUhsazFcoOMTGhMr61oUaykJTgXxkU44zs3eoQK
/i1QwKufsxpp3RHKPk2//fzePd2uV6G3yVEJz0qj0eBRpw3ZCn54xmt0Fj0VgCpj
AKzUUphrInNgNMsQyIUDDG/RlAjEYzqCU/XFJXSX87IA6QQEU7pQeWw1ROpGg7Fj
ndszP7Zqch3K8WybRlTIP6cITH/a/297AFmaPiFMZ2mS59HRLTNLxd4LagNTAV2x
2A0eHurfos5g3t/Sv77rfB82h4c6b4B/FVvJYbVN9CoW3b2lQ47qzMJNoMPR4IjS
s7vdO2X9jky6sQM3ZszKhsrHxupt9EWa9yuyjfgVeOZ8yBo27/ozkhLrJ5uPL9Ba
nwZMAZp08wd3O+rjclje0kKvV4rEEl0IDOaY41XNMUq7P0l922sad3A9bNwimMih
uErqLWz+0n18LESXXRuA/mF1sK47wZrYqVFq7temKoAfv6iBX4tJe9ntZAlloP9w
wo0MIg+qF1jrC4n/1sAEKlVzT9e3tvhL2m9Cx13Yw0645ugltImpItoBoQ9YNBCw
ZVRLCLN8vu/kKua5BgtGmEidjZwKANhRHAl0ENxAGPqkOkQegXVY+N3GaDi+CZik
/wiMHZMkdvmqkjARciv4zkpr65uTovWPqV51Rf3o1yBz7x05l9OVFmf6d9eb9soJ
8PT7394LQEnftgRy5Pc9BwSFaX8365nhjTcpiQkrmXhHxtJ4cEHlCJ6pUiRDht5Y
dI1+rYsS95sC2pOXn8DI/cVoLLnBanDfVxgQ+8wtAaLdX3yp1rxIPp8bWYcfg8D+
sZAnOp3FY9mxMxs551fCH2G/oJnSx50XV121/eto2xIfRllRNS8KKFYOPNhqDeJ2
G8CrLhL/wt0C4kIURn0NX2ZD+0UUdK8yhRAxeVulDYT2WhsEM8AuKCULLHtTOdFM
xyfnCk6j7rzqkgqmv/uyppkVH8jtOe1VKfWy3l4bnC+NvY4qd5dQLVlM8DBQBH80
CK+S1pIWuJeIkrhYmpU0u/f3Z9yMmx4aPdqbqoM7gzYMqsp2sXupn0Oy3w90bjrY
dPPn1x/CF3ii3Y/bjSmm1fl4AeXLvnHXPvHiIyeSHNCbMpFq2NSSBRcpeQbJYcg4
7ZXPRu0HIw1W5palCKtt9c9Vj6JtwsdIFdvw3x1MCzjTJE1Q7UpHWggpSFHEOUBs
JPO1mFuZTzKzDvlDf/U3sfeGHbLjRTxtM6VIQ2IrMscGraWgWzTjHjiMTmhHlqd1
dW/9AFR0ShgVBDTjQRN57jnf3HT3seEiN/TjPN3HOZlgteGXLAPq8kjzBqJIBtIF
TcvAnYiWVkRCJjGx7f9orjJ8JLU1g+LEqbuffq+olKptTsaPUcw+Yvl9MRRfeTOe
47HasP2uKX3vUndIrob6unRWo0kR1MOtQGJK9emldi6Ymk7ZYpZ1BsgNzaHv/Tj6
I1jOKEKiLuZpQC0GvsxL/35rU2OCTxkw0Lqe2wI5ixgFDTFzJKAZJtxEtENTFNXr
sQY1BDQlu+PRWFR9KDxpTDzLovvWlz+yZSOE5wRKx/Ruc0+6JVYGpw71uukNUaf0
Yv0xmH1in+IfVfq1hqkimKj2QoaahRnOyfHFnupBiYvT1sTB9Jf3wMGN4xgjqkd0
jiS6spUsiEmrfi/Hq2qP6qTcaAJ9DaWlyewfUW9b3lwkwfbcjLZw1vzHByo6FsKU
Ort9Vf1m4WJLGl1WPV/u9+z2HZwJfd9v4fwsOYZia8d7cseH8bXA5ypudphabSO9
Uzdo4lRro0bnf+v5Y2rWYt2Dsuz77hjeWF0DrfxBvDz6AFplNTgAUVYl6U2CUQsO
uGlwcCbAN7BkO9y0adFXi3YMPBktSLcqh48OQn99SB8Ql3SQFnWm3+gAuozO5dOz
kQLgY6toWgRKVUf310UDTeskQ1+E/MD+Dcp/EwtJ/IUJUjgIsqqXXjAcx1S7YOG9
RpAyqenvXXjDncR+FLPhOvcsbGN6BJI65yDM9FCZW65VviAogqEzk1/rh8VvdI5B
T8U6mZL3qrQntwDJCHn24lv6xuiixiTEG9IZOpWu1BvHh9nZ+mYNH6LSeo5kcaw9
W5qEN99xIwK7feorhFaY9Cu/zgiYssalbqNYeckX49FpPmi9jIyCZ3wLkvEjg01V
bi1rwA4gd72g9FUuteNfZpFesSGN/h1ncqHHxSGhRGcYbZ5EhzF0Rn+VA2IJ1wss
W1Mt+qQMppo6Xbq1vk8asVmelhksOrxYv+JLG8D0nwhvJN4K8PckbtAdmq1oQdtD
P+iQTyswDR+LPm8CkTLwmwLR9HkBAhE+tI7WLhYS35ZMmscY9XDnXWovLA/KjFdC
fkI5eq08xeiN+1lof+IkyTJXaYNh52+l9UQ6kM0hv9AQqJhmqhQy4hrU22KCRGBu
4VrGyWUGR6S1LWOjbusDRQyLFL0dh9voOQiCA6nZP7nZXBKP67IC5cfVVkPJrJz4
Aeid1K58azdWEIGnXEb3Vjn+6iQnJxyfn2ja4bQZ6lra5+i/kmgcMc4AEmi6FSFA
XBqaH9blKWHgc2jB1x5DWPVgdIU2Ilh/jI6RDP20H2ifPOAg2p/xmOrXIFcn2Dv3
kCucJiTv4T+m6k6gBU1FvsDkT1q7ySsZgMCV6C+HRfoDaAzGHO8UWS6MVZtYJPp1
HzHknDeGgUy4x/hTyUXAT9ugwXBteID1YEHoyxgWrMfU4NA6vKLTesxLM23BIb/f
triTpAuwed++KLKNLFDOMB/vf4bS46Cr+47S259pbdW7k1moQ7b3pV8TEUfT33NI
ftFfbUamcOCouOAmrmOGvRgB3jyeu0owsbWr/I+t2+o6y8B5KgHwnz3dMZ4SGeLn
Jfx7BC2cJ94INBNgmmSC1e7nTciP3TeJElGt9aTVMYa9lCjNBHSWS5BM6EVRztfD
n1jmkpuwURelfIK5Iqu8J1ESeXNvT2pxH58JyTaSbmLmyTaHTNvwWoraKAf9Lbnj
Kxy/jFFxng0a06msf1aAyP9QVlaNJC2DmtbDQkZDkOqmHaobzrRfaomFeyMPcnHq
6zz4P0lqEJxdctZZ4SDGY6Xn15d33SlMrQt5kKviQrhp4A2GCPJzMScFb9q3ZZxc
4g8WMXtxfY19B/KbmHvbVg5I0oAKjZTFgI2iPz4zDrVyDQxakHQnbsoJi3i8Uo6z
VygkFTOUYzX2wH2AijT5ySqXF9o/nWLOCkGspg6JAvGDVrT7VP8JtH2ET7ODkjSf
v1JxGDl49hGJmPnvqJ2VbccP+fb10pfEYDnV+CtSFNPmtTfqZ4KsJ7tAE4M0zXNj
+9kMjH/yk06ikLaUTrX/7LcGqHOwLHjA8PA8Ih5WFg8Uie1+vEYHYHQMYjjOxKy7
ajgMm697BdHjtkoHLOrFYmyFVjzkabpivqBNTXFl/mCBw4o9QvL3Whe7Y3qjyZn8
k+myhE4V18Owd0UiNISRJHf1yMDJ7op6hGg0sWZxMrY9Q5WyjEsfcyuoqhcx+0W5
xthz/NcOFLKkGfUaUrlf8Mq8KGSJo35x9nZJLrjz0ev2gPCqxynAomO1onpxUuJY
AbOJd9usispdJridolxcGe8fJJU+XT+7hVkS4HIavV5JKtaNCkUUwHzDW4poiMda
GYlg8y145qwabg5N/GxNHCfsW41W6j3ZnsKy5iJFuHBXhu7kJzarB+CqfLIo76sy
8imXoFXHqEqMONeq3aDfYTMrwh/Iv73hvra9DC5a9qyQdytYV+xnXtgLJzNrztFE
b6Gfh952hzL4moyj36MOUvTqbWyH2MJuaFXFICvwRZFQyP5Ml0qgwe6Lzz0n2Ix+
FrUAbrFj9IfX2DfnsqlgzlYLaBeFVvc7ChV/lw13Ho7a/n0j5grgpuyC51V57qai
O6NQ5xSJaxTvVxgvVmAfHa3FKSx+qrfXnOOz5qsHMJVz6Nk0hzXXPeEl+/tsM/7g
rqfWlbwnZfwxDwk2SVUjz+wOH7jXjERdV+hKyN5fTIBxJu7O8a6JgIFlyWbcsFjG
w232abvv9lonuJI99rMBvr2NFNQgaX23T2RGgu/cnNE61xnSLJoGH1fDt8WzrhEf
88x+jDj4NH/7NSeSOkfjmnarFhW5qZ+QwzbgmVD3B6nm4TKKBcNvNZ5LH0l2EsTQ
PzhNt84is9evwVkH/IcU0qQZLrOCrBbmAE31uMT2pzQVnArScVlM+Zb5I8C+/HCN
DrvZW++223CF7W35fg9Vl1UpPzn/ronwHkUAWNOkCFfCbzrBG05nNI4WXhznicC2
070IU1eDmutQB8n5a1r++32c840RACAlDwZHCJAXv5GE5kQqnW8XWqj+NSZIOhlP
BdFuUP67Zl3TL7nrQkohvH1UFUJcKk/rizXVwknNqlfROQ9rkm4KpLlJ4oDt+i29
E8y+FD+OmGlL9TfIZS67I3Ddpi7r8qWF2FMlpEJebO3OF//m9Ag+2D59Wts5XOPe
WKcHXvTRu0PFXraZVpMtZMSsRDVjh+13qB0L7mZu9PG8hXK+aV/IxvMNC6do1vfF
iNh3FdVjvv8Cvy7vj73qLVvjN/7zSPEyRh58o2umyo6W678svn8ZHEzF1jxxwTaP
dMfV0SjQAwFXLE0inAW49MeP6aXD9XeKa/3mk7jPG6lXpDB5NLHE1HisnX8+oXH/
liU9CPLKpCZBbCq9c3G/bZDW5aXto74v+xMwkCb9bm/L8IIhPz/w3NSIevajK96x
0plnh53NT9YxrR+FmOBxS3pQb9S9XTQsWIJWguDpoqS5aL39PaIjXyJIeaplr4Km
MQFBcYX6cmnZafFnrxcWHqv51ATAhwZ1XPYMviSD2KiToxswkuHAco6RhQcP0ce1
1kUrUa6m28AVDuhRlE/ebg9xF1dAlwzL2EGecbO5YX2tLK8nS1NThBgbcDq/Vqtl
5za0nfvqZZpZfS9icWLx26p4PqA/2BdDTRboYdXbV12JbxAZUvDyY7JOicgubPMc
V14laHogj5Gh1MHL5124WVWs3JwJGpx1ogpKSLm+BdLlQY6FxDd1jWUH4lsVOscY
S5/Q8pbd2YOST9IrdlwzAVxSbLfN8m18O7RnsgA9ayZGa+WYuqpJ5FohDjX8pKss
0ubTxxMqZ0KbRl9gIHljBrUXUrORsDWLlHi7da8Kv9cKqQKo6T+g9vC230DAh0SF
Qwe/yNGGuEIgFqEuXcB0A24DOpkjwLS8eiyybN15ytGNTGVLTYwzJUGTO3G7zhkk
RRu1nfogE3bcQWZ8Cq4BLIQABsgBRCeMkPNdr8floXFjBelFwNF5rsp66DIck8MW
0T9BQiRbZddvg1Vwsc0MnqaZthJUGazSQEX6aXRCnBD1OlO/iF76emL4yeYIL+w1
pCT7HCb2i51fgL2GOjw/12GAz6pOy4rF9zMnVEwf7BueMxMgRyyfqvN0vqLI3zKv
j8JAL5ImRQa4AfvFg87ALVJb23rvhFY1uTgSyofT4QavCKsNZUcXtJ8QPY4yL87e
b4w6uz2RGmFTyX2nlnHaDxn7LRIVfNy+YKVUtGBxevT1dmIibnXRbRI+SYu2WTi2
6ylLkn1P9E4TSJxASO84ME2Tj2+L2gOc3/RZKG4UrrJVJlyG4+sF52cvRGXsbISh
j2U4On0V1vRuSH073AQ7exKc+H70uAxUSEK8KzwBgFMzsZjVLUGCkRo/WyQD7LtI
vsWPE5TKijddPsgHwlKc0KW4Bt6fKdZlaQKukhy3UibW+Cv6bbi5iLOhIk//6ZvU
+3Z7I0tr0wZ8B91HXkkyKtesUGVqvZoymSSAD1KBX3mNQYdCHjf0kZbcvs060qRQ
7iHf5H7u5IynH2JIajOlbxIoC3VHtQ/brSD6ymv2uOqyhM8uVni+oZwYSOP0iECn
Ljk3pBfHzDFC2mIo7eL8qzAmiUydV1jVJyrYZA5NGhVHG7Q7mrUV1c9zmauasqh7
nUQ31yhCSuvSk1fId9XAZ1a0nuJTZOO5MbJ3kT1wez3Ji3D7J2vEyxz1/tWTaBRI
nEASmaga1nU138YJrpL0EUBBbqmci9v/CFYv5Nu7Tt3fasP1uxHPxXnBWZ3EfOIQ
uB4guc+0qEilb675WU8d/PiSyhYWLqnYgvKEf+GD90gZG4bij4kwRVq5IKMdQpcm
c0MmMZin0oA1FZVt4KL9oN06pK3PSSqdEHVGqLrZFlq/MHR7czPBNQxWIXvUDaBc
ZwKi0dPJtK6doF0GJDoG5wxo0bGRXZjWAdPXtUiu/01PuGoCqeY+mHj98cvvEP/j
Yns4wEYZx4a9nQwhYNktx/RlJgVRlPu+k2nyZ6Mg85oJT5pf+ZEdp8DpZjeLehEG
1A5CAuBDDt5dibyHkg/XV+vKCX3gVrkMZMRf+f7Tl29AUqFGdbocLzKAyBYdAMTc
HNMGJq/L3VuSNZlwuW4KP0FFh4AEmXbBuzyXRQBuMO6xh8P/P4rASsAbgxzXeP1M
B8Bs4ffBNCX38Y3bNba13ScNLEoNudmy8kpHMjDtkO4t+R7bXrtD75d/l2ntCJQw
/s+OdabEWty2EyTivv7LUcPoQDquXeYEqUyZxycEAEOT28DCWv1DmbE4wFjXku3e
ev44mjbUh71OyVeVfYOjL7tdc9Z9eg27TKNqNE0jgNlRksRUZnOrd1Hl1oNHqIKH
K9xIG1m8Qrn3VlfrJV4+4jiOsaFpx1Odrqof4rmfdbZr+nkwgkEtORpMJHCd1WDx
fQL/6gNBS81u+42GJ8VNfM6ZmkNoOMaPAAmBtKYD8tZmoroqngxsAwJgg063L1xc
X95YWCxy5qvMnuJBAmYMw3IN6WMK2V1pIkOH6cMKokhK6AU2Jd0EJbTMyLWv4mbK
SM44AIbSYPfJFHNhvqnnbMeVB8rXHNxHJ6j1JsqKmv/1ppkNbd2EF58gUUFqhKUj
e2j6SH1235mllgdJVu5FnWfMFiLveaNaSrsZa9XbW5ffV5KT02zbeCls92L11Btk
oTxlwqsBI3+ES1f1peNE7c6+hMppVZWFlvU0iqQGr06SNergkiXG0xrOGkeVMxtP
1sF0kBxZ+NaKRaHEOCEqHucl9xoYRUfnVVcUycr9A2E7wWBXlPamHhugJfoAPOPO
d9dDxGTZFRJgnSPDOuUbFX0/2gxfpIJHFWf4MIjrQPOecWD1HplHtP4Gdc46kvG/
lBEJk7WttHBOE9tziF0k8nVopPkaS3NlcuKwKK0j31wqcK/se6S96A3mvZl2lcQq
viYgNgdUiQWugU4f4G+G4qjBA+aWXged7lHNev7z7PHsdCWyecnxKkHNP14DdPc7
`protect END_PROTECTED
