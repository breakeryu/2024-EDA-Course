`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
azZVahuXct/heTDSDX6kThPoWAIaQKlMg0wFzq3rljuQFdKXw5Ts/3T/XJgn4tQn
VOYzRpQNC+xvgDHobCWhY/6Fh4B71Dcsx1g3BSDKZ+VxtIvmkySyjBnhGaIcvnwP
PdZMbXxLRT8TCOzMRRnCF5IZWjZcdtTs9w1I2nbEdvvPYGhQQ2j4qEXhwvBP7N8Z
B2aIAFOo9+NPASeqiR2tRKqNvFfH7mIiNc8OUQK7s6H6qo1tTgj3umZwMhGE7/JO
swRIL+yj5ekG6981MLWsgkutuYpoJPiRbm8DPXEu2m3KgUFm3fJUmYV7c4rWakvw
/9S/dnGqvZ1IvkxDAu+GxuUd8eHymLRZ94W0wLUEj+7eBTvKlKYQQNG5vhPLWTrA
+Qzb52i6jI9Nb8jv7d6W4oKQjpe9THWLG1UgmOES6YR+h8lopy0jAwISayIj0896
vAVJjPBKIxKBoHHvbLFKC4Vlfc+4+B66P6k8IwBRfbzl2r/BAILWGpEG+lyujRuL
/tLDMrexiR5Koax00LgIjt4k0qk4OkK9w3a8lbSSyILYpdutzevwLjQM7BfWdHaL
A0e0a7GXey6+NsPc0uFR/ipVaiovAB8gKXJWeXvzmYJV0meAb8GB+5CLha8FKlIZ
1yQI9v65hvTVEHojMbkmfqDPqzp2WkLpneunOIH5xi3h5bSXibLXn0wNPAH9PV9F
SMzx9UDfbdMiZORjxzHH2thikRccMZ0e3FodaBJlk+hSt3E2SbPHF3+uIKJKXuBM
celDXW0oye9YTLT/xT0JrWHwQLPzLxnLToLtTiCeKSUTawcO1rk2DvhJuR83R3Tc
FfaHN6us2UGkp+l3QjlKZ7NKBK2hmaec6YIRM+gkvPCGozeohbdRhal2fVGCp5XX
RmYnbBIb1JIeSY7Qbc8LNwEaXMc9J/ZMx4c10F8C4Jf/Il2HIlVipUYtPcAQkLFJ
uIIGPfYN+6hEI/G0/Z55ILaetPjlbV4q4nbYVd/YgwJAeQTLHn7IJ4gud2P1cHDL
7ufx4ufi3a2iFsXsRZKvtvDWnJHXWnAICxKahJFy6OQdscq2ZxrVIYMo0/euGhJB
CFmEdsnvfq9E2erIr5AaSUUHues8yqBEflfTBgJaZ+52Rk4l71Q23oYdJBbwsY+y
qMJijW0/UQc8z2xH2P60ARqL235Yf6URfDjmnFUXdc/HkJ0LTUGkR18Di8TdcUpO
nbF2oxi9mO0XyEPhwcZB5uxe2dtZDYrxQgOhEjyPH6OuXOGw6at1ZMZ1cYuVJIHe
HnzenbEE/8mE/1ZsKmUr7moqL3Kka6N465ErMxyWiq8Y4AU6d4pgAU2YQk63B59X
eKWcknII0BTxFqYos/Ev430WwPzJMbAdqHx1wdlfy0R7Efjj9H2afvr79X9mSQVH
/4IrA/UKnZtaGiMy8VrbduVKGVuHtIturqE/rtE4GvtTn3SuYC9JgWm1FB6l+Ipc
/xwHbDhkbQTSu1z//MVqzsIiGH+fYPSwnlb5fnpvtXdfe/Zly0slVdHeAoe6XJT3
ze0yXAWCaSS+Lbi6K9CBIgrg660w2TmqDmHwmCSkRQKrB1VOY9MCu23MG7daGIO/
MBziEIu5mHAPunGBYWPgWk9in0M47+nhdqOXFaYoDdGCfOonoEHZG01Jg1ucUGLf
cuS5j+kfmmVQCS61tRj3HUrhg7ukJy3tQeUhpa38pZLXi2lgjdnug1peAQHvLSN9
BtLls0j4CMrfSbl+h4dOZHCJYpMCVhBYpTvtqis8VrOXUPSkRzdfHJSQT9a7b/FG
O2gt92p38GyOh+vwjFNouFCd8e/9E421eTlDbdIT6d+GEGpl3GrgtqzXuVfDv1fb
DTtZhZv4v+wXncceACLg9FQBfIpG0SlSsxqB3TClCPdgDdofCjtlQ3N/p/veDLVH
RaZPUtobxauroSdA9mqIdI1FyrMNW3pF4kyH/e/POXbcddu1X8GqLj+0pxcMTR9M
DvK4qmMczMu16igWtlFP4DJ1UFh+5R8hd2oUN8Zolycu8hb78lz9BtxwssNfwaA8
x5y+hG0tIFDJ7t0gX/0A4a5IQjrmEw3mwSKeezaZu8i0YgSy/FUWBqkq3scRRKeQ
6ux0UOmOy0z782NR39sc2MG0zVerpX6klRwCpu7jzGCFML4PBOUv2i/OUMla5sje
h3UA5Q9NpkOlNVLimYA/2h/HvVt26bBJMKduir4h4qchb6osRyOvYDL1gal5NfXj
yGQuFdb78XL/9dntX3RATY0Bn9fHSIeWda5odTQOr8mXG6VJn2UyQtSZVUzXdbBN
v1ilq3z0sHxC4Xp6sowqKEO6gFbrj6mrgKhXMz/RJA0nkZoL/+o9LG8zvgAXo3pB
54LD9/g3c47eQF9rx7OaMQ/i2zabfjr0/CAcfarmyWXJmXx58iysQlkmtwhrNg8e
RBfYr5rvcWlCz1SQe5Vbpf/9LfmsbHRDGGXlQAXRB9w7ad3WT8Q25mM19003hjGx
J3E6UwA2VG7NNAFvxpqI/scwfvfjbUfUFaUwUTvbySI+jC12QCd0S3ci6josqAKH
9H3w+uIMAK9OaucrnClCazzcjkPKcC6m/Cu/JWP7ceL51nhowcX9TdPvKE++0o1r
NpzS/kpXutBQ7/G9noWbUgAlloucNVZVrYWutq2/O1RMe0aqk15dhOj2+7xs5Qz2
ZQki4FRD6aKBa7TQ/Spay2RtPIhLpQe5ko+hAuUFxT15vJtNKFZFLzdCsMfFEo7X
rJRqLm/wUlqrmADac5ppRQpYu7EvX/l6C8I3NLxjiYvZRm+JEHyW4+FAgE90KZhF
LapZYZPlSh0LELfxaKyojKsSPJHPQDw1BW5mxdQBk6E+lB6Uu72ZVflOggBaZ2bF
Ye8O0t79kswa6wRD2GMQ1mmI05Rk7/3MrbzIKBfM6rNdA8LHt0EOoZqiXwUOGBK6
vleI9/D02dS5F6szrTakcI6wIvuPL6wov+aD+lA9tGX/S/zs0rBXm5wwQn9iWrXV
r3/1UaNH1CFDm0SmFwH2tTaqnhY6S8VdxoE5mJB3N9VtBfx54Gj+aoxl04CTW/Mv
+21ejDdhHpXaOVRxy9BKJhOshdtmUJJRMdZramHKe8fOxEvll/CnxwhoplSKraiR
aevlo7sPwccUwSFJ4n7yyKtBHv3474+7lw5tUamrDnLWw9VAPX8wTUoaHps18K5R
OOcZR3TFO9GiGIBVy2v18ECF2p+fkdwelWd+nL+sI62K531LV6doyufl4yEIdmD0
7UIRuXnJXNipRTLN5S2RRLiL82glBIqT1DtkFxt91BwZC694VCS+mVTmCALTZgVQ
vMfRFGhwMHSCHYZ2hg6EwcwLMgs1zTuhIKyC+RRbPHmKSwoZCocBSLjVB+XWfSpo
GqGaqlNUzR2qqL+4rdkbVUwj4l89XKRQh4y14MbTowPYqbu2ujSLncOcZUdVGTJi
LUhButj35kev3TOjjSWtSk8LZAzjHIkJWDi2JrPWEbYB2Ve68D5eksQ8NanwMcuP
ExIb04teGiRnnIltFkaD7JG77dIoMd0/TKoY8dp/hocTd+kTeIm6AoQr3Hezpukb
JB/AQLE5UFkPqt4PufH/IuLLT2zOtypzXX3p40eeharjlUpHxijzA6WE7NIZMecf
ei1dBYWcgwAxJmxy+5Gj29Luqmo2jiWNGVTU6RTmtwYJWCTYa49lzoXGkMA2y6H+
/5TeEWv0KE8pUmHiD+jQY0AiDBSoC705+EaF++RGueH9IHjxDWefceaXypXj85QL
zjVBEHqduIvdpywMUQWkhzpWL2TrfUbBH2WDlVKh0QIWiTtxkd0KK8Vfn/4OvKhJ
Y+t2QduG9HRRU1Gd/kyLQJC4jkwkm/5StM59+0nIqK+SKvb0TXhRn41ONEvo9XgA
KD7KTFsw2K1NfEE4qOd1rUGdukTt7Vunsp6WIn+namhhZ80Us1UOZrMnPSpYJbD5
SJaA6CCPwZOqsPHlTtx1OnDomPxak8rDQp1B2mdhFiwgZtgeRlD0A+nvCBGiaqMd
LkxleTndgA5SaW8Mgp3i7877dzDZ/e8NT4IATR2d2cbTSMm6L8B84TkWpbJKEJIL
jpvkj1rwfTl5bqLlKNxPLSiT6str/XbFGQOAgQqwdV+UaAysDbm+90/0XngrEDNl
/uBeM5FRZH10nSB1FHbdsSpWJg0+lF+zML52w5G2BWs3bQ/8xxWZOYxc0wSO1R3P
zAilLvYkCXA7jV31c9k8kpwP6nxw69Xqa3QzO6qpQUzwHmU0FKcfjTE6YlvaVaXT
YNSn7Tl3JxqXxm/eisOm7v5DldOzr5nIVmQoQDm2NxrXE2+LyhHxmn2DYnzYlAs2
rwxzbhPODztQuMd8fwmJMEhqppLNtDECwJ6V+4d4bBxi05tvCwGIzMzCJB1Mjy2f
u0uyY0bwkeFCCln9AZRE/NGaZZuigLa/Q3PhtM/6qCLTme11Zn1ZlWa8gBBDSEl0
ZY7A/0VgPNSTR7DeecKigPw8sxst5eZZai6ReKjno8Z/J9uw97tE/blFOOhLkjL4
jtBrlz2lAwx/VokcMhiVO/foUnv3zLf5zSwYBmM+DTzT3oYkg6rvdA9Yx//Wr4v2
ePJAm/WLQgs5K5ss7suzluKSTSkoxbnVhvSK6HG63euQUizQnLgxQ9YdX3eYgpOg
Qc9aF3Du+TmoEXmfl8vSmtz77IWiiJhz0q19yc+JFgXJHlZYPMVxjWoUZjoMQ2ZI
YnDuDMgilsjw++9chbTFNgDBd2y9NXafnkIZ6bfI8csmtfO+1kmxbnbZ/1T8Oxu/
brq86+nj8Or8TDp3Xt5ZmpP/rtvTv4hIQCroGU9VXPECWvFeO/Os2hzIsRVRmsLk
hZnB1IvM8SO5EX4mY8qZSaktpGGwXfHYgKWZGQra+zmwXgUBEml1NqKHZqeAkw63
0VFu6ZwQNi50WPxD8kR73qnwOoNDp/b2Y51iB3G433A2meBGT5UZKLTAkcc5iFk3
5iSE7A6+6lgIZFQWtcgsVucd8DOOIlPQ4cVTpM0TdGmgRdatv7+hkHNAFXPOPseu
HNscSyxiJWfpAbH5zfXelulNL2jG5v5AcAWl9qGbrGJRyFhSQePSDJhNqC/4YmWC
VaHEl0I8Ol1zzTPWVAOM0rcfdzBwgdnX4ypRU1abqCCGtlnzbI6roxmY/6Pay9Gr
OPQoFtxbKgehTf8geo25QA4ybAIjkY0b/TfIwKpS9ctM0BHtprClgRqJauwMkEpT
O13qzHTHyFLKK/G4yp8mw57nh1WBdKDKqh9Oh4ozh58K1WGhxaF2nlYBnUmXkKU7
Rzb8/G8WN4gezyD0hhOf4osCFkkdLVzmj5T2EJU7IeVzEQ12HwAxDmK9vJ+95XOZ
enYb06xqM5qD7YLoxmcW+gWqAgzE+H7bT0OaVDQXZ4bazLCP2n5cvBbV4honxTUX
uyp3ZyqPC0TnDfKu3KprKSQ4flKhmoyOys/IE0PoPWKKPUFJ4p9SJ7eJDPySC1eP
IqPOJDMBwLU/spalEul074YdGeNDlF0pfqNoh4MAwRYB8k0WQqT6KirCjfLBe1E5
8lle9WRqYdn/OUbMMRd5tRjyW3JpQCuiZxxFseBV3sVXo6lfDcheQDK7isdB9lda
yMQ+90RilsvabfCpjc3/oNyCMxd8tdvM/i9FQ6ipelmX8MgVjmUiPrka64SsBvpH
fg8rhH68oAynfF8Jx1OpEilzblQPdB48qUXh9GMbD5ZXJVaeBjmXrWEHOig35Ln/
82dPp0TIGwonsWR0Owg+dh75hF5aQB0NEXpHtkPBPgzQ5+hXAJL/lx7Bmo47OBgL
k0GbctccWZgFKIVMoiKvIjJMsK/YFaMaqqASjR+kVP+MKZ9V20PAF5/6E2PdcUMz
l02aDFnc6ffAKm6pKN1guPAg3Ax0yR973Fw3sYfAL6dpwJkgMo+4oREy58Be6VyZ
NjOUbgoQgBthccD1uoAUgkGT+FrbkH/M++0sASz5qBrNo23mB9jsrrOtgn9EA6CY
Ol/M8MloVG/WZ/xPDzjPlca3YHYuqdx94S8J+ABV2jX4XAHwJaAACAQ1V/9x1P5Z
pALjFfqBsbwtYtNkQqcpHDNXzr8iwWQqBHyT2KWxny4mFOg4em/J33fq+svWb4NU
AX/HZ7FddhCEArNvFdpQvw==
`protect END_PROTECTED
