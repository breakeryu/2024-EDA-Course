`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94ysLEHnLU6iRoKS7zvHUf5LVkuZLRK0dGKdgUrgQflsH+rWONYWWgbQHA0dvGW9
JSOXEixt5HLXKbJPkcEuJmTwh6ARviO8b3CXNB32blv7wbAPAmQ0E7PIkZdiYRTq
io0f/Id39PNyQ6VchEk/hMr6Ja2ou0J8K6AEg/VtGRjIvPr+G750BPCBupKg/T0M
+kCR1JMn6SYEGuJ7mW+BCDDNkAknFZOyT2MEvsGD3m7m4KlrjAiCOiXFmck5Z2FM
2RHnr1yeqAwnG45wEgEBd22Le4du1Pvp++e8w+9rzHhlG87S9F+PsoHVG8xb14Ro
yYVG6JyX7xANGWzlpBylVeuGBt0qzMUQpCQEbrAirDUyK3J+W3sIVbK4L3ZnFfz+
vGutauDNsSfno9HptN9mZJy98YkZ6oWoqhxwYHTHE6puyz54KY980lVOYiZx/b8y
xQ7qZBEM7sXZP/4RJgVWiZ7BEYpIp1hH5eaMtoudcYpDHRQ27LByfnPa7wf63z9u
lf2GIAsH0rasR5BTTOjehA11ZNPA0THvWv3B3whzNOzqw0cwFqusqMTzuhzO5bTX
F8fglnkK3mWAslW3KGx6wMuAviYUxvqnFMJ63MALI3PiSro/zyyVnkqCpoua6t9z
aXd79y2gXLxfU/axvkSIh5w3tVK+wxBnsaTy6g54TjOnqoGsd8p1bdPuYfbfUETq
dIi2mI0X3FqpBnNbscXQUpkMnmzg8k+BMxnzoqFKikt6NiKmcMVfxTMhe8NIuocu
DaQIGdW5rtT5sTbUfST8NYCn9YvYQETlEJ4qe4eCzdTRm0cK1MfAz+zYWJrSnzER
dBJw+5XQyj/YZzaWNUyVUYHmADFyUdRaEfjq2hu5aw+a3FRs+5IG3UWLlIc8T+3j
B7oVk8I2Htg8Jvet8jn/R8w3pVK1haajfTYYa5EXZMv//EKkni1MhV9usLvN65Zm
5mduX1DspoVUQFG/Ns8IzWmn4B5d2dI0VmvKggrPQnlk+3m0pAhj6LXm4KiH4H46
Wl/nb+QMoAe9AalPPqfmbY7Kkc5kBAKhTsQotUOK6FZddIpKDuDn+LMXNydDoWTV
SBSY812jWJQvIS6IfWSEeweQWQQje5Aa3hUL4xgfWRluJtuatwwMwJusPhGenHfk
lWOKMuRarIicc0+tmlHwm4+o84Q05yqS/qMQabdJvabnH74k80Q7LYUGgA3c4cg+
kFSRVK7wt2s7PKBrmvGhY/yiw/84f8P8IbNEWOVDKEedBLseD/tyzu0UogquYiXf
saXO/oFXAYd+j5NARWUT9GXi5NKb0pxBOC08mx/gfepju9xha2ElCZHkXLCoTjO8
pH8vhVxGbWgvpQubY0BGFC5mhohmPrY0a55m+JlSLDaGjYTdRcZS1eWDLA42Dm9L
vI1e43sCypUiubhks7BjGA2OmuBZF8SFMH4gBqEG2YwkoHk28xdoHca2qS3U+myd
RXKd41SthOj/Q/ZtInA52M2bYZ61j+wuSruljsX5l/EVmlmcCd8Haw0CQyaj1N+/
/NZdZgZGv4QO4OIoD++CnIhkM7ajfO5CjLfRS+ckCzJMpzzrllozmOgERTuHn5xy
TSFEGefMKyFRF66uarN2sRbSeZlU2Tvbk6/ZKH2mNpjkbR5wsl1EOJgkpCb8+RMK
xtDbMFWbd6o5HvNAWIs3TDgozbB12hgvV4P2l0zwVjdBYYTfTRxAHCsGSXdan9/D
kLtAGHBmuA1QxNTImnczdQ3TioYGyJ0AIow007badzSizAIkEX3NIt6+Q/vuIixM
O8WHWEDAcP3y8LmwE2y7PktyBRjEBWIo9WvaG5PY0knQSuo6Qn6fiIhZNYCmQJon
WJdwTvF/JN/PYTHEZiy7PfY3IGGFZmm3ojpE8yl3aeK+qiVjgmxx7IJTZ+IsX1Jn
dd+j2j83TszowgxlAXf0Ee8+kTYGvKULw3xDgt0Ruy6IEbglGGEIzX4QKeDZ74qm
gz5JgWT8PBfM1QmQtqZzYXPjSXuhPiSh8+yyJKA8j/afqtHSQLdB8Gvlsy6Ce6Cm
jUlDAOyNZTsbok35+vLH1HoX/OmS173JwE1DtCExCxm+wS3UWavcs4itKEoeeKmE
5fFXJenLop4k5Wvh7OIOljNeYe3bL6zFWFtTY80T2X+Ww+vZd3YbLaka95vBv4NN
+rbpBGwY5RCBCDIXAlya7Gb0ZwRyGBIUrtrkPERDr05alBSIMhdFp70DKg7gkScm
IsFOdaSQFScGx+ycsERt5vocJM/IBcIUvxaQv5xJ9G8lDrIGuZ6Un/QvaS0Bg11r
nISm2W+Fgoma/HFs4OqFGXeDwHVTb1VpDjuMGaqAkfCekhxYML9dItPrfSGIxEti
aP+0ub5DtZ/jkfsC9o8bLO2mHs/YGel/w1enw6bAOQ/bkCT+2PKNaOzlk3JuXqAR
pb7k5Ry0To/6a4vOR+pXa/tpHVAB9nrvcxrbtTmjVRpMF350g07ufDHwZiDV2cLc
QZYKyoQ33e2LGIPc1DCD2U7r7f1ZmiJDuPQwLFPFX4jeRZcq2A3vblA0zr7XKgGj
qdMtnbn1TczD0ucXXMC1DvIJvJjA6DcEHzTSwOQ+9nFDN9DCNa9NkOeNuYZelUB7
jiSH6iMsZ12LZ4e48FLGB3AZpjngf5ELr5LogZPc6py8uhoE8K5wRu0E2e7ceN1C
VWw2zVQxIju02Qv12Im87zRyR3MknbQt6wyo4VkVaFCQbNbl7KmFK/AsF3ccalX8
Evr4YQzbrTm3mr07higFFKxmIEw39cV3RxZgT88i+8tr924av4sHYDNCuEF7a+Gk
K0ZTHum/F/0h2dNDy3mEpyzWPXA8aXqdx7iwXh2gryw8wmBbouHF5r8Obx+gxEwz
7XQq8klJdG5cFJzlD13P0G94AZejJfClHUXEbCQhDnOwT/Lt5jv+S6pt/Pa6vWxT
4Bfb7kZx3A0k1ZyPdg+R+iQwpi70YuvF29j1NLdHUdeEuANbtHjA1g/YCeRwUmqE
wgPXq5dtE93aa7Vh7rI+gf8Nw7xaVcw+JNlzeuCdFkrNhOcCc65CqRleJqKV9tU7
9y4OIC3GAKFdXotLFu0BIx8SpPLSC+mB3SKuqQJIx3/7Tb6+sCtipYyYb2homioX
qOj8VEoL6tNeL2jdN5MSM3gUgZCLC8k/BCo4yQu5FLrfdpNr3kfyUrYhXZn4czAR
B8StKtKo1ZAhp7dlk2zvyiRs0QKNvUo1tihCsgDQL0rE4zFXW6DOUVZTHEvBg1uv
HJAsFFqVFjXrk1lyGn4iqQDB7XriLB4/gSG92gG6jycV5sdzbm1TqTc52Euwa4A7
2goqesumidYWo/exXJV4ENmPM73pnwDtD5JLVB8fCLHRL+FVHI30f8gbRVP8pjEm
Yl5Qc1X0y76zappzcncAkWx3/Uai/SAN7318avvLOKNeevO79CWJFUXxSQD/qz8n
yAHv3Hy2Rhrg1fq537+dP2kE8ek3HF12R/nT/yKnxMEr9hMSc6i0BZ4mmJBSqsS8
CrIUoVCUvxBUn6S8NtFVmzPN3m4T3akiuCqf4X3ePxVGXEdc4TURoiaKclThxgMT
/tO0hovQzwJhs0Us7/bPWd6N/ftCm0UWnOtrjtwgqFM0u+Y/B44OmRnEpiqBxPvK
gJ9+eugl0LHj2sPHeyVK6zwJMi0TMYtrYcmiM5QCjsLyrANhj0fghVIm2x/vS/xO
3LyLqWTZXHqESezhanNezgxj6W4l59AvB2i0CFTy1hCuACIkAnuo+ARPpFzrY6Wb
7E5GnFSBAtGdcYBHOagNNUFe+YFnzsFcYhN9mW1olJF+tiyh8nU6cmPlEPXL92IB
Ct7lc1+TvWj7wC7M+JftW6aOvFj0Jcm72Vc6z3il2fShy1mlUZF4dEaSQjA6cn+U
aGg6sP+yaQpDxHQIJkS1mxVu+PH9eolG6ITjWVsqto/2IEFHmlmPYRn2sSGSFz+w
55Ze8A3t4p35y+9zWMAZHn/lTuhXgjT6FcgDcW31koesVFVwmjjK9NNcmbjJtixi
T/lT6VI7ErmDibBY8AB73XrZCmyKrOf3tjLA1ka10IXahe9Gj8LNfvHMbngm4r7P
y053/tMGlPYnxEzbpT7+nCmj0YSbcMfoLzWOyySZyxOiegkT7P2DZqNIHuYQ+hbR
S36G6ahTIZs88PSqd0dH1DTfcKLsT4XM1CTODkVbHb0N1ZnucB8brq6LDfvmmsqr
di3Hw67xWRquSiqCsGITElqKJZ4Ncm3dGpqMz3CObk08opm39GLToFuPBQdkw19U
uXcbWJFryxfqhbynhNoqJVqbJcS4Mg+LU1m7pU5UyRmZrEUAVHVNyuWKJjT+D/+L
WFbsF/VZFZkw6iWcRI4sj8XyvMwkiHxB3qdAIzSa/NisiuzfqpySUymR0lsUGO0b
2rnU/8mg0Q11mnjBIUtJ5Um126XwoidCtsGxLUzxsfXhM4EvDNqtQL2kvwqovXe0
NHBYFIHwqsOTQiL7+G/Y/Dps+ugFDuzfGjGmEP2p75UsVKqL40DIdXmPxzDYDkg8
THlyYbaWQ5NjYVDZew+fOmBIJM8Adw+SQp4D2TiYFk8F4c3xbevQJ+o+KQ/QRPxD
q/z5lZENVMZ3SsXUuiQI2LyhPn9I64XjnYR3dVx9rt/pY9Jn90+GszAWZcIyi4Sa
qDVKW+Q0Q/fxBn/W7CUawiC9VhZ1mvtqE8zLEqHNqlgaxf0CZfPcExt1ZeM+YYae
hzcgDL814YYJvgmqgWWN1Gh1XkQp6Br5f83b4Rzzl/SdU9QWRE0pZUsd6z2GL6O7
LrgAbdp70DFAgheAuOxJFge868+8B/rGlc/qzAwpyqkvOGHq+17hGOkXSQU8qHKy
rd5v76XovcT8TrCIE4RAxqJSDPI8kLtDzz2NdUBnxuB5mx1qqEhAmN/dTNq92+Q4
dRZ9eSKnb8h9x5u1MTHR7V6rIT1MYXpcYfhZkbMxoYazqEZS6/4HHWSlkdGdNFGh
tiewUE/eMdYMUUypTZtIuWui6IyTw/iuz4iAt1Hq2E89q1xgof+TFEyqt3PDW2R9
uPqygutqU0ZV1nE+3RKSx2ydUkUCaDvloWYhTJ5Y+nzY+n4UMt+fOoErLoMZ1Q15
UQ98gojasYzObRMqQ/MI12RZVVCPueXECy2SyZ0fJ/wwyolUF7s7DKcYSIXsBvR5
BKiL8yX7OrV07VUxYdno3TogqzbEQy2zYA4Unb7RgppwGnmJA2yB5+1wWG4rOc2s
jIa6ZAfdE5S57w5wcTuHzhWoIX5IFu3s2Zyd0IAO1TK0tZlx/63uztSrfOGj4Wq1
+2gyPq5EcR4Rb+qL2NLGFFcCoFki0zvThjcKTjfKF2xV728JXexwrxtFQlVIkx2a
2h0zINwTAu6on2NZanfL9mS783f7FqHMdWBTAtuqcOB44VFvtn2Yzqn3vOgrE3ZW
mRJo4XpxVe8jKfaVtMK/wQw7IVsBUbHpoThYpdSINcLSeKqTVZp1iFjLEdGOfoAH
lV4JaxK2OUVg09pcsziVxs7MWPsKznwuavYN0CpYdPdK/Tl7Y5mOMHHX0O59vPfP
w3bsRc5OAhzxEkcLgcUXDxnhqKayE5k18TfTOGj5WA9VjEXkdejLimnnjKhw8Mi+
nM79UbnGG9FNqiptndT10MgiQJ/TZcizY2IAhz3hZTU/trAencAoLAmBoZyVNdlb
I2H1o5xFMmMuSEfbz/hK7cunD4Tbyb7XvzpwTJnvJsI6jT39Pnc4PYG2pfjLtdGc
vQaN1ucrzrbb0azye8HsIlDBc2TfLVbJsXDeKRJAco3Z2VIsEB0O73Oy52tCD33h
Wb9oqtc5CnLXDwyk/3V+JYnkQbXgnpc8uZTJuRrXOOFo+4wI9McsT6b+VX9/RV/0
ue6mkEorG3i2apFU7OnbIhmP6zx72znRFCqp7VkHzo2uROuAXsH6oZkxdf3dQ7fv
EdUCLi4sxdVCj1e4WdTnCqK20D/oe9X/CCtLPn3BHZR+eNAP8yaRH5GPeouJOlwL
d47iuvwYDCnZwYkzmy3kEXg9Lre50eagQpxflZMXoGbCMFx372poLIAT3L8krX/q
cfvmYLVNyA0GHMaDvFtjsQBqUVtI0WC2zZ1WwPZpDpHx3ED/eeDi1FOSwOeE04Yr
6/IYLNefwK59UahjsQoYqJo+4PRiCVHT2cBMjEzI2ZmIJ7KpY6i81vNQfPOnbM90
Bot/Aa3xY3F8Zyci+mvW1rxSjMWEXjHszaFkB+1kqeEWMQGascu7fQEho9Em1aeW
FC7yKuf8o5ktQGtjvYMUlqB+yJQlbvGoPXRJ4xfj5mn7U8nuYiV0H5xZxTG0DBS7
gWRd+znMgS/03ezVrCfmun82G3L5aJKEqcMu9yz6w6lFP71XutIjaf7DkUeivkD7
8TaMbixb0szFnpZF7ET0Pr2foT9ATKBEOU8JWZgapljcX63ScUKcWE9F1oALTDJF
OebS2iW88sfdaTEy9lxWZQJ+UX2M/vdHvBHTPwqhs70kFf0xAM5TPES/o/08zAID
GZL58UQfHtI+JtvZ7l/zfeKBZZqBZDgmnMcLH9yB1C9SLWNwj5kc6n+MkfDVo9S8
rT71dIGaH++2uPQ5iAHt/rISZBpNELgdEHujgApm4Pxny6hbp/2mxuWzF2tgWGJm
Sl/a8KcVpwlHc0Tky12V+u9m2ZAc1eHFmF7sS/UCkp0ridhuZWFoMsgu2MhqinGt
5B6UgT3FxHAEnT7UbV21c8zoQxI9s6T4GaMgS+2g157hd3Alo+7Zv5nAfbL4UEEx
ZI/J4NNah7Oh/LZJIFGV9AsTWeYX2l3L/ZoKQbdPmFOJVck0ekMnGRIfcO8aarJ8
ZujuaopeA4waQUh4dkh9YWo14KsrTi6b+DOKegmb8W+wvjdptOC9IlD/ffQ+jUgT
qAUhfzYFDL6BsheHBXFU3fWZYd9RzNj/cVtHSfqESUBmS4ob5JiUMTGioEboGxtq
mNqOO91aQkwgRl5R2bFrkmiNS3Suqy2qI7Q9OqJuIfy7R5kl5Wn911409tm7KYAT
PUwE2N6HLQsCYvfgLGP/ewm/pvACq0DDsq6c6ag3HkW/vFsedyMyvu2/5dDca+Mq
3QWwGBmzKmuHPqwg67QYzjAm1a2IuL9JY+S9CXWhd7YG7A4+GEu+QHWG8Et+gXIe
FJ/qEzW8EIdX9avWHViiYbFSLptaOvaXgQr/OehAnNr77lMlzQv+aqyq8NUNoThz
LfOOKe06BgdjGdtNOilPbGOlWymfz6xz8XAEI66uPZdRN1APkN0JJYOfQEXtS8Ez
f/ikr6vVKvKJLbtnroU/HsrAKVhphl4hm6kWokcUNsw3mIujqdqlA+NIugucKFPY
CNBS+KipPK33Ttz5uHhBvMrkv0u3dojQIORCOylv/tO2Po8+LHJkDIPr4G/vZ5dW
ExHNMpRCr0gE3LH7LPyIGEbMRgRgEn7yfLmCSHdFfyAoGykoT7gatoPoMSyJ9v52
N5vxNsNqx9+GVc+r16OcinrL2200piWV6ZDF5DfiAWvp96Ejeql+ZuuClb/v5PVA
S+8tWNwpwUX3yimm123f7jzALRkP4MItI77l3qBC+75s4uOL+vQ67sK+4CeCYnCG
t3EH9Sz5d14K4tGFRocNx9NCj9l3H60oA6cNvMWAdCUbJGnUYDG46KUNp75WFtZ0
UksOlhcIeRtFqSBuqx4HxDQJjMHdXSL0R3i9jGDm0bMPCvC8zj57Z0PxFQMQRrj/
cVdnleTb0fIAJKCWbfUH+VmRiz3yyZF1xL+QjaNjlbAHM2GqTOaPlsrX/mj1OAB2
InBmAP2CLovPDSrc9A0SncjJvg3D49lzoTqRUnNfM/2Tkem7crESx4AEFk/gnWC1
2PwcX1sfgE/j85XqJfLBGdJo3I5oOROLQ1OJyTCaXA3vM7oc+JZLdzchVBm97Hhb
ppLPMC7zWW2yqmNj9KrcTiTpQJh/bd2ZcZdSu5uWOAsSqYFCjRd7VnV2IGySkLls
oS5gJvOPutzrSC0P+LwE0tGFHG2tjgMJPw+M48MLe7/dcGFQnRQJlvsg8XglCqu3
CIEIK2StfT42D2CnYC9qVRxobvkB57YKqbaUxjW/5mZKsQSySsqR4lgnRXLbT5vS
D60KQ532CZECE2gL4XMIuWQ4c++o0H3fIjNmEcoV1thlZUxkWCMkYFqOjvbhR6FL
5ra/B7sQtKxsmi/Ewk7uR/KlSzTlnTBGgBikbgUWAHNyeRKokKw0T2HcP1nbUyWU
Qdfkbj7nviBuXmzV99SrAhdCiDPWavXWG3QNNerYLUx7AAAkNXPIjlrZvJM1pVKi
ZJCD5Dcy/15aOFQ+xvokSpFOLHETWCO2M+yaG0+676NmNxlkwDc4E880WvWFo5ux
iL9ujvArbtjsIRpDHkORKAXKerDPhrptmRRwbaRRc8RTqu4HScsLBAJt6C+Qc2Hp
ERc1q6f0cTLsHGSm04QEDp8INoCs1vReledy94vM7lt//ROTUf6cYxTQDMo7/Ou2
NWHsfojwP8WaOY3wpp00J2vXzqcw6p410x84+LlNaFXEzyCpn33TnmpOo9bKpfcl
hixLb1TW8qv1YmdjJcxGSakFiyFVlZO6zd/Xk8YfaQ4/FZO1H8QJxaSZhg4fQN7w
SGm8DQc0RSvoNwWsJrODsclSkOdqVhXZcYbA5tRSvqvRq740h3q0PWmdoenz7sXN
xZLovHdfQhCsEWEXJA2+af960BMSlRqjCz/9UC9j6NNF8/RQVNFB14fbrLjAfdt8
oRCp5QOKGmtcaJOVkmW0wTlwIcFviYAB/1XR1vbHTtYX0dewNFJ05WIcSoRhqQxJ
5ZCXfiglQ7cOj2elDYu7TltD4Hazj6ahqRv3/x6v4Oy0Q58lIKpdoSr4XZ5r3Ico
V7FfT58LFt0Oc9ySKL30tOSFdMkOQ4+wX1aEnqpfbOdfvZBiC0lb7h3q0N7BFPgD
Ubd9yyBmCPDMtn5d4lzdDgdLsdMHkzl7wQJr7OZXTb+3WrN/mAJn2jpH87F1JzBU
1NjSE6NGcaA6POcX3LT4WT5J7kww0AUM15CyWQx3aVuKqxsz843LocmStfx5ZslF
8iuLC1Yr0wYls2xq1Ke2773z4AaW7daySrEyf7kvySaQrqyL38+OMcZTeicn+zw2
oxeFG9/Hwo8LOMtDO7r1VpvNbB/4QEsBmlO9ofX/Fn226eW2hW6jhkPgHpb3pGSo
8eTGpLzXAONWacjk5eBI0fCEYTzos2yyVm6SeiSOb2xgBjRJQgGDK/TJihJvnUMx
8AW9kNR2pGorIH71iYg1cWBMLFqAgkgRq3PvNIkTpM4OqG2Frd4R6Yha1RdyLwdg
CXeiZjYcZyl65LA1VM01p7xW1G4gWqSaG9/A8BctIuiS9EnbK6CWE22tgSob2Gsl
nlF1K55EXUx2LPlEihT9hU+doU4EKjAAtSfJE40N3y+as9AIc1G8yOB2NUSZ1JTJ
hcDdZG6SC2W1I+2kLI4Ox3wWCGna77IRqlgeulsVMwekD9woVVgsmyydAloiFzfG
7M8s3+fZFOn22tJzR49ogxKtkF8/QUaENAJM3huiv9pKdipUh0qTpeSjIwYG/s49
PHqho+lBSXXfXyvKE1F525i+DW8PJjQKfNGpNBr4aJusgdFQ2MRz9cNq8goqKfkx
/TQnySKe9oQyANtODLk6TsftwViwcGu5a1eXJOv+mQ02q0jNLkRKBaIMWbv7FPsN
0ws7G+Ne9VZGozd3g1UpqUoqgH8UkO7hANyNp3a6JdJMZlV4JH9MnAD+Wa3SE9QT
gQlcBmhtTHBAjGK6UaQwzkt6fLc9PM/SFtO8E552t9wUBMDwopPcvk3W3V4IRCgs
sT7tL9d3OKgIlo/32M4qbRGxb6+B8jOsqigXoj9HRm+kq9RhRzQDXmmep6YfC0j8
DVY661YEaicpCBjZkZtOensPVyRDWrSQRBugJrQz8KZ44dCKU2fsUTk35WgkZuMO
/+ju9gDRb5AfxDHjDPVmjNeGlwsGr574XBHMDlZu1QJINfbva/5/NHBbViT4tzx7
G5imjU0P/MPBrIQ/NiQafDVmKS3Fd6O7NdvooFNd6yICyYd+2X9qaJZCtATQ9rIj
53yntNAsB5YnmHwjf47nRG+5nug1DFCvPN/M/wqlBSjf7/kRgIy2lPEFI0vLQNQ9
qlTnGsTA/hVqdGlAZR0GrSDGS90hmZZAa0styRJZ8fvPxNbIHvjJ7Z4dfnRlWlSd
IwBXLasI8bb8b/bEsEUCw9np3NQuVzhET2piu9Mt7FCI+OQ2uzI9DUk0mp5T4Muc
LlBrQGNftnBOT5Hj1/TH0+1DsC/COoA3yYZ83F8eTlwJUUPDD3Hr7q1oODMpAj/C
i1oZlYI69E+Sh0ptq6I6cUyV+mwttvS4+5nQ++eIbiIaB+RTpdnFyuba3zXs5Bd+
jjns7j3uPXHc46OWZLbFrsgD8IRygeQoVhNr9GIZXD1VV0PyBS3hnfEX78u6QFQK
+gbA3brwpupVceJ+yVzMEv1Pr76L/Hz91Gg3H/nlIxd/0Si4lvbrF+DTLbuWvKzf
AErqYxpY0Y1hUbVftDw4nTom5GY9otcIjTrfcYxZL+x//nTCya/BzEnqGGaglhIL
TSoNuyQGT4FrNHmWkLjK6QQKN3THZocUSWJrrCt8Hsu2BupbAnFo2FjTkUHeaukI
EGxdELF8EaOBatiqlI/tZbZcmid0EEbTadKFl9WQUlWrGeSuLppB696LKLjaK6zB
Rct8aJ6UiAmTmUJWIDEUog50STlQfoapHic/4y+/xgKuU++4YvwmgZ3kpsy/y36K
5PV5uT3gSgb7QZnpdAzm2y+8GAfqux+pYWLmE1GXmV8xR2FT0SaUIERE62HUpk6Y
jkA2Fko5aes+sanKasQWn30GM2kTZiNFwb0uuw7NFkA=
`protect END_PROTECTED
