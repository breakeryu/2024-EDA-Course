`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYq7GWc5bs3DLax5Q0bJPPiig64gWYnoIPPxin8A2JdEIB55FY3Pg1JVa2nxKvE6
kL8S2UsX6Rs9/X4m8N1QkwK4So0NjI7JqfDi/17LGqDZFgsHMnplG1QtdYIyQXOJ
uCryxO18dMqjv5QQ92Bx+HAGIPi5XSIr21Ybg2smFfBzHnOKNHKmtbw9SM3jJjHl
NRYcbSBuINdFZuFgMX3AEN+/cnBbLulIkQoCI+0AYRs4IRsh0RKTsx1nYJj0yT6t
1SXexRXAlPEkldPx8DGeXi+cd+fNIFlzLE6CZ5/fn0180RCVJI4CnWiYfKBv9e71
G5wlFeO0FHzfWG8mP5ZWZZNcm9ZcPmJJB7YMEzwHH6rh+7/piTM3boQONudsUyqr
N+DPlPxy5DHfkXSgP8RiBmxxmIj7PoH9gBZMHvvXGh9EzYsOUPyzxcKrgZUS3gJF
qeDZHLsox9HfixEZvEJ7Hj7rm2M9SPUW5P56+VL+4VMRLwnyTbe3721evZYHJttC
GMucQhcKwEA1LAVDjgJxSRI1jJyLRvf3dW+j3LgyHVyT90f59xSy/Agua8L4HCuQ
kwuUwrjgN8hAsi3ci1NAcRqVP2EZPRsUx5MC7mbXWn6AAlsd9hUQwk5lCg1F5Jtf
XUBh3qKR5haXYSI4FYr3uNjFsvRN0Z3BrPavBkraGDElqjdsQIkASNjxiHOwQ51M
WIk8nDmQLdqSbAhiHTg2R8iBurWPVJXvZ9oA0XkORRyLBiq0WsdwNZukygjqgOQL
5r6qv8k/X3JKY/cAY4xo9GTIftHVGbyVHsabj4ndgrrmg1fMhmR+v1xIjCRL+w+Z
VKWG6enTu9PUVB7uqz1VOdDwwR+o/CcqxtuYVI/OUuVp1S/Ffq/pwxB/uKr62aOT
4NL2RqkOFgTQN5NxHg+rk53762Fx/DwblCYVI7STxj4sRyv/m1WtYaehQ6Uy5Wdv
MPhv9MSZUA2E8WWenx6M9bp4dr41GuKO4/tQdnq5/pJOfc4vKzv1pYxsYyM8iOKO
Q9u+x+UEyVsQjLO3xcfU2q0dvdAuPkSBYD9LRSqHNDHEmn/xwEgOvyx92Q29jaUo
7tm3VCbYGiU4rwa3d00/NXJScIlMPICmWhMtp6YEmysPUn48d+z0xSi0Hag5mlyn
vfd7jFGtHLDvS6a+eyR6CG+XYZE60U8+EXFH8gJs7W48OPHXllxWre7v1v6L8GBO
TFx7o3fGD/8ArVVz02HxXpj+lA7wVBlf0DwVHUEyMyU9jnv3kFBlbjVPlLLVINe6
+LtRgrUpk3ykIacFFSPXgaK5QUHA3YBtb3CaO7qMJKo5EplX6UUaVTjm1oQiVPS0
M3qy79ElSbMZbmzz5DYrsTOlowI3QTObm2jIY3MDOdne3cmePJ6ZcKStFKTGQMNb
to7FIB2WcW9MVw3cUEN+IfrNGbP9qGoKQKJMpntWBbphPnZXlIOuqhuL0ns5xfA6
027hQ3cHiVff9t5q01xr1Ac5J7zOf9UNRI7pGszeuxc+Ju62CXg6nf5x700I4gCS
I4YGJ+2jUBImFo5MEr1TlFUmoNyAVsghDchkxZXR36L4NYEQG+rDxvIto2JX0aVJ
8Ankrqchw6SBKuJCryP6dR5y0mt0I/8MBTxpeMCpLEn7RXojYcguA17oR08dNsXG
RuWdmbsW5QYX1dxNseUJZF5TX/+aSxNZiaSydVT7GEZVlAYaQZJ7afgF8qCDjTGt
pA6kGeI39A6QuL8+poyARkz5zaCkMC0dTqw4P78UXAZNNvdCB5RmQ2MTbsup6d//
IY2Ejgj3u0n5w04a1CE9V3tm4gDk1d4PtvpoUHQaEO6ZDqcXnvSzV809U7S2RBG5
ftwBDe0TLMM8Bj/z+PIRpFHYViGzl7UODZvb7FRlDnk6Vlep1X2qOlTF7C8iP3tc
epjCweRLGq0ZlpzGFH1xXa8H2xAvl0DsMfhcUEoYx78Lqq4aKzHr8SMeg6FDHqzX
wE9Dqyrvzca7R8N1gljpWS5pjObT26WwDgh0KMCIG9NBHHHKzET1lOZiy4S73T8y
9Rnmh1Jg0RLyYnmeTjbPs17q9eqnM+rUg/COsnZdvFZQnkV/0igTqBfm/xBoj+zZ
f0ce9ii+fQPbkmtSTqklK90j57Y0ZIH8HuMWgzWW6oxzUmZdHdJ8koXYY6EUi6Mc
rPMp8pt1HPx1q4+bKUkBrTZJbvx7j39wETtK3sS91/itUv2m1I4MKlSHS5WMwwaI
72Jty/6H0inqK5mGPTrKjwG50U0qf+KyeWe+qTgJJxgVWnUhKdWJ2tUSe6GoRtkh
l2wQeMo5QUGdVAjoNJm+VXQy3+UaI6rNafQIOgqZa2ovUq5wwgElJiLdX0VWExUH
NnX8myoiIRijDSxuSswRYNTMGTVyIqZsgXSWdUrR/G1nE6YpV3E4XzySRuIju+gV
vD/RUcU44C+Qsyvp7d5DGg9b3AllmkdvViZwpp9mtCo2+fcngBW1lqfnHkX2++O3
XyTicnnWT2TmP4WoDHxw3rOnPrcPo0bPcYwp5HQNoFMhxvABuu/qOibYnFeUqME7
GSTWpWM5rIwlED9zE+I1hDFfSCNyr97FF/5ndBBbm+8cddmNaK9/w1Msybei7P0D
+nJRd9K+cUFwj19r8IYUnUHtDG/SGDzW8O0pHt1ScQRnsJa4EejU7rvLdm8qPnZN
RA+jKkV5Q/zEo6BguA7RN7HRIfz2LHuSKRDmKI7PLQfkJ6MmBh/BgRj3MYPrK2dk
YqLi4yQ+OXcpyCTJif+c4I6L8As9RikRkIM5LHvtuOOCWAPC9IZyJGGigx3Zzvd+
lc+aOu45JyloLwPc05A/tjoo6tJQ5ncBxp0WRnxaiu+zMCynST08Rmr1fwBmLPQH
nwa8ZpoOizSbzyK1GihXxPvoUqpwaR/L56X/eGUOgjekYfpOs7PIuAJhRv9AlPor
kbmLsqcwxsXQfR1tiGpnx2Y+yMVq+/p8J8YMQnyq2C5iFtxxLzZYb+BM+o7UZKpy
kQlISxk/AHbivtPKYeefjDA+6Df+YaFGPGmDm8x6CyELbeCg7/oz7VNEfec7zqFw
9hzMSDmQPzK+ljOUXReuBS7+gnrSGqm3HkTf/Qk7rr+1nQMSyZ1ATF6/hTKLVGJl
cRRmqmyNu1MFoa4NttSGaHrYb3awjXPszbJfMuZuvtvRHnLdZStLi/ilizjdNW4R
u9pIe90uRtDaixulLJRIOLvPfDzsHx5scTr3H1ioOcvmpS0tWdqxvqG65A4mPaWS
ZD6COf5SFrWRqEJ3LO/RHveWr9wQMWqdmbSA2rL0yIdUtp2tMmF2Qel/UKz2fqOj
8EOTm1oZetwsyIFc4kg/dD/uHRwMB3Pa0xpmC8831JHXckzcFSKdT7vG3dod+Uj5
Dyk47254sB/fZw+CTIKqM+d6VCVHJ0EEF4vlYexxf4lQaPxtjPir34ZOzvvvlr6K
zHL/Ie0gR0VID2BByPIRyw/Zj16eO2vyXpt295UnDzv7WLN61ZW3u+vfyajMrUmI
6QFoqnJKa/SMENBclgqP9knvixUOBOg9TA7PY/k4C/RMN3rIAboO2mzl8SvNYZz6
meUTpNF8jnEi+TttV2hF+btb3QB2HjxOzDmxmIvp46ob1g40PIzlhnAqSrLvwiZd
asPT6kpiokzHgHOywbLugQGGBzD76F0FqkzKCMEnmhcPambUOPGmtGGZjH0iI15V
PGN3YR/fONeKzi+cZBHxrD+bph94ucfCwLK+6sQIbatJaNxiQELrlLu302kKMfkr
ySK9J2/hOxpvtW5lmhj+GPJPvVhNv02alxwSWax3XHAEiBfylhK0shs/YGSelSFn
A3vV4iuSNQI4s763veQigG27sALgGC9FMsU0YEeg+NsL+xu5z4XikegGp3TEyVcU
IGPFjmezSJSCWjyfFrgV3398qh63wVpMzqTvCRyCB+Nshmjh6rjQw9c1wRgLKEuT
c70O67JOnfl7MzQS720DkxOZsqBeqdVY8sySI3vQpRQJijBxR/BkOYwLxyRDX5q4
wZ6Lz6urH0/zizd9vPUVFW+XeHGueUcGqu4MvBcOlgz33hqYthXRrjicfwGgI3an
25O/bhtHAYWZegoFnOgs7oIGXKBm/Z0EAqngrCqV7nW2J98AacKRn3Ho9sbKWMPM
7n0opEaCoLHLcSgDiinlobQiX7U1l2czIaJbJHL6bSFR+7NVgjElig0KNGiTZ7Ut
0bFbYhzp8ZiSBH22hK3ff4U7d4of2o/vNnwSAXloBEimb5tMoMCN5NC9I+QurdjM
B1hVBX1vK9Pfn5GFNMd1FLQG4ZQObZi9RsAn0xIg+XJO92na4nPjoNfwaWXqRmiE
b6fpW5iRsWXMQp/Zykt+0Pnl0fXu1NhTq/vNKjnNeoy+bm3PB0/QcfZcRO9Fo8/m
61TP1uuOM9utfBMvL9+EqNORi+//5kPRsyIVLzT16yYKrQENaSCyHedrN7GcONpU
GYZ0kyyWR/pNCo2PLVc7rwpU8TLnsPOII8oInosNoRL7jvrvneqi6QirT9FHBqOl
aSlGv33gizLLipeLjPC45SOZ3erFr8T3TtEixs4cRBrzTth/ObCA/zxe2uRlt2SS
E46Eyh8v6MD24+LJMjNX6BHElWc04aajDVOjw0ZzA8YeDkgkmMeonBQdMzkpGxkV
iWHMRjb/yJy3adToX1kP7EzjhY5uwQVt5DqYLYOUP1aN8+3MhCXy1U9zFbFBVULW
MZ5NBY+0I5rWcBfALW+e2zpIlahX+USoOi7NyNyRz5JddQL85mQ0y1siWnhs3/JP
Bv1ZRWIBJOHId6MYhcway6TAJ18xl8XTdVUqbo6yIbcjj/dM4Z38crNSin7pPQya
RZWhMdhsD+ohnIMy3ELyYVmYg3RdHLmDdcH1rbXzL0Xd35u08L6VPTerdUZNCevf
Ug4OHWlPGwPLMaXXfI2j8ElydDxqBhOnZta4OaIhFtfZEc25ndqYf2p7jFMNvXcs
NjlcdE5rcC9D1GKvkUU8tRMcG7XZ0RObict/Dhp+WSmscLHZoFQ+dDseYUiPJ0XL
FvjaFfmYQKMCliciFEC0NhfV/3usiqM2RAXRa3OWd3/Jkl5h77gibgI9tNDgzVkf
56iQl7qBRYmamyG5c/JZIiyzS4tCTV9PTb1sVZV+A8FsqalKWAzNK30kSMCyOTKx
zpsYItyBZuh4xctSe9NwgVCRic2v9UIR7QgpS16dSOYGNpk+kT14kkZdFhGONMkG
kX2LcShN6SnZrKFnR+zhWU6f7BBeDnCnH+HjKy7Tq+yHskLy9AOmagY6UY1vpAQ0
3AJy5jmZqHGOjaYV0T4cWwbRZtiPoiNXko4N158C8HyBlBhk3Z69gte/9NZ+sRk0
MIc5xQULRH/wJJtOHY0dhhS08i1M1zt2HeQe8OU9/bPZBWi/ok1nSlICRg9P8saE
yWv3bTe7ob+nfEr5N/VutGwbAvKzdAOoI6TDn7wnG82fPwKUrLs4Zrfcthqrnema
gZSrVBNxQfMAC/kCp48eWT+9WoEhP/UmFUQiOCAO1OEuyv/LrH60Ca72fnjrfm5K
LFLbsQOPqKHu3SZeCC2Q5N7Ioa/uLYLZhUGbWP/Hw6OxyaFpfuGh5OjRFCphInkN
tiWXPeQ22TklIgPmBIlxYE6iGjVnadI7cwzEkU4R+nQUFtKhGtvvbF3SSHDS8q7R
fqjXIND5v5kSH5r+jGfoOlMyBzk+yLAGndaP5G+AgeNpjiadYKLmKwh6TjZAKlJj
5x3pBz7Hc12lZvRpI58KLFJ0Jmwpvrg65uBzRg+e7uPFHhMsols3C5NZpwrCQlyd
ZV6UmcMusA/X/iy3taP31zmwnvCPcLgXM6i+Ma06wuRtCLO8R1Z0DYHc4YjdTsHD
Lb1HHLGaFOEsS7JIcmvwmC9Rq8rJQFCkbbKClAIfYwy9h8kfPlWhHmabrexFeBTP
JqHhDUbG45v1FRb2HNa0qjM70PmRSQCws46qtP5++aQkphhbweWa7Bo0TWYbMnCQ
nLpTmTg6K1Na+vtZedzzGf0C2ML0q0iOkp0DoOIIDVDGegY68NdRlbm1hYaIKbWh
jFXb7ornwdZjx7MAcTH352Lu1u9mCmla2NS4Ub+RSw32FtKo9CK9WQw6UUx0FtlR
mXn1bjiKoOtxYi9I+26dv2LPTHozCORyN9hk/N3TjP0dHprfybZNP5lJUIysC8tA
ZJPp3AmubDoQgZkANyvoqTgVfXjvXzgAW4RhXmlsl1hn3741BOczFygJZc06vebu
9AtPZ4SF3a6hJ2fJQDdlywv71SqUJlHBkiUEtZYfVLPyHTdvz4LsuQx01D/KyU8w
JKlFs7Q9CyR/QsbwP+9H239HTLKIj7lu0+Y+TqfXIt0e5t9+8W8y7rkz5r7kvrf2
Dib3rNPoNx6CAgYr+1GkbGoQ07rXW5oa7vA1jIBp2yNY37/I34XKMRdtJufYPzpf
y2Wxa/mDK1DcZPf2zf/+/yTrppL2WLh6iZ7PhyD7icMCB/aaoEQ7DX22ZyT+dKvH
IHZa8ib3vsOONWCQaz3K3yg4ny9WwtWriq29QXnMF2sbTcuExwtF5LEleM1DtrL2
vTAVpZcldhDSp9F1FO32RyVFv4nND3TNR+iUnQkDHJVWEQvM298iSlf3VeNsogsa
SF5N3376mUjbTUR/5VMeCwvO18HjZuXpwLG7+DgOHqgLtuiIAjsrqwE02eYaLpXd
PVfs9eUa2DCSKGCrNZzfq7xPHuRzOVEYObCX2VbQ9Q5UEJ0BxbISLCPPdKwxkedN
BRY0YlIgEPJhra5hqz2yBpVWX2Jqw8v07psiHIWasu3JI7pidp6M3Ud/domlumWJ
kX1Nzz6NJ5XAjeg3AXhm8MZ1sPdSsRvOFIum7LYe17q9Rh47Glt2CQYhlrNjlZDG
knNHFwUC0kFzoJuxrQ5kP24QznF8G2G6GOFrXaRgyq64Zyh09B8YK1Wqe1S32D6P
a9JxyY4/5F7KGCr4fmmabdAcJvsQ2FFjS7b3ae3Kp9tBqQ45j7lJ4xkUME2eh6BQ
cFM78LTHi8cqaQLONQfVHLWr1jNV6KoBbcE280qKrePSf6aZr2ZXMQsWzSr5A2nG
aFP+FEB7e1mPEmqwswTDvhczJKKU63mnAXDB/V3erKiJhp3MKKJQ66zjhikr7Tnx
0dR45HBLc4r3HjqNfwT3du+a+t1XhJUxLpbWNv/PxvmVlj8Woi3/A9TKITspJL28
TvrKK+8Vy4dFU4fR8YUwqjais7LJ+jYdpBZMOJVqxm0zO7R9ijqwClJWVU7hEaS8
rz0rTpMzzhwzAZCZZBX0UVfvi2Mf/9uxEvKACbTZH8QkndhDizVuOX/LVQ+kM2UM
H0/bW12hKnxA9u7nZvl5iaH5RhJJ16KnDenJvl94HfFd+n3ZmvhLjuzBJaiUK94m
jSDEFE9rYT6tPGSTKTZ9zkm+lntAJhdr90xueC/wuXj+QpCROjUGba4K7pBmK6CT
FjpRbhcNwt9/Kq8s11ir0Sl/LAenLv01J3HikRKP2nU1HVwaENPkxdHoSgNWetYz
AlCtXuL45O6ujv5CEEOaTtv56VyepAThff474f2bgqcIGgQaz32YyZT7++zuK0jn
eEtMl9ek6oLtTgTR0ITLqExV/48rMwm/Piw8k0lIjTB4v9jXJ2Ho3fK0SCzA8IBm
Ap0RazF+YYwliCIB4EDR8XOPCpBXOJw/HmF8aPGiLsL8V/+3w2lRwdS7m2ML7CN7
iu/91XbJSoHaGk8QR2g91O4e5U2HOZdm5eAf2aI3+mJOW7N0needJsRMHCt9IJWM
zAwLjNbpav98O9fXmf1HcAEfX+fVVUyLh5x/9NzgUdV73YbWp6ewzQ0bsy+WD5Fu
h/feU0mQy6PWXXrsaBLvwQkie55DxdNES3x5mOisCp+wdXp5ET103FrSjPWN8WQa
DqmFqRvbu0PpoZn4cbIb+auxUR3oQXKGOXoBQZC3x73s2ZbG/E4dbQ975N0lYb7h
iZfnWk/bVfaZKgz3YsWdBvCMgPBFwiBqJFYbHZrg3ra8FUL4YwOrAoX1Z3y5/3+D
VFhMXIYQIxtAGyVHksm7IHzn/DrEIAeAKOTuz0BeNXXZG5HzL+Oo/IiYwnDz1Z5A
knG4c3PATwSlwxb7zmfhOIzKziAAnX1STDPp/h48MlgtxUOnti0rIDgz/cwyHiFT
ksDcEXXaDvbfr8xJocU4NQzcUPvrxjE32t4LC1iad2ZBcJi0XAswfmNVLleg7CRd
pK0Rrc0rTMqh4qe7UQRRBoEcYuqi6moxYHk6nqeor142lQWmuU3kObTHEM6VwS0p
MdK7/UOpXF4Mya5u8NYxdXa1v4cXcskeDhQfNGInXmmQk4N7ZAJCklegyUm0I1Cz
LUJF98IJseF/pF8ZpNIhytnkH0C9PnZZqO58UE+QZyUq3iLJqyM+VQXDlMy/vbo6
ahfQBRi0G/d2fS7SjRJmCGK5mpBK8l/mrNSQs1dZ/NRvAtrf6Ug4ODJPYqxuxe1c
ou4cggVgHU+3iNJLUnwrU1CC6vgAqIQP9bxRmiYQ0WsSycRMyWZKw4mdov2NS4vC
yIpOr6ztaKjT5quZf6X+WRc9GiLknPEngeXsURBn+devJk9hXKEhF6HL6Xb4N1sG
+Rw/h29lEkbcwe7IRDD4wY0wCT4QcS/8VTSbtUuEogfHmhNFWLWduUvV6GYjshTV
tDEZx1ALBUXWMwMfl23sCiESvO27xnY5Yhni57zGNZq5lVOiJKpnE1vSmWrCK9rd
MwDn8fUd7ndz8rCcfCf1RSkVfVIPnNwLPieyBeHX/DRcLXkiiVb25K13pLysm1iJ
Lw2Gh14ojQiDiPufsbKH/SKylqPztCXPA8LPdm3YgG90h30B/CdLS1HdZXOa3KLU
pF8sl+8Ugycp7A7PeqPoZPzmuLP+uGn7WvUSP68MaQPDbRUIIrJRa6SqZoH02Hwy
p93ldlKDXXcF4sDOQPYZelL/TLoIsZoMiup3MgBjXJEFh9VmzZmhpWjv2q9RJN3Q
GCOhjFJj3lKHbf3PqO3OOVWkwM2Vvn+wuad8Xyh2s4U3nibtgcDSWtAYhHxhvCZ+
cgwA6uoi1NdGVV3mmThZp2HBV7w1AzJMJ57CnhacgN3i+eVHJp/tppf7J+DeCOx+
JB/KOaud+Fruu9YcKFbm1aTQp98MBq2PMXbbCDjfs0sDIt5M6eZhRRgWVswA5sZZ
3bSKFDBTPe8FFSzR6OF/+A+/YCEHypKPf4M7kVSI+PVTFe+IOzvSGig+tKHRO6OW
TVi8V2565wmsREfTgz4NmwudUpSTY02rrTzGog/XIHb8BdO/0mkyu80gKdoPxa5R
/ogCkattHPrCQavQbeeg+mN/wwHmY0i1BkG575bml4A5b5FxdGqEzGizxDgnkflU
SGDrVEVX47VbR+POE3D/jrJp4qf+kqY6ZTWMKMEu1PiRLtOAngN6lwaKNbwLRsGk
PAke9TC55+qePO24TkxxHmGQXaupp+mpBNv9vwHKleQDX3FAsAi8BvEZQO1zPDH6
rVlTGgpR0Zx7gLDaz/yL+IbS1VuZcA5wmteBMoSAqLpySQw9nuYXotufe9yLWGnG
HGBAr8Xm1yUKUpCDMjRNIDTQULVVWC0v4hyQE2azGhgx42lYwx+YmawGcFa7KJC5
qXIKI3F4TqcT1nZY3HFZkAE245ak06hutre0sdFeft8SkBX6ePb4MkZ1d4AOJfvA
K5G66UF/WN0/ql7xhIgIZPo0XveuPhz7/KaVZ5O57M1CsYe4/h+IfJsG4bJBIuTd
zLMPwqkar9ApDQIpFH15qCAndopMMeVVNevG+5A1qCYjuloQkxdJF1OYTPoD1dbC
ZqDUrzt2swVxnODPj+4xjF3OtucxPPIz2dxTGh9QPri3oGJTXskd0SwS1E4A+Anl
xeaYQ77Q9CGK7ntJ7XoDZJfoUSDpFLSEcbX9wY7qLjBLlsQCbZLZlLdSRXunS94x
Kd948wq5WC0iFt3o9SV6qIWCdpBPTtkaQgTj7exOQNz2ptj+OvWC12B1X26wFMaf
VQBJGXLF5PewkwGuLv4lYAs05466bkLoU4rl8vp4hYgLCA9fPYDWdA+pQ93Lmqlh
jTB71flm6p/TxJcj7Sd3TaXxPP9+zsJWO/XUz/AOlzM5Sl34WXvlkspyjHGrNGaX
09k/J7MTPPJyyJCIsb6qmYfHJget/AQs/VJfjBJrH826kNatsi9nsjoCXCMo1+7e
gRRGCnsofrweOhEJfemtQLVDSHiDM7nm+1DJhrjJwdAcOofgcqv+y2HUd6nkvMeq
yro/KLrgmjdySFKdKmngzC0HCvA5Ru7dRQBSh/80NSLDJmeeBXbWoNe+GmyLrf7d
O4UBt75NViDvFU0dCJFjr3DpJrkTlawTXvw3ghR7qRJJhSFZzUZbz2g1fOtqyIy/
3uHbcqerHXmEyALYXaN1a9yxa3WVG5S1tfBuwM8N7Db8p/NiTBZ55Rl/MmY06AKy
dIaADUv09wHTee5GEtQMpxLGPZ6UO7YHlYrNJdj/zYEmcZTPc8eOLJvDlQbRqIfP
+REgwqhfOOKcWpWY4jmTeAY+Rf1XM2G3+Ibqy4f62AqNvnxNcDzBcnydZ+4BotnC
usYdorX0mRa8+nB9NuemKh/1WMK+up/HeqLIw63Ajlf+OC3mF2wiNpFg8geqofoH
SYddYjoT3Zjf4plHH27PIUGEnQv/Q8+hoIskzwtK8wvqNe7CW7dOa9pMdjLZ56J8
o+wf2QBoWaspMDa6syDe2orS3m6kWFG5DLrkNx6NcgsLwfptpANev1MsdUuJCQT6
Hwj9YTMPbNhPO/c8DazJZlFFpdC33RFnUfQcBkWIz+A=
`protect END_PROTECTED
