`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VgELT2C0MiS49RjrVtxfbMZVAXmJ+gzBtuVhNSnQ4WSyui5n0eMQ47p6yWJCk9gU
di/4VrCQcRN4GB+/HBCS2PDIGjOMgab2a30Dn8ZkXDu/RPUGLMKVwuzAmjAemuuY
yIxKMT1wKU6Ub4aFSIv3u/sJ7/fA9omNt/gU51NArb1DvOrvbi+AFGG80mkM333x
VKSJZn3RZFMq82VZClqra836EWjbQiR9qrBKSozCDXg/cmIW34LCPxPgBxqBrD+t
hF+3jdcNMTSbwAovhpaqEoXsh5070Mi0K/jgfNoZatJy0SC/x5Bm+OQqmqvP6I9d
1EoBlXrHicp2gnai5n0AbvHB+fA9+KOUy0cy8EBCV9NCELrmf+/GX1iQJkOJyK7i
JhR9MZt6C+I0RuT+wxOV5m2oCiWKyzYbjaZMZg9bwyFXQbDB/dxVy8IyoWWgFfg+
bHz4tFWg0b6tg7pwEHyLQyeAkXtDRiDtbSjCD8PShSt35w0ddOACRc5w9H0pncgq
hVwSW7ggs1vqg3wDv5VyvqRCqrV0lClqYUGIWqxLgy+ImMMx+rJ2eT+CKjM16h5C
tFE/BCyTJUF1WnBI8pJpbEOnpEuKGQlpfbwSxFbE9pc+f6QSKkwGqzyz02SKWpg5
AdeRTNroRxJozlpSMReB9NQxbkBCpoQnMVN5d4lkRwFoQigiLtYIwmwScKgRf1iP
aeOi8ex5UIW9s20y+dPD7Sey5/4b180Bw/6zKc2LadEelbmdBPtcj2ZiSFXGgSeH
dho30lUlLh2IFkEeXEVqxfMhowFTVpQYUZO877bmKv26d5qhfuOlPO9T1FJRUZTH
9maIk+PIna5cNooeMZ+dgXvaz4jq5pxu3ALhzijf1+S8HtCpje2BgWU+w4xuLu2a
DPaX1p6aDqYKtu813CpyTnD6wwkn4Pv9VUQRlVW/vwTIhKznoXzqFyezzUreyp5e
9M0FRvf/RCqc5IZkY9pz11j3ZmXgEK0eDilL/2xShV+EF9eBFCJinkwK9UqqgQmt
ErMrtQTTRsPrkS4w9qHst0ZXeOf5mp4Ck7Crg/YddETIgS+qqyuFlEIQAlqfXexC
p87x8yMN4AAcRv1xwlhMFI1soPP+AdPrO8sNAeoX4cuCngJr9nX6OnfdZdb/ZLQ+
lCynhevrRnKSmtyxfJtFT3aTIisWUWrHavSM7Ilf4StFRN2jA1S74foXWTwVeXas
uGmDPjf2JBaAV14FCDpn4XtwMauofxKT7jK2St7knb8qxl51hozQRqoMWpvEiYn5
fdxqDdvDuMgFtFYV1dr3y3fe5oE3SehuNy6bUdLYJNslPnWP3+pzkfNFITibfIvS
LKFdGwn6nUyvkfBsFh1jjlyg0cKx0JdkjwXpBDKh/5Lw9eCKMEl7waCKhLYFoWSl
HrqAP5heRCaUxsA6xT2eaSQr2SVoiGk7+o8CMEK1OOSidz44l/33oG9iPrVvywf4
06IQtV59MJELEJ1NtK39dAK5KoGJrQnas1qzeSiTmo4rNERM+z0emCsX5uwTjwo5
2HFhfV97vIt+vJ+WWUDC8dQVjMV8Kued80j8YiOEZJUX4UhO0QTj7UEpUPO080TO
Hz1dWZyTwm9idTuL8qjLSwBW3nMcgU4YGceVRD2JJRWvdBX2wyrj88+xicbJ/Hib
eYQPTLNrv/4t1uBTgFlaN066hzGFmXAuLWODgq7TxbqDwgf/YcUsTZebgZhUi+eW
N/JvFLVuzRTyfuKq3NludhTza9JGhmvlXIVKqszIzGQsxaegAtmB7Zh9xOjkrc5d
sZvT3agPBQ9bdWXVMrYk9Gz4xyi6mu26bTnWWXZMLEmdQktEwanvfCa4UJE2EJHN
PefvNFVBzhgQB8j8upyo5h4o+JItV63f30g4/luzKd4VC9/31+iXSWtdq0biWj4M
FJxYA0C53UWR17s9YUBGvLeimF5m34LcB4KgQh6bz9B7P4d1vqOS94vPDXL61xsv
Opv3LirXqBagLqXLZ1rvlt4gOUH4Ur5nEn8Gf1e+YL/R2Y/zZTfUyHfjvInzzvNh
O52bYwlSLfewoosNKQQHg2RTGj7bFT+LCJVVZ9i7luPta1lcJa2Zgcakxv4XISr7
vsEmO8AlyIE2jxT21fG0aJ7jPnTg/FFEvy7G7vzrtdZsFq/q1mM8e8eJdGfCtkpj
SMTEEfI3TJlmpOrm1Cjq16pPpR1rQQVsz+5MIDKSO3os3OvJBHjWXhox7T4w6sBb
sx6RUKfNcrwivz+AP9/bdNKG8g3V6fsJDhZCavKTCW4j0gr0REgfXZ60nPM8Fbzg
LA0vHgNVP6HH0Pzdpnl0LW7NuivVMWgHVfRld0PqjW7EIXrVz7T6BylU6lT9ZvFj
sS4WEwcfNTJu7PQ0UZpFzQIXKfEQdPwraRg8oBxH/NMoSYOt+DrBGM986V0Ql5hE
6bkYynaOTHmVix4zND80KX0ZwIe9ZJH+Tjm+ZGf/7y+s67P1UaLOe3V3EbWBk1Gb
LcvSwIpm/HnAJtI/REvEAq3s5/d2U+l9Ludyz0Ufcn96eyh8Y2jcT33H3Uxod/yh
FTO4fjNtcpG6loUFW6MM0xopfozcgKxfp3bnD8OLWVv5vBRC/7MDqwiadlsHcIAE
XgceRilnsMjxwHPXTuMMygyn7mBVQTynk4Sxq7tbb8lHGE/x1pg4oZFin3GbPzMt
B9KyLUMAN94nRvhsV7X6dNo+LEiXgGltiylZQoIGoDYTi/1w6LdIIW/kUaGYSbEJ
fyHp8pbAd6TavYahVfXANdpNmwgKwn7Wsb0AbahC31rJKLXRdGuzzWXzu7bAw+Pe
vJH8O7PS+f+ywCsaVD5R1ByO0pRP5GtKxOYWG+z4LjW/CxuV8Bh2kqglT8M2inpU
90BbxC9R6wpJudRBr0OUlwZhEiOF+Lv23jjcyJl7HNaqMA0RFg+qAih5HPO45aFz
FA1bOyxXN/bVGW2FEqKmnHeTJOckgzDEKLW/C2eFB1I1HCBKyVaAXq2SbJB9nNvE
cky51A8YncTormP7zCXqmZLrVqhfbzqxj1bi5jPAoZabyk/NAxo5d9yueril2eWu
n4HFw8wxya6xt/wAhOdUkcbHh6tDzYTpwr/tc++D0cyR3+ns2XZ4di13YQYNfd0R
+VAUaRf5fuFr3OpLo6/aZr6bkapJ02z073b3QBE/9u2BkAohUYidO4an9FaJw3xO
D3byC7xFOKGrO3Rx6PiWp0P6mTDis/R5A+PGstjZ+6qzKt3j63HZpEOfNJsYy0Yv
UAB8PLW8yJcJOvN+9zenls9RUH9gZHbOjjuC1T6myffTrprwLtckjgU5myFEzOz2
ERlzTSLphE1vi2OuIKWs1qiut0rR19fJIn0rS5kuhNQJbxXcBMio6O0qXBsUDaRN
BdStYMIWZrQz6vLOG3yZ1Q9h0dZ+vteX7iLHZg9jBNrqc1OPI529iU4l2JcbxZhx
/psR4KKIm7I/5pCXgktHZN3nVfQp8sXVq8PE23E7R/vfrVivym2Vxnrl6FT+FErF
TV8gJQzxj04+hTK5SiegPNiB+j45gMLogVFv83Q/ixUzZnRChSSAxXDyaaFops4W
RJwQBVOtY4Um49bySITK+9CGwU8TIu4INHeuu40hXsG2v7oWIChYmHhy6i5dmqI9
eeJBYfY0PDBfzdfiuf3o8AxoIrmYt53xS2qLFeBeYwt9VV1PsR79iPfFQqvVzg1o
6ljqd7grbaRKv4OIagDnDbMdv2m2iv4jF8PlbTOcPiEgyzCMar0Qts1p1wAG8shg
TSpna6gPOkhUbhNDbUmI6HvOiWoVtCiCMwuqQW264kBW0b4fi/GFdcjO6yE/mQiM
YsqAfVo0pdrSppj7aFAruy3U6c35nyjm8t6Vni409a6Oljgw6y6XroLAyysSSFvH
ARQv/ZTaXRWTKvzg99a0kS8MY/ZTrD/00R/AM225gHS2lt+8yoEj+sQOj7ghlHQ1
w6khgDotEp4N1h8DHUAyMXQsuIVXK2PceU1YG/7rIxPx3THMFz1hEoNCE0Ve4IWU
e5d6qJ9avNiovVIgkHCMC6cUVDDniKBMKKAG1x3owe7yJ87VRdv4ddeGgNvoa6aD
OfzofFHuePVmG56Z8+XXedgBOI7cSc5HagwGlmnmjlNDXUapuxjmpESD9uJsSGRP
6aNolnutwa1kX3AT0v2fpIonuhO88M03pueE070jO4LjCqJQ9ouuD5rqIsw1dIfg
Qe+/yMkf1CEFFWPO1ByfHzp7rl/u2kCiZrqeeFMtZeDXoAxiJ5QqrGVo3Za33hku
6zn6hSiu8Wn/p9umWRD6TiM7bS5C3B6uzzkcGUw2V+wV/gLH0Gx0dBs758nONrE4
12I/IofzOP3qsl+LNmmBItOh74j10JyqW7Hbu1BT5lU83gUZIi0o92gNRhWaSqKW
47p1kBNYmbVySh1ooTxQTLY4p2wTb+LQ7MdBnJCqAdEw5wjPVofxwzgcvouSj12n
2hzLCzxKDZB1guwISko7nn6BfJ8z+Fc2QZoPESaIkSmNyB3xwmxvI8iVe0BbisvS
629SITdZtgWneRp7xrF7pluy/Jx3ze2d35MlmGYWLLsJtwC/N5DDh6rIVF0lkftd
L8XgJMtMitisXX/TI9VYLUBR9eLDYXadEtXTg/rpgAIWLNjzwtz/Ng3qmCDe+ejS
4+gmtHTV0OicQ6QIGYn9+67ptxgH8hyvFpd1JJzb8SRVkjdpdw8kt8jsVRTxnlsD
Sagl+M6JkqDG6xhbluaeCIeGge6a1bNpOstVw0CdtunFLf7Cym1haHpbgj+lQDu3
WCYrs2UYTT07zC6Bkeb0NrA4KnzJJLd002vL6Y8D/y9sE9dY3sYRhlSLk/g5CDr3
Rdrzo3h/E3YgMXzneT+1EZAfVaeQvQExwGc8Y2btUSpQDfvNCh1uEDlU5Tk66mtt
qHJT5HThQYIBIesdwbIhTgO6DXuNoJFLXPhDkgG6eL1pDYkwDzg0CYd4/YcKv23l
yJ4+B1XZMp9jPkahHTKvMRkQmfTrq8YXS5zCSWlE14Ozom4i6HLiBf012PBATLgX
rxXDr7TUAO/WjwmL5nTbOQMQG1Zfqimc73EdYJ3rbOC9/i1o8cBbiXOGZWODsV7Q
K2BrSx2yTQSd/tZphANWXqWPiZM0uQTtgYmJHIgXZTzHVB0sPiAn6CvOQ/s4t7YW
O9ks8BGD6IOCK/D8o6+Y4UxjRx7IzP1UV0gmSkx/U4eRhvwQ6BzkJli98xwcAOfA
tNw+mGwfcqP3Zl1xCyZEfqsRE0FB8ocj2C+aYjpgRfayepgx50FIhjvsaktTlBJ5
d6meD1wFCGoOQXKN/0hOpDhDoI0kt2W7GM/Qu4xybhqkTBVQHuE0Q7jH0rvJd2bU
r2hDHvJBiFEq0lE+NHof7exvPg/7ShdVM8kI+u0U5neJGG/ykON5z+wi0vEeXNBi
P67SLCwMN+eWtH10oFrKHn9FX+IZkPIVnwMEwi47tMD2dj7aFSI4yamZ/heS014M
9hYLC7YuwmqWsBdPFbOb+ipVVmwbCI61OXKGmh4uSLcJfo5gBqAgNBuOlxnpJlQa
BKMsryFheEZRc1WkbQy11vv3R0vF6wq2OOlS1+IzgW+YcpT+9VaH+UycY5MH2LXI
S76ia+AGqOKFatgQtgedtk1QXd9TX+SXdV+dqszp4wnLAJCE9QPlB0KBENXIFWP5
1oXpVTs7O36+0tdy4CZhGL0BoQeEzj6X1CjQH+ker96uxxtSXkJIaCw4WJ8KB68H
G0fh1hH+RkVjEiL13Hpy2r/1UCw6O4+NKmMtiBXrku7NcVh9lTjx+8O3kwU6Kfth
JcLh3g/zhPqgKZzciAp6l1BMWsRer8+N/37GhXFrYJTzOLd5BCj4XLc5IyiWnxGS
NYbEO+JmfmtCaUbBVep/Y1pxbeoPFPy2Pj/Z2MHXbT/btDZFWP2I0x0T2ortAAA8
SRnkzo9kUaWTZp8ItXIK4StrE6944jvveMYHp0aNxNcsndl4uTCN5W/SBC6x3lJq
g5f8Qm2ezdvLxaCaCV72bAzsrOcUrHZsX8LHnwISHNEF2ZiKT4hMtu9qSqYkzurK
JVYl+MzbXYF5jsbpjK/qF8nwnlj4TPLonhc3Bu7hD5KQ0dGJXXmB9EyeQ1116Ech
+1KC0GcBgnVEArSydiHse/sg0A35LkDcLj7mVrLQamXSKtNFK4h3zJUNo1bFp8dR
53GjgMzc5B7GQU4z2KNcSV99Gj692J+bimBgKmHeH6g7xOynMcqs/dDFI7CJdooG
T7N3FObg3dEcNvrBj0GyBTb2Bjk/H2L60Iug7Rp2lBM0zCQ9nNEH662jMDe/ARxD
of2K5oCCy/2kwYaWzq9J9NJyXnZFx/kXrIjfxyY9M2eiyHqn5znTCe9+0bQxRo39
CJut3Oe/4IWXFKIzDgXG64iIP7pQyeS6+O7pTWQoGGipgiEwr6R1cR+AOjo7ipyC
gnk93N+S2PQLTw1JJeJTsWyyPhPehVhZpw86alyNtgwEyB1assh0fiURN8CwQRnc
MWymgc9spO2GIt8PqtnrmhjIOd4lQgch+CiU8vIXbqw/AYoKmvGZ815MTTLOUnG+
j5hx2OlAFzEN71vnOIl9E6ps1U7n4TSe4rH0YoTKTy1QQ4gsSI3Wl7nLL1cVmxGC
rYMf8wHkIIvxwsqr7QO2A/2Y9IyxOdQVh2175DRw+R+LftymrTjJ9HCWzzVkMtoF
x/MqjibloO+FWQAtcBMt8YTd5c0lDdf4z/a7gwOxZx+amBJIqs+Uh2FPyFDQkyRV
vDRvzj3fycJDeIcIlqTzll1hloQgFF85LOoKkiZwQaT2vDBSaKUelwU/NbWwJ2ZL
WkpGxieL4SXtqzmaFK5+VdFayV5964abOodOIGM5rjOHOK5w4M/oLcT5FlZ+4/z7
gJvkpP6sT7cFdcyBvcJSFAJE9dSJ0rdfKhFuTiwb5e9n05hhumpnGs5MLQZrGLCF
1VTE1YyBaZ70vejRIZSKBLte4/yD/H2Yp96W3snjCNegkXdO5YT7aQ+ue1HiOC+i
cnQCdsOrfsNk2QQnncg574YG9GXDs4TmZsiVB6qFX9UnEtPxYFxhYyr4W8DcYDSm
/yOV+elQVKHLmpxXQUYs6YabTQ/OhOUA0/ZZE7pTI8gzS95rwEhurWb0RkmCPjGV
HlUSyMoUatiDYgKSYEswIVoz3gTYy7fRst22G1DiRDrwAvpNL2FbXD1y/BD7SbU+
xIpXCle3CPgicaGf58kX1XWDZGh5hMQt1AYIEQCmwoEtoul/YN5JLknM6jEGJJbP
9nfctr/6YGYM9cJQbFtjBBBtT336J61Y0vQX7GxK+HxbsGaGugRrIO4N1uBoAbIB
xizBOsG6AcY3hQzq9UKS2A52qagks/WBKF44AsDpGZDv4BuU2zhxXaLZattrbW34
7nAUQkO/wVemcbKFTapoK8lep7H9jHZo76ZEXW1A8mAiLuPmZiTchnqVEt7yPOy5
4XaLw6aasrQrOh+Y+qY0wFcWjAQCCUH2lqYIRHmTWuHUAk38PYbECW/v5TltkNCL
X1Fh+QQWDa70gI42twEIrmCkKDZi9HOmLC30BI70AZ9JHqRVBv/kdU9UTiCHy6mV
/giqYWbW4PR+pQ4gq3zRgy1jRv18gjNgXbFLbQpkHLtZ2E5d4EfnjUEBTKYdQLot
XBJ1qDf1QTSHCcGZyafU2n+HpiuH+zp8+4rt+QEVSnwG6yZ4+QiSSC9L/yxzllcw
81bBgtAWh/cCtPKaFsK/Ledeb4eEzpqLmpFUgkJurPuDVr9iDuz+Lfpq7vvT2/9Z
9yZ3SrevUVjJ1Z3Owh1UCT2g1MsZmS+YjrBfInAhliL9xme1glERm4QqoDL2uTve
O7d9idTjA9lw7xgKtVaNbWGALReilAcqqOhaeQtpwgk5PcKONdpHCWR3GuyXdLK1
7lUdhaD/P1/gxmmw2aVa9TLOMsQPisvqiFLX92nskMwEbCPcB+6mCnGNjc2w0JlQ
mEIE4LHq5cDjHfwmMW72jcW+PEJWS/o2SDDxQQRJN7M2AKYoFAE5QfsisOJOolC0
suwz8zMiitcF853xEk1+KApWrBn5uYBgIN1/E/6/q1eFv0gfI005vIk9mMX1oxTQ
TWSpIKrUP8Uj6NmPSlDW4xxhrj+N9E4ih/JDADC+/ZPjhCRkQ6AdZ/AVOgjHIqhI
l2BXjFk1+bMkxY3A2f3zlk97LJ61NZpWGmvMS9uvf5TTbsrKP/aNUFIeHUG9UY48
jVcaEeh8GQuSTnNTeffRWFq4vT2MMRijUx2YgjbtkGfpdJ1mmrOF9fKnMGMRPirm
IG4GjCYOxB8RaB2hiKYZ2tgDujLBnMdVoBFjmEhPErlG318qkXHX8hslUW5wkvlo
+Vw3JKnCGLI1UQocx3UIOp6eeHtkxzVXjWTRb/2BGoS3oo25QLq2kOYtXpeaDdeY
8QXl2AOlN2DJiRG3Te/FW6fTnOKS5QMT/TNIFfufkWtxbaPohXP0CSSZRkGz3Gjf
099SY5q57k8ylmNd+uLMhHbXYLF+SCQcDrhx76u+YVgjzu3zqMBIDZjhuSJ03hgY
QZsuez0uve/rBdr6CBnQCC9xPUVCdPpOiT6xM3iRtqSfaKUIX3pCCVYCpj0HDGii
aMCTLFpvcpIpGpbyQA3L8xeLH/tWqKqX3CQdt5YNwujGxO5mw7OAOaX42mv9raBg
L/84ti9pb6UZvNsy9Xr0D07vbiQZWaaeRMWfvYaLyGyaRJf5NFHDj2eThuiFSbFB
z/c2C08V3lZ+nrsXdQTDYxDo9buI5TIJG3dwB4rHMwsoe/LuOQ4G2vicCCdD4SGo
qB/v0ALkMpYeUwGNw2/DdOsUaiYk3NHym9j7ay01IXCtY0WF+R2apz94le1FNuIw
3LlrTa46H0wssOCX+Cpi1LkQ5Sw57xXENFqNkHcVzkgqXi/bd3OnSVl6bcFmfhlU
+edAAEqTJYyXJNnLwHmtEmGEtY6DVd/a14wDJL0ZrSuFmxYtZJ7v1zROmiDFlMfN
2SjUhhmFrSb2qd0sUfFNhtLGxXMZ2m8sMsUhrjTstd3RHz1UH25efFtIz3WU4pE7
lluAPBJT0RuaNTcdP4fiLdWbiVVyBhKq9B8iPD0pgqjBVRrvuGTGSNbCzuE2eQe0
y5nhR/ZAPhym+aaiUUTIuSC5i1Asu7CBVWH7HS/baCfAMf1znQ1Dqoms2A5bZ3Rx
zea5hAmSCXov6ZS/Mkc0i28BRmKuaUi6+who+Z+qN1qcsVIpn2PpJ7pXq+ZpRVJA
7ilijoCgMBynukz78rtUqFDZEbH5/vMrS/hbICbiBnx7xyC/NpGnby82HuuMds3T
7Bs0z7kKiK7ambqmXz9fmMg3evijjkVcLdMKtleTjc41rQ1lXa4kh0axnkxYjNrU
PQozdRtjCPu3oMsNpSmW5gDbi/ECo7bOI5dR4aQVsCOLR1PykSG8DUnsi16ZAIhL
XV3bmc7S9gUWl4lTyvw0ClRpl8BnbSlbs9h7FkEpqiGS9d1oHDlYif7ucfKvfHTE
C7mXSrS++UV+SEbFXOtpB+gC6hDmHa/kJlVRUEVkKycOTKatsn2JJGoM4dBqij8G
kSnz/pyUlPKhduQS5ca2ZACtg+qt6IY9N3hQ24uLshFhHF9DKTJUEgdTWQE3QL+I
6GVe4L/Xynii3kT/ZqT5/13W/Ga7svSw9V31CM1mor462TyBMxFtUIWHB1HzLgri
hUCyNYzxlRanrL1eL+ifZXX38oXNMwWxxQ3XBiivnwWDv1lKABn+jMg9eluHIg0v
VJet0nRRF5N/bttM8o2/2qf7x6qsfHXnKTDQU6vXHIHBjCYVGRhocJVzK3R2pKa0
pys0MKmEX+2MlxCaI8+9mAkDitsa8mS0I3K92nzgCovBMGaubf2WzfyyYa8JbjS/
tYsFjiTGVmWrZBc6PHB8Hj4zCKKmscMvJCG93hf35NGnY2e3j4en6TpmfzLreK44
TpXquWY0UIR2xldNsPdk1G2RNGW9G0MccRDmnjKEzp9dHrOycATCyKzOIqeObOk7
ef9D4pB6bDHgSlSgChWbpyrdMobZsRBZ+XTi1s+StbutsWvM3SDdb1sm4ZN7FLGc
AN64Id6HNyNwiInT9nIuL/Dim6AjjTUSe5er4ascHnbE58MewdbaHKCZEmAxKNtJ
MwrfpjAR4UNCoUSIprwptSn+EZFqKwITyTfc5NXuuKuerOcMqn1WKLiKk7WeldTc
qmLW6/7rqIYuCwaASicf74FbCgIWFBi+g7G9CtHoJXpGaTkhQZIRiWPJDw4FwmQm
DV038lSkZcZqxtTEV7ZxVdDku5K/CJD3nkICQ6VBZJqTme7zfclDOfQ0OkLnuhwp
+goYPWsV5wiFJLXG6ywgCl1XjSpOp+G4oRPSUliDsuJn2wknesSWx0FjKyh+xcD5
cKFMKK2M/kcyJXuc1yCbQrecDqOWyK1Gci93Sl49aGEIV/vOfjt6ecVqYnT/zj7Z
NfHMkjms4+V5lEhyKm1CjZ5AWnNupFX+G2duFyNaoHuinbtXZzoPMbHM8n8dBoUz
62oYVTR7nHe5/4rYRq/C4H66ntZiVBwE7/G63rLCVQeIi3JIx9ycpQbUwqscqHhw
JskQt2QpSPwQf0YrA8JjD/OOBkXwWUmPClF5H11UaXdxgOQaV6lmoocHXFaenYug
Syog+ih1jbYe8PFUioYCPfEwL7Uk0ssFbZxN8WuUSJwX0aul9tQex56rZ7N/PScd
KTgYValc/VpjElxjdTASKLwBJiiC5tUyzhRhT/rcx8rqvViwatYFrdBR8pSPNUoO
60lBr0SRzviCSfzwMOb5wN2US0jvCE/aYXHhFNQHXZNVGnwt31WAPdBEgFFcGXC4
WhTfrT2mnE8HvuHUWe5sYvTAVDYRH6n5GcG3l7khKky31O2dw1BKf7FU/tqYU21D
y1gdouf76fUynMh+S/Orp72Ixw9+F1MN5WU47tm8HM+0tjZ3pwQoC9dKRdkj/Hqi
Bx52fGLmC1C7GuM/S+xrjd/2WRK/hkNswNBs9e8ChE+Y7fKEfq5ZcjXOSVWJHdij
qfkePQOil1uGMWu+Oy7utGQ15rRd6oURmdDkB4cWp7n1jYdpDa2XtS8zQEsvLvaS
mfzDCYtKV7cdlbceooLgFkO0kYB1WWuwHpxTzCMWSfqgH4B92mYcUxQd4gGTRwEo
oBux7j2Uw9N9/G9VQvss8YS034iBvc9YlN189T0n2Z+k5irba9D8fQ0YNPRuXcjv
O3wKbsmcJhRenkD0Oahtf1bvpKMSdj0grQNvrZWx6eagtHPRLa7EuL+U8nF0T/Gj
KIS0ImQaDdITMieL/JEpvpKbEp0UPIAm29fv0q6VWtJ4NXCjymTGHYzprUW+nKBs
tsvSE3DeKJtPG+jmbqtcRcKZXWULEOloHN+BLUphbhR7GFgyhtAiCPadovomN6kS
o/8SJiOe268HxI7VVEIKO+MmY8G2AaolOZ3fWXrtXdyWfa+HDs3kZn9ihAO3tauW
YASg/Q/QN3+hRkkmiqySIBrUNCq4Fj8Fg+oMiVrPgb0Td3jno/290MhbPkdKz7/A
ayVFCip7awPodvaHkfat+4GbvordR2lPaUHhyUzjZRRU9RcrHmUX0mwJhVIfTHdq
iVBP/qAxAtzocxMMTUaFalrcy9G+qCaTSBBXR4r8njGwEQmyKOkQURWFohwMMwyf
TonP3cyO7vS4PpKVuWAcLdrCB0SKm/UNR1DuFpehdjpdwlHAhSUZJ5qrCB4UDdli
sIOOkvO3Ib+Rf6ep/IzMg+PworysFSqKcdKcx1hK/sR4nS4McT2cQYrVcsSnB3aT
T8c1QgE0wPqAtzhFrQIadvnZI/kzehp/NTJ/me41RjuZMnH98xsxhpDYK2b8Ilgx
LrtLCIEmPS41RrIIu2F1Vmm/BzEpIXvl4uwwldP7jv80Y6aCFyECnqmOwa1NA9g8
YtAgy/6Ag4sSN0D0LIYLgWblXaKIolo5RbrMvOcGG54NKPwBz+Y9vYqEnmVwRx9L
TSVxkx2uzB9Zi7KSHDFf9zRVKtrPHLyIUl5ICFnWde7+dLytg/iMfL880gKYfv2s
FkGLnQnTGzaMMbBNtKC0m720wrK1Q/rC2MUTizKUx5+4E82vwF4fI63vULw85DgY
Dk2NwlLdd52apfhS5Hat5tnP6QIrjAeISd3V2P1n07+UTEsK1gNBni8Lo+WITI3S
HudxLEIl4ckyQl1av+En+M4X1+RXnnRx5r0HRYK49/PEnxGuXdlTPem7t6q32eBY
bJ9MiKNjk9fR26JC2J3VDcKixeVb9G0lv7w59VO2cTkosgyHTxuCiAC3pzd6IROF
7zJfICiBYlObMaEpoTk1mEjQ+QQkRKJSTP/OMmMCipRR9AGaECJWb7TfBEnUOUUB
cnnsWc+4XmVcWAlALtwgjOKRAqoicXg6x3YmVvg7h59AVPQx3MPdv1FiR35T880O
pseZKxiEuxgfM5EKuywcj8JxJZ+U1fT7aYIIpGniTRtQo+Vn1kkvV9Og414N+TVq
DUEX6g5eJ/frLxtK310mGJSeM3g5eS8Kpwq91vGkvXBF6yOljm7BSuaBrwPFmkaP
cF32FzXfRgEaPsQFiiZOvBlJaIT2EGmQwoUuyAcyM7hTNYF3e6CY38HbZr2/jSi2
piciIYyYrJzQmikxcVDyqQ==
`protect END_PROTECTED
