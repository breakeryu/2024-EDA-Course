`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RAn7p50GrZo6jhQasEx1TLl83u2aAo33ISDdHhS58OHJZaRLPJyT4AzVnJsKugLk
qzDaKup/3MOTcv+I2d4dZT4jooMOTIBirosubX0v5HbU8KKpqIalKh6rvjHTAtNr
cllsjkq2HLc5nHCoDzxTlG1LdCRdAU9vRs2QfB7E8gnePsp/HGSGyitcs0nj3P1g
Ybbh6h6wXzHFoZqUVBEuBDPu4I7V+WVRfdVhZYt89uNb0iK0nZUMTCyAENaT1asE
NTOF+cMjTjBr2X57+yXK+kxHjczMASi7GqESpBXnVm5qK8ldDhZXkp4M+K1KUxAn
Y1N6Xpl/r7FMHDPjP2hXN9oP7Mcmgs+DPYoRd8KTn4HxkZkJG85QfKiMDXVX3Qhy
AdjDHcnCmS3jUy85gKWEpk2u/r41Dh1DF4tIdvU3HsoZp9RweWqem0/Pk3o5mHKa
Yyvj17sd2ypWgw4sg9a43X4dVcO323yyxF0dT3nFLG4fk/sVQEhhJvTlQzK7xJxO
2vNoBz9Y9VPxOZS60IkKHzjZTHHbE+vNdQnJqN4PcEEYnc88dAg3tXY3Odlbl9EZ
6+7CeiwIlR3dXie6LDSr1l+y5lQ9cxTYpIKb7jR09RYHR2CWyOSqSScXazLYYWJU
AW1nmmKVjDrm+ya5SLEayCt8U6OwKQYm0kVbO9wM8B3GXQLAi2050MYeoksaYv+A
lsWmfWAf8ai/6upfIHytOs7RUKNdjPbwFy3JWr5mDKjQlCRR+C1PtHHmzueDBdV6
yFnSmif5+X39YNG7m5xrZrs5Agw1auBAaCJR9dfkwbPpJqu4zHNvri8ma+OClW9u
+8pWlXf6C3m/8fVsz91OhgifXfSSk6UObTRM5v63lqc=
`protect END_PROTECTED
