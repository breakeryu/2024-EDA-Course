`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kh1ve3V6vhTwcfb+27Uh4qYob/MrP603NGN8UxAk0zrMwA9oh1lJF45pHzAeBzgp
iDgL6Au+2IXO38Rx39UIxOb1lOP1zIH3KJyG4aZLzhmQQh1caaVXiPEpDYOTyv+O
YOawq/nRQuDq8XPOm6i+SfWe1ig4ljSA6f13560W+j5zokI+ucjSVIgt30DEyR0I
h2hkU3yPl//QhIwC8oiBvc99PEXZcXgYv1PS+2GNM3uezh6Etx3zukcpRw+TZ58Z
HUyRIgbGEmZV+FPjUIL8bNBpzDDgPWswE8BdTzd3MPlJtHePINwzN6+hTsJWSFVG
Ui2k7JJcXyJaVysbwovRavhGX2pHf67YwF11fzx0yQULO+YBV5wq03iCdtXxQn4S
sg9WfjK6RqIqLAF8TCH0v7es2M3Bc47XUboBaDa4dXzlPXFTCU2bxGNy6ZXvQxKc
6XsQQMiv7Jr363dUdKL/kSQI7b76Ewr37qPOFSx/OxacFnAyislYp1VXZFwiQ4VX
vvsLyvccUG4zZ/kLhe1wbXnO1+01Dnjc+K9s4dVTxJHHP6HL5aF/yyrvs209VcCh
qXE+2JvkHiqyCBLO+Ghoysba0nnUQfstDBVXLNEsyumU2sI10Uv09g6Q9oiPJ2gS
Kz8aRpkMZKKq0twWbMHXAZnC5QD2S/6BAVwJpwO6jULQaB7Agij5n56aiNV216Df
41Shj/lC/naQ6+dvKqGjxK42YNURb8KGvqsktAPyS/UQmxX+KwWWa6LqjJPP9mUD
42jtMZEYcLd9EapwKo+ShZcqJLWdP0soqmyAkCf7sVmqFiiZXcpSMtglr7dQ5Flj
YRAnAcfEtsMJrH6b9BysmNbXPU5vxt8iuTI7HI1tqvkrrHcxiO6qB5lz2zXvSUNX
ccE3nzv+RtLq5/2Sit7XAd7cc/0Aw3xmFvAHc3Ri2K1siVjZFxxgph0jDsRYnyKD
nReRNsAeTHDwS41QJbboH+fVtSrQ1eTqhmdKr9jnnzdtyrgd0vJ2TD+f0G60rx7M
l8NCLZJjA7JZhGaexo86sikdYvrFZkb8QZkjZs7zQqSPDxzeTbABxisXE86FWfLG
EcXmz2gTX+XZIEbTZgzMUzA1GkF/Wx0W4p/O0lbAxt6NK82kzQoSyOipKA1xrsDA
wvmmC6PeJiitB5Bs4+MXtSXQDGAdtGU4DG+wKvUoPbXEU0nC0foVK8HaoyxtpjJe
px62r8N0Nxa7O2zYb4HsEulbEWMYL3ERLUucG6wGUfSXzXi/xZKd5iSp0H16Ohid
Bl995GPN/ktnQsS4/t80f/ccb8QkgXl3HnKbZhH1nSHr+pwh5wl2PYtMmfWZmUtO
n3wy8YdkMRPU3J5qGGjI4zr5MrN801FkDUnp2RfxKraAgTp29lIQOZ7xxfsrkVO0
SK3/JOXh0CH8lxj1++YK2CyRG0mp+/Nb27Aqnb2VwUnq9x+etvw0WOz3ijh+XypV
9yEe5/V2zXX8qzbKJpP6zTGuqCtEkB2sJuyA/eYgGAF1SyZ9ClBwZLfjLkV1GSnK
y9V+3DXO8He83rv3xhKy0+LoC4xcx81Nlyc+OGrsh/y4rVyxcplFousXhl8LLsWr
iSNXca+2MgYBP53IyXshQt3uBk9aFmpe4TZWklYnveO+1oicaciF9KKjzoiOwdv3
Kmd1UiU0HyB6BlnUM03tnPvGZ8FXfteA5GqiRxtImv1RqyEHMKEsMQZP3WAU8ME0
1O4EPd6nL0wMh2kmFRmSPid6oEXsjiFr63nqJJnBqn/bTiBgdHfV6Mor7Z/HkaYX
NZJndkoZMO2Zw6JrJJ2JGToY7o0GHDZywrsvOrBV0KZypxfJoKa9gvEhwAZNlJ3l
32e0A5tl8ApNicrnQbh2HdH05fiphWUxWw4eiCAq4UeWhlVe7aUDNhQStaRSaHvR
EmiOA/1rEqaOgHc5r4IEqdtx7Y28naBCL6WiWPlNkSa5fRniTD/cYKWW6boK4dyJ
Am+R1t736nxaXdJ2IVWaayJZTDSFoau6HgBtWtSHh84jioR8koUr+Pv0+OgOSA29
5CnILdRTdpK664J6TT/SxFtwzU9Jl1MR6peP92eg6kYylaCTl1rjB5S9Yn+GCtE3
PGrb3mvLq0UU6GV/925wZ2Ck+gWB+urz/E9GZrQmkaiiX021AJgqltES1nR6sQAy
wtQCgvQ1SS3FoYNsXJqLa/QJRmtPY/VrRil5pTVGbW1KzfsWWVVb6PBU69vYl5DU
kjVbduhwUA3HlOhPIoVhlzew+y8ptJXYRC8XY1XvgZ1MJzohziSYBEqUpCG653UF
NVzkiSNAv4aeNrjg2tRf+uBJZhTtFy9QxDK/gYYFrsfZXZ5srWqRx7m3DifxrrEw
3UdQGfquB9rn8Dfz+y6MJDawW+OWXEC+53jlmh5DeZNk9xZGBSEe0v9hRz5+wxHi
m/4eeRslSospk2eeFX4xNew0lVuUXrAF9C/9NqX7rY9dLJRnplC8cNAt1mH9VFhM
Hh41U+1c9icVVqb7ixPJYM27wwj01UcZiiL9ok6ikj3Dox8YocOYBV7dcBvQMAoE
OOYDfLMSp6+eUX072I7gYCsx7Sc0yMM4Di5GFk4g392/dh0P9IcmCrPgB+0wTGgX
AUYfekufdQItw4B3nORXxdTJ3gcLIg53/hpD21X0iJ0J7ZKFS2sdOhq5zDrjBjZl
3wH3ouFNhJPkaYQ8sfIr4hEm5RwRQqaKU9kq6pQtR2cs+mZuuAAOGnzd0GV188BQ
gmxBoA0PbyPUfDhxTReQpICSifBQwvjm2Weve5CXBf60fOui0et8RdowFU4s2IEf
Qq/90pwyKagGFWMRvlwpKejM50f7bULgBkqqvdtBM4XcrF9yoMI7q0M2hpP8lom5
4/EuKjM0IHsPbgS3OXiCAIibO0yYLmQ9nMRS5ej9GaP74aJVNJwKDfquRYMaH8gZ
2deooTS9uBD52oOlGsqZr0QMlcxRt/sv0CDg1kCcQC1EYpsPBOiYLYb/oCdp9bur
MvXseaqGQ9JCPZCvODTlXeNLWnHbVrneiKa/J72Q/tomsbCqOJAHAVCEsyWtjkNL
itH3iOYjmKIbLAHEbWz0BJ0kY6cVv2lI14np0um+jHX7CEW6vDZ7psrGdqwX5bqX
eRxF435a4RSWq60s+DYigudm7ENMCPGEFI8lCJJHYNfOfLajhLkQOuN2aWI3o91x
WXLGMb+tzbKEU02UFi9GZklI1ORD3cN9aI3pgJAuRgxU1S55ohNyD01KfaJPVuHX
G21NQ1I85GgmH3cGT4TNlW2zFyZ2HXaKad55y0Q7DGNHkIQmAE+7VI4E5hUhbPFR
8qXiB8ocMLLMFzk7Z9bvxGcs5UECixpKKj/LZ8UVEkPU/YmWTQnLFGqK+mWRx+ly
JoeZqysj2ekCsj4+b8r403ZLnT3bDvOOhM/TLNEbR4GKZ2QHzILkWkGYKmTMEg4B
LxcuMIiS13OdLdeT/kpg0ni5ryDP2eRT2N+H/JV17eEUgNd/dRYWhR6wnfxIlepa
qXi7v4QqOHfdmpmZ1RgO2FLGPppwV1NyRyLv+BCZrx1dXy7A4xpioDbx1QxUa7qa
N+KU9V5rjfELeVKKhKwjXAyE9jmoErWXCGcLk2QmojoEvQiWFWEbkk2dnvyYpOAy
NDjXPDZOx3eiqQXinEMTtpvECQwOG5oUXfHI9srj7cTZF2vNqPrZTCUjXiieXIBT
WulZwRaaAffpXWd22piOL7hfTvNT8mVxDU2lQFrr8BRbd+1qYM+fGSMXnf0pTGYJ
ieDeU/bEXIxYAf5q1FhtX0Re2lblg/DG973U5dd8yEvEkTCU6yj+tXviuZsqOn1i
OJ6rMMK4VsTpYU8XMoF55WdR8v4Dn2B6eupBe0pkJ382iHplNb8xcb+dch0SbI3K
CcHp3CGyZ7f/h4IdaukTllStHDGunUzC1GHCZI8EAWejI49jplMZfr049xxDb/gj
tnPyTBD5HpHtiMfTj8Rm4Hx/qYbsstjET5UxEG4jbg5Hif/UbJ1cROuWPwwGkWxs
23PI7xMWmO+wcH116PAVno43HjB8GxjGgu+7RNNL56edG8iCXU4pf6cCNxZiIRJW
pCc83/MZS4QhDJiGP/NCDKPP9CsIQlOBraXF56vdLZpXMmGXaq3S7vWxLW2eZFdc
c6uKq6cd7VFYj/HrRQxP2ZM01bFiYlHMTBAdH+mm6mz7QKEOUn5aLOTQVDOdc/Pb
P44ube3eFMZTwA44xKxXYZxiqibXmWkJcqnC70nT/6Cx4q6z2KECCtLePj+UbFjC
LkHbPqaIFFM7wBR9u9eam8ZJhCFB3K47knPgpXVIGJL2S3tKJ1a18qoGjf44Ufn1
ZDKJu6KfpZh3RmOmDMqsDbOjV3yw47fJUhxVzJ7WpSORIUoBeiLgV9ZqPd2NZcjY
8tCH0LKOl9NWIGpLcE5gvFoCnr7V6c2bq2lh9VlSN5szM5/X9Ka+V8PmuE9WYJEB
l+Nna7ZQna7qkByGsM0H+f8YgzGpm6b1j8lfb6y+jGiucm1V/23oEAmeo8/JYdev
zUaF9oHi+pcmisYf8pYNwKuUkGNdDHZ7yOzjjoukighgCuUttqdf+qd2uEI6NUIW
4H263lkhPi1jEGiFXDit5fAYyULOtzaY55NE0D/KLTMlODhQLdvx+YSSvimThzqq
pvbJ+pANzTpZLkcSd/j1RRiKsNsNy+zjzeBmUEuCRDEnM3/1oz74fURnDbJpA8pU
S3IMwIm1Ncy9O0uyHN/P0ONwv7fF+H52Gqc01Q/OjCV8yxh/nlgmWBe9liJhoI0o
PZaZKXhGEWFN42FVRhV2tTL9TTfxX33kCYkXlBh0OafgbSrlby5IXbt+ABrJtSAZ
JrY2AAVymFKDGq5gZYXv3pP8Gd0/ejvr90MstG7jqs0sepNkB7Q0vJiOFjy364dR
2xCnRslarrs5P6HmWM3+3CblmBUDA1/6KvmFfQh+aysPdJhxCJ+42B+O+Bl1RopP
OPcRjkZGq9Gab4WFV4gXWuOo93e/RuJVhq1mo9l6NAanNijJoxk78DqQXlzPrObv
7aWh3T4lhzC0yrsSSZgcTkx7LKsSLhTVWH6V+Oe07uqxEVTlMcN/qy25RJBhYmn6
IYDAZhOSOHqfUCaHL2phQ+Yum7xxoIkENU0Ov6/VnG89tcy5c9+yyzA7pwDAk4Uq
VtuAabQ+vB/TY6bwwtuXw8/11blCWfJaJ3aAII1Vh7n0UT2AzTM0i7UovcF8FOVs
vT47cRI4y8ZbK239cqb9HDf55u1HW2930Qt6r2fGcK6qcxJ8FYkgqa9PftxT/9xr
SYwjVscKq31vrUgQ8Vh4hr+ic3CVVDbhseVNkunnJWRJrRPBHhLk4wsHmGYWFCmo
LOYcmyCv0mTKrBIVvWvNoQuwXgY5Uo+1kbBcCavjOFYL/2meZPhFDrlawIVLa4T6
mZLrtAddwrIhHkPbEx09XqWbRhxB71GcI/ZIgAYCLfuQe93g787KWYvaB+UOuRQ9
jnrqey+eVkORJKR7G5telXasMhc6IWcaffRBHZG6pQsBQA/BUeWQq0IEOeWE5vkX
nFouDE4ke8ijqnxmE78yNL/afePZzngTp4VrWXopLARk2OMpNZidiIrlaMTXBs+u
5UFm+daUbNgfC+b6uhJ5WCRxmsz3/KLfdSmm3g7954yIM5NVcx5+2h8wlnRNaRDy
IAG/yFCwMR4jFPPUS+biuXEAY3sMTSM5u1Qqh6SYLkRs/5V2DECv9saIzb+XFgSq
3D+LY0QkwbP0Fb5HkDUMwKwQe0nUeEeiIrtY2uYV9MA9N6tcDPo9zx6uVrp5XHeg
4NkrIPni9TnKm5tWhX1Xrvm/tVDf+YXcu5pxyLbVyW7WNT2DurIW53YO/94qDqAg
TnHtnDUtnBAGhlrLyE12Bsq7s1wUV1xFG3fX2byTZ5DXbdPFvXevD2wnKPi1CrDI
+8YoDc5XphgEpurJ/ph4txpbyu7Vjqmj+i3klZq8+f9gJT0LV72Sg1Z0Za9QyS9q
D3fH4WEahrJd7TKf9dRrmbEgs3K6olZIBR2tUQPlcwCjzXolgLpJKK89SIhjXkRR
I9ZyVY+WArzGD042pBrZ6tIPd0lHjAQzQu6jn3gnTlKxrBFUV+0X5z2RDzxBUBHq
83Ihu6bD7HBSGGCB4ArAGcr9GS2FHN/ut7ICN5YWuiBllYh/b/GCJ/oQtQYDeSHn
3oCJzrUqypcCq8H1Jbunqk78EXSwrD1pjRsR2ZwXz+FSGF/l7meDcPOFNrMxjg6K
vYIJ2aEaZIio3kW24posACgKrO5zsgulyMGTfPtZtaJBkIr5i69+VI8M6DfhgwPs
hblZKk5Ih56tGQJOx+VtsvKwoDRctWA7cM3Bfryqpoi9WbXFuw/2iDsEZR79ceH6
BzBZVp2vbi6KZwOEnY1VM4U69RFHPx9bNmvW8YS+csPXh81dTIFBi6g7DNOBQDZ8
AqeLj+4VVgZsrtiED8VEU/Tv81OEFQMd+oTujDA9Kq+iWV/ISshvLtYOzJW/zaaP
OhHmK8GKgmQqcJNyz0blU7DC7yjDO6TsEHdbPQb3L75qZrYzQjMtBpF6H/yDDiHO
OsW9TXbSrajz4hpudLIZyf5SRa6jGmHd7TjnB5Wq+PKpM6Y+I0+GOWzlE3gm5LcZ
N4q8kPp8pNeH5QAGwS9R8igCjtD2bQVV+jiqqWHiDsalIfO7fT7+nKE8XkvxPQ5m
5CUTvcxn2DjkGVFwCYemckPqPQuVutum6HQZ0w9f8SGciwrXwf1aN5/qalaWg2WU
vY21+Y2mKFsvehUOk69ydATA+mC2D7Yi47XBS0Fb3BlBsyT7miBjFCXBoBk9fTtM
unsmcH09+JJE8nY9frVOQzbqDOJUcZ0Ui6Gsz7BMzfSID25WTSC2Mj1YJCvZf0pl
PMx2jjHlpbU56oRziJT26tfYsUa8+emDouTilOpODzvMMNfc77uvIiDIEDdpKtsL
OqiZeOkNtKj9WRuSjV5sW7S2GwoYnXnF6wZBzD18D40q4Vlu/2kdJ17aH0Hv5FDd
eMvxQfU15QOvyPpupYKIB0sAon8QSIjZcG9lvDJMcbrXVSuDQW3EP0+v5QH53jrJ
lWW+j3MNv6Bhap5pRtCtnIc+gfh/caAI/CHkQwr5SN5jMdudM56k+b7irrywLNPL
ruoXUM8FKnuS3pH4cq5FE4u+isma3iAwAYCrW+a89ga+/YYv9jdpuaWh9GkWDmd+
7vNmNVmGdITc2ETxseIgyyw4XspcgbrVzt5gtE5q157r6mjKuqwuCrMd1ABxfW9i
703gY2BCfmZo2yv9N6OWbNOq1Vjcs94smy141gVSpvn789dFLD+vE0xr2G83lqN9
LeOwhMD0kRMg5n26bUVeeH/vKWlYIakQ4oGV/ecQGj/32onpqbI/NBSbx4RE7d1x
jEJKnGMPfIYTWnqIWdXA2TZmiLGm+1y7qN2sdgNPXbpn5NzDCR6vSN4DCcTkzVAU
+7wn0uFnX41gMCNh6woKN3GkS9AID+Qo7AofoCOCYH+XX7Q5jEq51P4PZ82N1TWb
Q35tq+hIzFTo+b9aKIBlzUsiDOZipRiE6X5PAPiqeoKlUzRs9kV/pgo+3NDDxTNo
n/MEjAR7As2YwtNxWX3mgKXrlUY5aAY4L5sLysgWq3ix2f56IAxzwlYoCE+nnA9X
1dP5+d5dQKKgRVO7EdKztfAf8j9Jsbtrtd6JxUIwoClKvttRfYnzUIcvB0SuL3ow
top3WFCGEsgtoR333syN7NpuOR5zj7VWGwzI4TBwj9Hja5OkNJJ7214b5uk/LNF8
F29+C9NFOeSXpkOJrJqYizY4azfAKB8idEtErrkFaIFvWQbd2i1JWTVviw5y8tm+
q2iBJ2Kg/CNZS3jIkbHTunFucU+vsqQZwOiXHUMbu1SEV/OsIjzcdkeNsstiXAzT
S7hzvwG1K2SaY75TaueGkHuagN5WQDbEBBYysUEfhJ6ncDnagyMyFAxM5H/dRHga
tXMo3+/IfbEDD+eC7DSsPx/b/uEElCwyBeVNNJpUjfEBhfkx/MPWeIMuOB2usZUF
2vzeqn9M9e63JrJfXeEEGcwGLmII/IanCljf/b1txGD3fzeY/ZZFmlCA4e5HIlCz
8j7ItJWuGEyHifo0PIZ+J6yfu8wyiZjr/rJ3BfEEMmRLdlqKIJttZ3wjxSpjlrO7
TyKtXltB/1v3up1eaXYsJH0j2GGY4ZcTpzYfNNkzQHGzVXuXcQAa3C8GgvljK7tW
WpJv4BDOLid/PCvMKID4eN+0nOmoyqeJHERy1lmGwxu04/GC5bI4UQIVNyV3n5qE
ntlA0WIkbfx5R7Pt3ktXxUp4Sns72teM1GbTOh1SokrA6sOYGWHrlYpG1u6nLSjq
Hw0pE0MGFSMr5k10g/OtrtPLEpaxnLUscQHQ0dECScdWAAlEwXfO09Cao37S0RJy
wdK3r2uVm+8MJcP9p0hc61dwlg2LrxF/Z5Mn2I9fEbuy8/bJa9WJKCD2dCKP3f4e
t5nCxttkn+jbqBMhx933uod1Miaynz7UQiXsI4TQYpcKz1fd9qcPbjOEELyTG2i9
9RXaMFlNw7KZBtPrNFeEooxCAG1N42eQpt0haKEf+7OAWrilqF3c0RHfZ+hnpfKo
iyG+CTjz8pGZMClEWYxLz7Z8u+j29dJM+Ehn7vA7npPZ9r9VV/2qNcNfaOsgdp0o
46Gqjn4H+kiyZdBbBlaTCOsPj0dn+tPQuUec/gcSfpR/xoQPQimci8Gg7O9Qdomj
jFqIcrUngE3qxBm0wddq/A0iReRLXyusaeeOUAmkkZf8H6BfUrYvvK8EQ41IrTan
h9I5wsb2Mns7yE7k2paDpEfTctB8z0Ur6KdGl7HLmbGgXJMmq52fF+0LAdIf815S
ibOsg0ZKCvBb9QT5FddjbKM/r5Pv5zQ/GF1A7gE89ASMMkd0ziH4oyJMaG1y1DWk
S35wLw7pAqOQeM9Ow+0f1+SynPNqbjiY+2uVLQywsOfcWVL/bwaG9qMk7WfBzC9S
Y0RLtrkJ3rS2FPxZI1HFJFncYW6vkOPm39LX3ilI00cH17YrhuWdeTfKjLOscK8B
Q9dESfBaHMwCQ4DdCyXQqiNEbvOK8pGhTOQnwF3/a8XcPizS4OQzuj8fqeTG34M+
xZMEb7xJ0nK7lPPJ0DgQxdVn33W++D9Ayz7YDc07UnPY9ZAafDtSMhD9W7tR7nhJ
7YvqCXf11NttJPFF9egEOQ377MnpyFC/INhkv95Sx/dGHWQrLJqIcI5uLY3/het1
+r3GluNhJtASY8lGoAKU3rplCKL3LtRTN9kS+gFgR7rLN1qeXYvvs6K+W+oCqGN5
Jq9auybf+Mjn/IT6HeymcYgc3PUIrIq8ZfDBxeGysCg7Xs82kdSfo6JDVgDWbYyY
VOc6hugai/Ii/tD2xK3OqNRcTxAgMklIha6HSn7tAAPwUQ3/eUwvmGT+LQjMgJq+
YQYh97QSIKjRCrFrSR4E7FJd8XKuTpuEA3ysDq4OVYpGBh5VrseRZt7x+hHy3WeI
CKPbfbJ6BVeVFoMXPz1UkUGIeW7ROMpEqJB3oRt0vSzrtezh0fgh/9J3DFl/FVQF
8VmGS79U/O+E6fQYnehi+9hAIGM/+AY/6J22NCchiRKI5KxF4++5d2Hn7HlFcuWk
CncN7Pgqx8Kko1lvvPr+9zXTm+hX0FAGGtIZMMrd8SRs00cemVessiiKoCGprNaz
a7DjwmaAEvTMhma5DQAW/SvY0I+axQ+s0WqQgsBdyWrH1LYIQIJJ18rRsH8IWX+G
NfACqErNTb+MzeiKQgMhQ4Kb+xlLi803lGg81N8DuYjs/C1mO8rWGPJqbZ0jejX3
XU55hp69XmRsvZj8pxd8b7roCSbPn0AiREi0xzvy7RyGxk6T9DmEPOrJs47PnJv3
ZK8i6BDUVRSDPb2BDvrR1/84pmT8a5x02el9cVTZbhoI1+DeSG0IOcdoKnDFNDjV
+XurE/acIKmGfaY+knqrEb8fLffDR2LMFAboQiH+6DMo9pCZrdT5jO4JoLbfBEeO
Ptejk6cDU9CYBlyQTMweFtGTcAEzjeN1WZS2OXPN/3GYeJovVj2slRrD+LOY5PUT
48Ay6FGasAIkqdTiAFwk36Xu0Z3nAZ7ZtUCLySFt54vYC2AS4bvxP/fmeX4LNRQS
yvR8uoRblW3p06Nk6Pn/HM10qVsnwzf5GwDcOETwmoCsWMYDDhfeyIdq29K5vuDV
57at3d+hrr6CNI2iPKjhIk4jE4qncuEpbLGuLUiE7C2Xk50Kv9r7JR5I7HQYPlW7
/Y2Mhl1udPbXZ/hTdAOtGS/GSlv/lfaHPgZO8X9grnknlGM2gdCGpRHUXdqAQW5/
3ebxFMt6DfZlK024BywkS2fl5tBlPrALCNOhXuihlMF90xD5fPoPFb/6KfHna+9Z
P/Ys4iBgySI2kiwXgvJFbxrOZ8hv2/y9Afmllf+/ab20oo95A0NFFNTTX/qu7bFh
mASmmziVbb28AuKBAlahgIxuFjd9RU/91wqsy3LL1czUXpJ4U3lw37QE/Qhxk5cZ
9AGtu1AmEq62niYt7hJfzA3VqcQaOOXLVylo9MoqivpsWjWmxWUrnEP9/hxGOJXu
VR9JoQNYSupHxi27XI5F8+1HejXniBGYGH14SKip0UHXydp45ZuQllOXZu8DAe2K
5I4rlGfe8UhzBlNK0tGUt1/o5Etj6KOn5KERY6wd0JfAVdMBxIhLQCBsb7e3EIcm
PQnwqDTEAxnEgcCLB2b59WOzg0dT7ybmY96tEM7KoYsGNaQ+6v/seUVICYAnhcxS
yjwCqoVNBjzLp/6qM4T5e8W3HSYlzargPm/Omdh35v+M9x9mZ1it0AU+tOP21kWh
MtTKMt96fV50upzJkI+SqijSRiULe/Wr+KWkmE7OXNoGjzi85Ap5Sp476qKuXC6r
14Ian8BnwYSzg2slSg7BE615nc2QcHcu7i8eu9Ddj0Laoa44F2pyTPSYG9wDZYP2
usWY/xMmwS9R9txa6BZK8VLHPdGSOnl6fH9nSq7F9ZFQN9DfxCPPo0bfr2H9U8W6
xhbCpVEaM+YPGsqgiyNvxAMZqvublPFDIQnmuNBmnuVh/Y1OSneW8fy6QfYRhg59
lMcjTJ33ng3vgENuT9hd67SgMh6pkmIu8/Gtv48BPTO9drQrnHl1x29bSQPQwuHc
976zLqJ/APgfmJN4k/bFfZb2LFmF0ODRRfl1EQ66l+vKEPpOeQmGj3ifTkaswqBj
SSMLvLyvxwUzNmQ2wIWqo7Jw1p2W8wkf/zgh6OM+H9fpJ0BoSawNM4leR1lJBIlv
F7/k3eg6JCpB3iJzy4gtX67tnbS9ViOlIkA9HHALIuLi5WiY1vu6m/h4f55zoJAo
pNSAjOTcf+fAm9asgUPkX2JV5wV7O3C9v9ZCUm14aA7TyjeGXgSoC+wRCXTCo8yS
KpZ2NUsRV9OzuknjcX9UGLRo8r019C43eg9Ioql4ikB2771XAvt8f9dptC5/bpme
4sj3lfQRtSDbo7VNXGCpT1rq1cy/fmdYLT870tjc3FY27U4nZ2mVnZfg/lJwpe8u
dJaNehOD6PXWBTyOiaPLT9HgD9npvDM0uExmfy6vWRdUfUaT1JzLR6bPgAjmfmWA
JMMHlLQyd+6e4/f/gzjJCxMB3Y/o0Zc1KZa+m8QhuJYUHyW5aPgEYKg+HEfrq9Oj
w8a4ZxsaFZPhncRybfIq7YpOabcs23D1rz4hQHf0H3phJQ8s1mOjTQKRC3jN+WgS
x0BVpuUK7t6UtTMsO2Gc2cuQsHew6opsvW+RHAnpWzKc4N+ZWrq4MZHHZxN6RNwL
KK5rCuMht5JpnF9atrhkKlXxf4pk3QB4Bdpia+Ok6pWzuisDbVQXn4WW2CU7yH+T
xteEOVzaCUjX9deCVArLan+hSO+5TIP7b1htEiDQEo7lOlamNTiSZ0N8rWwUn8iP
oD4YqkPM/dm5zxDZlNCll2OOISbyIuFiVQOBxN8sXbQuD0MGPRM/iPFIv7ASUXLh
BLzSIKw15dXVrZphnjcLjHLhe4mEbacmZG0g1OHhTqcljIlYBKtfeism6Tci+QSU
Vh3LguuDKzh0YxXP+lCXSOhGGY+RmS8dwQe+Yu/cSWTB6diiYrJP7/NuAs7IFQeN
8fELZlRsRwVtx56fQTflsY+C9mNSbaa2h38wknKGrCJBA2WCkdXlYVwyUI79wJEm
TLVi6lDhu9c15qiiBcIgJWVe5x9G8eLO4Aa8Zs/0HM4BP9DvarihIEVhAXU9dD/G
eUYT2IaqYVtFNJIf1UoBubbgjUo71B3Kzc5ovF4u4vqG2zr13r4IrwP8InM3+SNQ
cQ6FCT+ZJT8hPIa3y3KHm3ZWHnzp2B7QLu+axp/lFaMC7+1kHDEdf8QQS24eeCwd
A5e53xQIsvD85hyDe9zmSJg7N2xbq/1JnEJP8fvfxMsNEFKo8lpB90KdyMq5WERZ
DTxrHfkMxVxHiBmbYuZxTluggOFCQTLfVLDN9Gp0/7tFOcAbT6luqGZHhiPiiFIS
WVIkbKta7M4UVEQ7blTiLpMYkPEp+4zpqzFBsROkkEeNNpcwRDNLTCN71SWwwQQ+
SmPnQBueKpBw+VxnkPE0hIQiPaWxrrw9G2BlwchiV14SI4ZDapCIWSuDt8h3NziG
rYFtjXNh92I6BAc525JrbBHkP3So0qqgcH8Kg6FsZysLV7ZP/JgxwNZjHyV8NLod
lOQDsDtFfblvgs3mpX2zzz13OwyfFTrmDfEWKvV6zuBtirPywNZx98mbawsGRxSS
8nwS0/dPaXcT61DDVZ38KJL2cCewNkGw0ApG7zIfAce/ZY3qjgekWN/4kpWLUeKn
QyFfHbUHtnbJdRVbQ+LkDFIHrM8sKdsYpKewpDFc42isfEOgBAy/iREkLgQT/KZ5
ZZOSWaPUpFl7+Ezgde3IK8kvmqOozBmyQ+/FhjUnfZ/R7kpVNy9S9N0DU8vll72c
TYG/7NA4IdG22TsUbKIwcujuWDVBKp+pwalWdhXwy/8+M2dFlCpopOgWfaenSS5h
clUKVVwsbleyvPAI2r0cSSkdXNUOEgM0HgjzdtOG2+30EG7FLeL33jjVV45AYVxW
Z5v5+B2JsGcPzDjoHyhF+Rtx3vhGF/o7uX59DF69CUP/vBtSBn1iJSlKMHkX82Me
rvdnDQsDX/4LM8DGv3LmhS2m9e03WL2FhW1SdN9t06hx2G8nByjaP3l5zHQ3iPCY
kQ27TmkKuHqMViT8J1d37LVWoLADqxnPdpp3l+f/C2GQPdFUr7coJxVwy/azq3PX
CRSLI8F4Nt0PjIx1wxAuJw==
`protect END_PROTECTED
