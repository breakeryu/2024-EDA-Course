`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RRsuFp8Idquds6ujBVWpXF8gCUa8InlcFY/NZBB9kZKkPdb6NJcL3ng58du8MwVd
h7Lupqs/VjYexEoummbfSGIXyzDSABukqnMthNBP9mDQf2ffaRxOVt8JIlOcgyyC
4NnD7QERlCFX1zQAqvzOPIgn83ntdruoP2nFYkm98+I7fouDXvH9zv/iIU2Q69AF
KWCKDZrGqZ32tq4x+vZt78nA14RqLVwM7dJKUOBDHjhYOvo2fhwGKhCthfUWhh9U
XA7jNLj+EZHe2tV/R9v2UdMM0KpMOF0th28nGGBIihjzEaiojxh0vgkd+pTaWvId
dri0l9Hj3ofvwr8e2mjh3+CRM5W0K2gvU5jZ7dO1sMCPVQdlBHa1WiTunMvfF9GP
7aU2oLYfVGz9GS5MHhLSl4+VR36SHI+2y82C57ezsqhwtbjNhPunMSoL32c0sQLQ
MW+74yZ2lZVdDGk90MhfWt9qpF1+CTVAVZy1KzJ4NstM2GPBrJPCQwMMp4Mn0BR7
69tw6jYZOpuzrS+bpf1eGvuI1NcWTyIHUYRY3aAgMOAO09IPxbH8Ngn2CoSLUm2p
7y9SFG8npDwBg55moeNIJ0p4ry6rKF+LKYbnycFZH2ucL6fPYDCYKx2I3zyBuSro
uZaS6+PGE2WL9jJOVk+ZYUMI0jZExhbzOTZgKtcE1b1hXmgIOFv/L7pdfTfN1UFU
`protect END_PROTECTED
