`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6JP+vMTrd470+CWazE4N3jeW+51mjXThKlDDQDkphRYVUE9MhrM2Xx8PfICQVYxs
2/ZGdiEEAuLGSlUeTRhWdy8/nI/Ugy5c9kwJEP5qAkeIm0Ou86qcO+kqDgaJ7QdU
R6li4gQXKaZWrQlHyGIILsE9mxGsuROTO1Qcz/amycuNEaGDz27R8NHg3S54m8KF
3CRT5BRa42QLljniByNvcMrwZKYnPHtRGuEryetS96QEM6Z0I2yGzIsUT77YAWA1
Ogy1JUVeA+OMQXB78kvf1y9RgxDNMSdvcjdGsxSUm8pT45DB7yUd7MTTkeM243Rq
sF9GIrsQY9siP9O442iTbhPstWatn/DFExMwG4sx4XlrMDiKiHe9HhEQkS0QNJGW
ojNxO3yCmNcjKbuG5Zpt8iNXQ5uuEV7Ini9TBpT/XwMWTAaooFLzdLXGuPRc4770
/Coynz/NbsHFn9fESbzFclHwdcfZ9YYWx3UZAmXxPFabk30R+ePa5TlZJu0RiYtT
nVeKNBNz9Zr5rWvjDCqspS3GiBbzoLFqYTzf8AS/X7lnw8To2CZHGDce5zMNJurp
OTGL2q/1TI28VaI8MnJWG/LANQ9DTQMLBia4Hpoc4mqS0FzfPhBjaLNxTIczkLI3
z01SK645Z13gGuyQiO1V2Z04ezxZDEj3hr6CLmZASeC5XG4nAloCE8YGXA6O2uxL
J5cHX57c1LPm6y97oJoKNDX8Q8M6jHxFTFYiZ4FDVS1qp/RJRm/rkXXtmW6ayxDh
J9CmMIUhUpjm/j1GLK8LQS5/19QPgeeJpRew0iiuBNAkPtqY3KqK7dCH+Yc/XJ3V
WM7ncW7NlfXWDSJZh0OogBAmKPMa2U+xEb5xMEBbMRh76mOsi+VFS4WgJhIiE2c5
Gjs4CyAr0QgZ19X/CMxTuYO861WKuet7N2rPrso6WY7FUF3z/bNop7lgLpmwNCkq
i9TiVhjTMOLG/SEuP4Yv8GnsI+sNeABW561gATryhzypn0WutVYE0cUeE1dsHsDk
YdT5aMmSOy24oFeSOZzo18kiXii0fBW4dntaRBYEHzUcwUbm4NWcuMGngaS8Df7K
o25kCpK/HMQE4Gw0f/AgolQBgE8siqsbN0jWU427bd2Q522VDZGu1cmetwPV7avQ
EBTQdmxNbk4nTluPx5YmZNs/bT6HOWzg3wxLTwYgO5PtLM2vCtUh4S4Z1M1uQi97
6V64M6YRKyLF9yd7paCDI01g/gFc+7ljTmGSmPrdY0AqvfwSiCtk1wUzL7OzFT9e
Ri+D6l7OrzMIUnvrLMzXop1GheyyQAvdejafxxgWetD+SNfESZhmoVsniFJOySeq
6cpyYZKP39ZetClFN71oYKOi4tpg3jcq/N7BSuLTYLyAuahr7gh1mAzcbDDXqpwH
WnSB+YxNIBp+1szz5SxX6xDJ1OeNFIOfF6Lrl06ZviHCD5XsMogTpNkFxLAx94vj
Fl+hl+EUAssG0xJxL6zAHE7hUhtty1t83+otH+mlYdZN658DIcLhsuEl2tqWTZrq
UP2dJMnbod3xU/w5vUFeFYMZvgcuSJH2sja6vEt/M4nDA6D7pslICQlBregxgo5t
YsaaW6RsU0i7cd/+Em0t1iBEHdgD5+4Eu5zwejhhimF/o7kRQJyYmUx6qGoWHOEo
o1K6WtaJoZyYbcI5G6Gf258ngcEleb+PNfCZfg77gb1owqT+gHH8W5v89HiLRtfI
2D+p6YzBR+vFakdpzc+OFFkckQY7XH1pkvmxP859ownbzAt2S9sjOT8sy+MHa0Kx
2dk0dbpe0C1IJAPdsEKV49TklzzArUdqza/28I0OH2AAjAKL2CF95WY6FVLllWN6
tEOHxTOrObCRj+CAM5jKT4jufAlWIjjsd0LDMYRcHwalPO07StDcvAhTgiUeuajI
zWpCFdIltGcnYpgdVCzlMqGU5CZMerMtrWZdocPjZl3V+e292DghgMpJToJA8DUi
VXCAMoDrZSNxIf52M5nc/Zo8YIZyncQ71f3nNVqb8vP6wjGyeCqdKtHOxQDKzXQ+
gJAxHpZBsiAltozonMUU+9lpKLMy6vb890IIcOsnBt6sjzGzP/2AGst/HQcW3YT/
xLdlu1yrwG2F8xo9eQRLWukNDUUQvVyM0+A4t6nUmkFMqi6zMy7qJ3IsSGkBcfIT
gwlgD9ZSXe7DYMkCOMzHc986RwlxC+Lm65ooq1gKMxsrJrkbaxQjq7bcH3wGx/b/
rES6ZwtzKhCK6V8MUeywCuemjFBGsJwfiPlkPVaDna/ckiBvKzDPTmbbnNDLE7yw
irmQawrJGcXLaAAIHEwi4BvSfiGDPKAm7Sc7lZ+9uLVEwjmS3yN6j39gcm1JXP2M
dht81rxOwsVomfl+2yE6CBHjKpC0BMY/jF/Clwpp642RhVn8zmZYFZPchMOcVj6m
A6/h5zOwB0NvGp7AMgLCMzrucmAi9LLQlOkpj1Zuv8i9SKBQIW+JkXaW+KfTIAHC
a+zQCTixnb3+ICrbANFye8N7H598LG1vzmxQsH/eyorxg/8H+OQxHjcZ+HVjGi1K
2T50SsodIM3ywALceYeawuakWT+RdXaIRYJCI0JK+RMLKlIxLHJe6SpBftqGscFU
CuOt4LYEXuV3x+EmhOkiQUtRMKHDPCzep3fMrMOEBZnXHY62a2vOQwFDy6/Io5Hs
xRe1SCSVyZ41d2tqwiAR1Y8ZwsNdlBWRFW0E8tdu+n7FIOvQDOxhne55PnAKiC7W
LBbq4wxMdf8kj6rsvaX2xCw/+BIJR1KtZnezDYhH8CHjUY7IlXYZvzuGbPKkFdvB
L+4imURqJYJNr+F3zbbomU+D43BFBZWnrVzIbEhkV+YKX5b9U/F0UAIElwpMBu6Q
nvoO+A1+STC+QSXUasycAxxu7auc1uePJzTSV2TEzZ8JOj2peljOHmb26q4ZWdtG
m8T6TTTVFondEIjoUbVoQ1j9UG8Dn75CG9Us53rAyperR1Fr8tWkg63UzKA7yqBZ
VdHi5fo6ondceh3VFwIJK6YrkjMUEZXabxkxaFQftwP4w2IwTWQFvDIGHNvS707B
5HsENlbXn4h+dQcv+LWSbZ5pGJfNjiZbiPAD1tokuZt+z85wJLOexb7okNc7dl9Y
mZcLxKrJvaHSBw86J7IJ8u3Hg6YQQ/W4NjbrSpChc+XNFKr/rpZVW+exdgjiVU89
IU/JYnOBCsNFQgL75YIk/Fj6NFMwLyBVv8+IrNQLtRECiaawBzEShDjB0IBZJ/P1
FQ7XPYxcm85eMcLzqCFyggg9Q3nUhbNXJQASN8botpvjm5xzGclQSNutFN8PKfgV
RMD+DvL9nhcjeUcxYHO+MNAH0duV93QExGCsLAAjCvdSjmNx24xgjbqbEKkTIjH6
Mp7J5rHLYgFXssWviJEsZMD0P6YICwGbH5IUaUBR8aCLsGVpqh7pFeH7DBrLZafF
tmLUWrnWsE+PljP1oTCJfLPAcYRBmPQpROcHRQbwCRyeJ5MwOWk1+NE7YygRH3jr
4z5WTgCc5g/ox5uegtyo1tMlfhv4xl/w2VS4bjbzodEmNQDkZTY5HU2SYh9xUBeZ
WzOebQYASw5347gN9nQ5FrsqTr+NzIg+9HDPmuzkvfjQKgXn/VTyeylsIoJoh6JK
BDcH0AOlDoqWsq2ty9YbFzWozRXr863ur2VFdBa2LJaPxnc1bzmCK6ekFFC065O3
eotaIAaf2xslRMvzeRrxjS9UDJpIJzzH5Vok2iFbcxS7tyl7j8iBb9sap5gbunws
SbfdAQD1lvlMNIemSY1iLN1szpNmTC8hhmVBi5hzHen0PqX9z5+STYuFsPE4N6nT
8KhmfzWZuk91Y3Yo5UMHGpdlcWuuaIIAk5zvfjjf58f4r9y3bGFCNwiJF2WIjg8i
IhYFrK5sc3Y9JWi6GHA2JnoBX7LBRicXx2TVCb5lT3vKedhYiKJB2xT92bNiMKKL
BR3qoBj14D5ErS+sGZIeRzjDHHMRhJxy3keUj3xbff5nNLtWaIR2CzMkSUgAuRgS
qJfQ46+RHD0WxZO7zdMq5SAPfsFnzS+HRa2zLQ3it3ii9euTp6kuRsOElxycRmJy
uSgLqFAQiCH4aJ0IKuSaNkYXOAilX3SdPI6ua/cl+jVAjA7Axbq1kiwuCXcmrdio
f0LLiU6pEN+e5mHTuZuONm+nJS1KdBFJVpsUP/8gxGeqqImNCXefrcL7MeTr9aBO
ceD3zy10r7qW+Yj/HXnHLL+DB+j+FTnxdGUnNzcKM0y839Cz4ISKPrxmwDFpkXGB
ijvl9URCbMqoZ0j/kgi67HQRW4i3kWQLK7nreYxcyhr5H7L8zrlIx2wDVrexEIfe
BHBR00oY8951T7lZdoRJLOIx7Iw5SICVobd1q3CXpEWhb5QKNBvWJdq7Bg82+glu
Sx4X26KAelccU4xqZ+rfxqBRIFBJmK+NAZRHW4UbxX36laH7kIGzuc2S5hIiUhdV
fIsg+XmR6neMYCDbaxcKNR3wx5yYmujLC2bXunLZb/Ylt22x8RDhxe4jm1V1RrBS
Qrc6SpMfVlgqRA1wadJPSIlUMugfcBSDbqcUFUa2Uy7j+xMUydB5xIyuC4txOO43
AGhME40D1QlBFOMhmtwtRjzEAgY+flFeUv3yqEIez4WE4EpOJ5jdjiOpQHcPPviK
9er9+HAuOHr1FDvyhTMWv9yhV1XUMfd/ECp46tI6FVvXTBomjbs8RdXwxexNxsqi
s0sJtS9XruIZVmlzcPgdGeQa5XAR5YIc9+nYMJgRI7MRK8/ufJ8Q3p5h7NGMM6if
m9heN0swKaHVm8KNf7TEjIhWjlHvCgBjX0ITuODsYznAZg3H4l0NDtvOWWttxCt/
44slcSQt4NUt86qZ0FII8f/Bl+30bjryxh3W0lfR9ZK2+JfvcYJMfHQl+rXBStDN
l5HOvDSw6zTx75m9CrgwyIxvIN38v5bPv1nzXlwSWCe6K6c0XXEx58DthtvigzKe
nwqS4Vxvx7MZZxXzE2PzGxUJNhWgTvWha3yb8uHbc+UB42sMx6Tv5q/SIWC28+LI
7FvC+wzwMPXDIu5HkGWyUh6FS/z3/+UMgAgzV8SUGVkRarfM8skEVGvSL15StxH5
JrltFE0mqxXt7ON9RMeDF/bYHnYQNz1hufBIORLyR4gaBUgtRwfs08aS2y0u7gTC
T3719mkYG74m8yY2YkOcVMg3RzctdE1U705wqOwZo5ugCGpdvJWV1YmHJbb72DOq
xRMu7WSSA2mn60pMuDs1qX/pErD3X9s5aLLMUbNs3O/qRhAPYb4G9+EcdNf6EsH0
JwUBGADUuKSH/Hby8QhakSkTF2LVDG/GDjfg04TVRSbaQ3jTbiDpykhojusYFDVz
iny8JCuR1xoSFjrooyAzl6iVKCDT3yoMfhJgG83XgAdyQJBMlthVpaEGO9JDxLu1
wGDfLPIaKABRWE3EEVLWlQ6OH+iTHMfR9htkkL4eZXJ2b4x4LGeLhsVp2eLPZrBf
OBFFLnpZru9PO2Ty2uxNvxpB0kWgzcOd7W8M2gXzwgxuer/m2MaQILWaXkMtJ33W
tMbFmaHZnBxGf3PfmtTnTusrTa58YN0ssfn4PmXg9oS2Wr7MPoT/KyC7CXWhBYzC
XD9/1iDZ1JNJMg9qBziiRTq6I8iTnxdIF66dZTGzmIsgHpZ1ezlV9CY10Mx3xL3p
QvQV4qnuy0zVb0pTjm1Bh7hTAK6FmOFNdWhQy7U7aBX3/utUNIdZMDNF9CKTeeqG
1q5XH9LQZYigU49TiU9yd/CeUpsELatJqheTQuc5GDD/tlPuHwlT1LRRi/u8Rgul
eEBXxuNv2B35yFTduPLH4BUtUeIRJ/bdvdg7nWucGPJzeUOXhktCmrNBbjx1Mx64
AAgXvEmikHL5op/GqZIuKLv2+v3OZZvDYngiVrFM2OmXGQTeJe0BltKECegJf9M1
vjrI0bi0k0hPMD5TXicIHJFeTo4X++52ZB4WSCd3L9AMqRkiz2cRYMzPpvpvWSG4
uKsPoXW1IcpjOm/w5XG871tXaeM3GP27FrV+ML+mzyWeS7YuuDY6mi+mnMAHw53j
sP64zyWT3c9QshlCOFl4ubjWnqH6lH48JE9leVQ6znaucjiv9HCLhTqs0sAXKHqr
ef/i227HTOt6b9jR6h62bV5nCH+7+GRCAD/YjhgXLR+su6UFEXjkheKgWwfOn6IO
sVBW+g4B4T/yWDL2WBuw6WJe8vwntXUqDeu9xndj5w3uEMKJmEzA2trZKapmGSSA
7gzovBnzh4M8B5OAh6F3lMT3d8N5hBGQp5DYPhUpKtDLQ26hzPytxYtCgpga7MjT
J8T5R376ZCSYf+EgPk5HYmjmzfVfhZ3bbLZUv3I952cQmaOeiOKkfUxpJY/BYykf
Zq/5/sYEGbD63nCVfeePVEpZVmwNdapAgAQd+qA9+i7b2SJtWA3MDRk9ATyS/l4n
TJJiIzRPRN975IV3MHxQiG1PlKxMCvRdlCyYulghGc/vJcTGbqB/LN/6VDrBOVfJ
DfeNiNC9MJrHdc8k3hH75r8GZahKyjJWxGmrwz5oFbSbpKABEkoxe9TzrUcce0Qv
qS1Bg0JRn4i/QeDlcWBlChD4ubr5+em7OPFzfNR+YgQp2PengFTDzElxm3PKpJdx
I1uQd0QqrnVx5u26Kdet/pjCckoDwPTVswU0GT/HQwbWvzE4z5LiQ+XwPAyN3VCW
ftjvX7b5rK+k7LsIdPlJIHERY/sl6bfcHFKLYZaaStDcrObJJa8Eapl6TdYyDIAm
2fqt3n0ADwkcnitf0b6v3sLjN8gkL965GLKYl8ja58+MKkc97hnIQSlN4MiZ9zX3
wa4LgM4HUzfq6VzXFjqlYWX4jrgMs/zGY+2V5a4Ml5pgY+3DVLV0tXMI8qGv7KN4
fc3vDEgDhH+vesnSiyrN4R+Htqq22TaI5pGoupoHavE0yvROmuOm87Bld2YX3Cj/
D1aTQbsdNhkHFkpyZrAuJcvlw7Hg8any3stGhKuMW6/p9QhupkLD13qsCF+Aip4U
oW+2n7+kNUXjv6VUS+IzgV6bjlNEeMEZjf573R/U2XtMGKcTrQYTvupsiMirj5WH
9zHXGdZt2o2e5Uowg6hY0Hc42Lopp0YOvuFJeNqDrcxaxGoKA7yCVfEdzPpA63sf
p5xJOktefT716QpGja8dnJJPSsIWHEAubTQmXM0pfvai5ALf+dbZf/7VLWQ+eD6g
daAkBDKyHyjO9PRex5o/KGo4MF5RRkSqpDi1KMVYhmPWtWu3PZMUZNNdOr+qXAaf
g6OK/oG+Kdm59eRgMprG5g==
`protect END_PROTECTED
