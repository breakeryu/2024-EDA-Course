`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ayH6w+DD5xAidXHwqN5DoSPtHjNhI826iLsP06AfO7v2hQHHVqRFLrtBx3iYyNiO
mRXw/4mFBmU1nIrvjvpCWHRzZjcLVWjY0YYa+/7JlHgC1JY5TSZJ9uZFl17Ory5e
p24g+H/pArken73MDot/MUV5+ecHR8Dn0YlwOmcMAlNJcASOH75yA1O7O00T8idX
+w2pxuX4EgZuomcuV6u5mWty7aT7vivUy5m/1SY8/t65JN83wD/QrWLNm5JsLUMT
9SCNFeQ79yUgEgXrxCS/THOxlufpvNT9bi01HDMSG5mrEhwny1k9kccmfVt+Zqcw
Un/0pwHfk1Y4K9eTJYm5woOEe5TJEkxQ8BjHgKr63gRdRN8Y5Z8KI5IplEcMjull
aP5conhsvR+yveOFdBAVP+MhEtvT9mgI+APKVhXlE6vEIYIocDeViv2CtOLQRgQK
Mty8IMXVo+N8VamQOyvEbssJmXEZNBEO0cJnKy9PIqtMsmceIJKbDhL+67PauvCy
s8bu6xfaLnlnJSS7m3A4IM6K7wFLhe/pUrdlWHLZEt31YbrsKf+LCaQzWbdc3x2a
QWww8LBPRhAhokVHDOHi35CiQxvsicjxMtaOljduHoFmcOnma1nSdlo8tFtI5oDs
+RHfCBwgRQcYUBXwlOxbwU2f+8mc/PaF0Pr/bj3K/uKBapW/qYL7BGa741MapOwL
Q0xYVTkR45gF0KzH32skBsElo/swDu6QdZy8f+Xxa6JcT9iPp5Rs/RfBRmHYEXlX
fbmtD3RlJqWFNoIL6rqfEmxAwwZgzkWtwofRgpj/Kj0vNTSOS3fAVAktZ/c9WHZo
EzTOWr3CKqAl+2zu5SKKWHFsJjBhy0QDJjXIS+2LZnVxQsGQ5+pSnE5Cgt8JzUhr
`protect END_PROTECTED
