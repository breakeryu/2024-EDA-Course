`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47WubS1NepnVW0mardkAD2U4q4Y1Nfbg3dJKcSZ5/Ryhc2tpWpewxk4TF/ac5gge
3YjJXL+RF1dc3PhSIHBFuCkRhT41q8uxNDv5Gwg4i3zjoaMZ71nVS8BLAYBAQ9ca
oQhhv/1B4n/E/YP24npKQz+L0NPlUxXXGYzgmQdhsgwmRdPPhhnV2SZo2aLAwvx8
`protect END_PROTECTED
