`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2v87ImbzZVBuzirxDr3urlOAwWU/OmHxv5d4aCjkHqrbG/agVAsgczT/UmsuhSN0
65ViI6KCkLVoT8R9NS1WnZbFnFlwwMWX0Cmo1BHnL2Xu2JyOkOWM4d0mbib/QUBr
6eH8UmewGzPlrHKmySFpxyjLQdlxr+IwEKTrDZ8tQteGgyOgmsSxEg0JCfjRksMg
ZxJ0wPwWcDehAgGPpn4TYDFI3E940fz+USU0IDaPmlwH3JsQi4OeY0T8CCDL5LVR
hwAdAlsLwFa1Ix7lkTlN2KubNJw6okLCqmiUIaVLdJiYuLDgOwR0X6D3+YCWa8mJ
7IkzZOwlvvMYB87v02z/8bOa67gb2RU5WLBdlPP80rihy/h6TrZwvmB99OilJseg
/PB7VwOH+o7LEVePGcijTevDEjBVZhI6Abt5/M8FsmyRjBenY7bm2gUMKlizrF/s
sW5nxh+Ty28EWIHfFRIhHWr2ISzXoshTBSh4LZHPlI4RlfvZJDFyAXx3rr1rlKVL
fNniBERXnBp05qybkTyj0v+W/QHDuN5HSoghwvClS2Vr7KGjE+n7uhzE2fYxzRUd
keb1A/7Pc8uqtsUgwW7F10A0Zgv2EfC4pIGu01BfMDroLOrcy1p8ls/ZXN6CAw2m
tY8vogJ2BmVkop+EsAlmBh/e2529YGCfUImaLG83JlBSPoujAzDMaOKy1ScXzVlK
g3pw10moRWaXo4W8Y6LwIglrIMlkxdGDlev8au8lNEaGslL+tE+8Nvp2i9nOyI42
QcDvtwEOmq9UWLQwQMnl4HVIYHc2Z+2w0fmnW9CJC/fPAHePtVHb/yERrv2yyOwg
MygTG0L3KJpNPcUUD2FCaS6MVHYcFd5Ql22Il6Ft4v+022tL57jqhgWAodxKHS10
uIuS9AEy6Lewwx02a/rz1Jk3ugtnb9LvwWT3yQHIeeXULn8HES4nbCTha/QhvzZd
5RiY8T26Y5vOoQyCrCIFrp9X4hpM/RSH0sacyrrjxP5G6BTsbbmdoPMpPFnjWrC2
1r7wZx6ishqPSjSVIOP6gs2T0ZtWKX+wVlrWUr1lDAckva1o1Uf7gEbrmHngk8Vt
e+FKeNTZpI038Vsesxse8g+eQgR7b+8rc/KzHlQhmgn+Q46yNTTGfY77HBG7HIye
m48m76igjOzi/OR0aQZBUsF159jmacC/TjWNN5CqE8aLA7fywnSk4KaNaXsjyDyc
vCYIaEmg7ccuCEFCBdAcNvWKaYTmBdGb9QapeHDHB+gvLuiGY0bHlFN0YpihvVEQ
UsxFZJAWq+tLSdQ9Eqn71xIYESh+2iONzO1LWeWVXBqSlkJZ4G6/3IVbttvejZw8
rgFg1A+JVQMYCPPWIRktJrsVjrI+gy14TqAsr3c7UBq1Q3X/NNQFSj8gdKQCqF7C
Rxkjs2//aHFJqULQtCCa7IyLhZkIrKROuanVVvx4K/1C6SGcblDS7Vn3VgRGXDRM
/n9xYY3RxpNjn+aGdBdDf3+0NMYwRE/lOOCpQbW1qLvauinJ8c8nNcEv0KLenYdD
P5iqN71vnbfSPT5lRPGxxuxcjj9ewL+y/2ojjCSxYrU+Ad1mE6D2wc4xBaxPMEUQ
KWbogz4J1RZGFxIojrr+LBUjDB7zcRwe5xhpYgKivHirsRQA3ePoGn5v7kvbnOnf
Htox348aXzgkoi9mooWr9FqeDW263kMT7AT0r2LRsXMECm5iFsIQkcNX/mPAKpQN
4alki1Bi4yKnKqlYnJ3VUaxb0ucE9BON734X7+KB08FUq9QCrA74LEWx6dyIBivP
aq8ueeqWjkwTxlEaKHAwHJdOTYfSnbV8vIsLN2RAjMgZ4wAc8jeWhKaWNHTsER0E
ndwlF3K6aElYQxBCpvvz203jjhH1FMZXj039kjVjrFUcMJ0Jgk2daedwO9DbUnu/
UaWynDep83w+GFthl5r/qhmreLbdguo/lpAUtZ1AUoeS9kDV/48Nsgs/9fp9ZYKx
SHbEI99ENtpgADMHbtA0nr5NX9g/P9qSiCeDbDoompbN4HFZNT1pnWEDazAstfIS
l8IjCwYXsnNeiH9NKWR+xtI+vE0eryURZBEhOmkY4RlWanrGXEHFd3U3eYlXRxTX
ceDkh9QBxww53rYHtfSx1wO4nsLY3g+J6J4Arn/di3pnrJ9C5YDKgZcCV9SEpXQe
YuGyITpA2voyKln3qwMEFQLl53WT8O9lJ0yBpP1WN94rC6H9UUm1Oe0qcLI/ch5S
jJxognCiF/r0lQbrT3VrfEqf7w7HpOA84e9tAjcOmM8h+XSx860qhpd3XMSGQRnE
ucbXVwy+J5zvoEnBnCXbrinpg0dSqiciCT99XC3foAI7CDEbf4vvo/jhH4rErZGD
L0oNzz+eHx4GodEGd/HPKwNWsAChmjqi0AzCPonBvBgIfBYfDRnAPoEXTaxGxUk3
dQZSXzHGOpiTT+T0tUk5h5jL3AislPq1u+Y1i6ZPoH5F7rm5J+LKCnbE2DBAKayc
3+aR8tAjkC9rPf2Z23BzhZB4MiKFvoXg/DL83Desw2/WoQ0ZC8JXs+KnoMb12KeV
obS0QA/piw6otjrPZtTPyEDHE4VgBAEu0u6c4gTJBvSivSekQnY6wdwJZDOH7TlT
lRFTchS9/+NePwaWsYS+9hinlwg5gQ6A7Rq5RGqH3m+/MimbnmAj2cPLBJMNXnAc
9GgGHI9UYGKRcN8+SgqfJm5uJowIAfB1OlvIuVhlnYhueZQ8a3ZXcMTY1qlPI97T
cPTmIItcXHGH8yjhLkvmnwD1QBu9k7ahy36ZvPWg/YYWbz1U2QYfGLBI1Z3n80lQ
ElXobSs4kjHMxysYSwOOOLGw9o8mMUDMSEZRuYqzY70rw1Rk35FXmiy5a64a6cpw
+kZ27VHlfqg7dvvYnKCuUuBuGp3ovOWdNKTfqqvFi4NP/Ok2NwFGz4LE2+1bqvPK
KMP895A0HMVQlI/oaLZj7XKkmUCvcn6y0LdTzsy6U94+T4X+Wb5u4WunVQZHygm9
iKAcXcaMzUMca9DAUxabzi5N76ReocdXMGPaj19bfMDGz9yMnWxSKKoJwcw8oGk7
KQmYJJWdrk4blsJj/7o0y6beRbU/mQmLVvpM58XBQjkwVyO8Tp3nqcROnn5MbOsK
BI7nYZBN/XNWwfdalw6adms2zj77RHuJfl/LQKZkH+P7GhDbayg9j9X8WPifUQaF
EE7pHVmGLwanMO/tyXSUe+ghuxVsDg1tglpeSvXSzxUOZb8lBl7dQH8jAgnwNBqL
hOlxea3JOOSvo27N9KuxDNL+oMKVdbsvg2qjEFv7fiBmO9Vjp0Ab854DC8osmx+n
fEkYj7vRPe1cyUwmoRO4PufKRoI2/BpgOKU/lYvNBPFDUp2vLKiQXXI/famlAA6n
ha4sHtcRZbI6/wuBVmsEYqC2ko+ou/pMjgxfUqCpwow4jpzy39cjvm63H4SBHZ2C
fKwRBvTIklof0G8pBozCfn9dCKv4dZBWBKv9zUWfuBqzc0YH+dB3oMqw+H857cOE
rdJQTqpCiWFBioCwMCprL4ZwWE0ooXglOfqNELzV11en6fLJCFlQAIAsdwns2uu9
xjxxV0rHSlcq3PrvcBjgN+qY/DE1BaGKEV6pDy8FAyQcKoMpbSPDiqRE6OX7Z+UQ
jzdeyMYqLJBPub1irQPZR6GnKzBDndDjppanHcdfwoooNxUON5e8fcSY50t1vIe4
3juSwdfDKKRgSCefE10o6ZOh70IRIdgoCxjpToF/mguYePChNiqyrF/b6i6vPwDp
76J8C8RmO3R7Qr8kkHJdyCx7W2CGynTq4SDPkdJLEI/DwQExIp/xLCisaiKXScUc
dUEj0skBaElhpE4z2YIYDGjcBJx/i1nKTGHQHbwzbmjkvVXJZ0rn72BZpCKpBygK
10SD+5Gecj5qlncpYGzQqBbEHrDdQwn+AX45D/8rpNn4L/4HOhL3kypgwyLed9yV
06d6pkbiPOR8iY1r9n1UYV8oVGuRE2y6pK7yuQ8ojZvn7DoTAbmEd5pDlfo1FraT
6C0sTz+nm22ZO3Po8LFTRUKrcHt/e2cn9c6c9bI8lOJMBGwjU3mPLF+xKqJKSy0Y
SX4DI2drQdDGGdyLHlS8oo7+CIc32DzkFIijYkgvrp9Q0XNAVeRLTXQIdgKHiUmZ
EZLAwc//LkUk9022+Vd3lEqMgCI3nUo9qFnrnAisQO+4hN0F4V3GAqNlIdIV6ult
6pgRI3OqpO/rMuFaeoHvSh3OAmXD2HQ4425gOnYCmknGD8wW3U/6hCU+XNe8WfFR
YaxDgHwl5pR36fCtT7g409LeYuTgNC8WjaYIGmyOyOrJR2sytpqfsD1aEjtymBEX
kxcBMn/TPKvUBX08nmbM3KDfTLpYYlW4bJ5IQ7EgLfRM6TY2gVWzm5GINm7aR8eb
nua/6SQDqcs3r4JYHz0PGUpGIwESY4duzSNGGwF0GDjeKyEAoi1tZtWsyGY2wTxI
YFlAA8HUWmpjvOjYncoeCuS1UsY8Id2EvMEmjPJd96pWm4HnYNFHCZhNX/WyI9x9
4/uhVwGkEuNMlMa7X2fMSb3f4p5YnoB8duLYWvcYa9bWswwCLPo++Dqt9PkAcNJh
i6F0Q2eONaBmocnzPsdmmJhNuD+4zTAUor3a5Lh8DyrZUxMIoY64bHVgRRorEiUN
QZFqEShFC2rECPgbQvtsbc8Q0XkNjhI6xKaxEel4dIwZzBMOWgWBMuI6jSd/sFnp
g3goDW3Av8kix9LYNHSE5NbfAVc+5KvW27739LGlDhJht3ADZkBAZAbnbMPk4Sth
VxFrZTNjqzX2noyVho29krMpVfN/zId0soJ8j7Wv6RxJUvzIO8yxlRbQdytfsiRT
15Mk9HhgX2L4q6PfxC3I5w9TjzQrRP4Q3o5+fiEPRzhFyX0f8/44d5xP+N4ianb5
HAJ/q+uFYm8gQXXfWhVpyysqetVcE8dAFZroWHYXHgQewbi+5flQoY+2wh8Qv3/U
Ocap6W/+sADTnT+5aMoArEIuHpQtyWaX+go2mt3CN5IKsuBnYMGkqYGEbkiUdtp6
BOiKdiYkrrKUP09scC1hr4vW1kT5njY8Cpfc9x2M/aJAADiCSlH3E5Jv0BC83MTU
YUCZ6zqXwiU4ngtgiC/vJQRi8E0WxRXJbNxoPIUCMXfzyiqRecz6/9DIsS5jWwmQ
L7JUmaankTc1/Bp3toLSWYnWzMUWDE6ypjAX3HUtfyLdht5C2887LwZmPBHv8qDK
y9yg/+SzoKDjR9bhwzMccEmY9WtdT2wDKZDh1uxJWakspel0wx/EesoJpLozpGh4
+Co94mRMIdFtPsL/hwoDUv4sXb7EA8WO5uTabJ051yAp0CUy1lMNouXjR9p6koFV
kEgGLn8ABC7N2akTO/1eR5z6q1wqXiuV+QJrJKb9R80mlSE7BUHGGw3BWe0rA1jV
WQzR24Gh/bonxWMlEZqNqqY21RF+vUeEC5lA1x8gvPc0yHMst/zzO7ihWJwFL+zx
AnyUXyDrpaKg0LnFuYede6oWcfmY0z7nOHkBgiy9CPxuRr0b5cLHhbTc7WpLPvRc
Iu2BRjlDPj7bvPYPiCQ6zOB9oUKsxC8SQt5NKxo3CkFKQ7/EFeSm9oaFIlj8zop8
zd18ESislaWbfzolfWPH1TfFh4Yc66riBjPAme8HeIlTtS5KlMTpZAYSiqz6CaNV
1Q48mAceCDK+lhR6jhFQt/wyN/CHL0iqWqdq0hj5SiAeGpdf8DMYQTiPv9Tyk0q7
nS578XrFt+955DVCpc0LfOmA22NWZkmiPiIzdzmAJZwpmX1wxe7cNtPsvsI7adpu
UT1nDG2UtkuVY4aIZZTObRu1cZnKU+uxM01dVrNpS4kgMdcmzDT1yzSByeRptmKq
pkA/ahEMxBFSRq5zgoHNNCZD6RSSKHzph10ou4cDdT0M4HDZfZ6uwXEIFqevFTTV
Y6lFImN0PrwjEHawGObjY6tdE7Z1gVj145GhyIoLL201VDdaG1NJEi757JDlyzHf
itVpIHUelV5dHizPrhtl+7k/pHiZulvimJM/gApvl48sdtROGGWTJGUjByv+Na8s
3VouaaZxLgJl1OQwQKnFT8WsXi6jb82plmYmNHeVJGB4rs975TtxoWombiBw8e5C
HRZFZf9ZNrjf1aYVrR/TDJN34O0iS6BV1u2Xs/yOrRSu2gR0oGWG2QUbF5l+vZDE
auGQTdnD3VFBlhfqFncOgT4rf2/37EcPI//zicy6N97JF3saFyNYfAPUhBeP3u1j
eHugQ8m21PdZO/SHOVTzhkVnxNwP8MsReahasgzbMZMbsj4f6N1fDsXvxWjdWIjL
xcy9iQ1sK21pL17ya90EEURvzGiK5ztfvMOCIenaF8BQ6C/4bXG3d5G6ykrddFI0
NjN11Wkj0fU9lII73UkYYTNw4WU2Eys9/hUZk8qzeB6U9WCcYiaB7EdbapQvgMAz
B8OmRJg6TvnWv9tj1yTH/hWxpcxPLpoUBBtNpTOcoVHTUMZUYYDzN0GUai4tsJNu
ZQe/BnI1e8ncAahtE99279neo279j2ftgWSevJP/KSXI8IPPZPtW7ElRvd74RB9Y
65+h7NvDfAQ1e5n4IIlwgcBw1QGOwaoGqyCzc3TBp92+0Hv8ez3d5whZlXnWr9dI
gWEcVlESHMf2VgUDo/L7v0YUF28LENpYbGoprtV+0lIH2nJH0Z+yu4tUpuss2ueo
V/MPO9I6Bc5KfcWx10upl1bwqdWmHADZfyj6u0kHRmiDurbR9reAvge3/EoIsJua
wJ7SaM+Qvq4/Wda+kOu8LaMq941BXommU0upveJSPhAwnOFelYbcN/gViBakun/u
y1bZ4a63cMkYN/D1LKRSTC35XX3Ur505g5Gd/oRW6ovEhdCWDkB1tr+c6DBU/bR+
c6UAIBn0xF1/cq9xT8HjmOvPHb2HOeMXexovzu2Pi7pwUGPxN5ZE99e7Qoxd/ATc
QgbkEocgcXeqRXQy0rlzz4kV+XtwSKr4OCbl8hQZnwEuyN/LdN71KGSBHRttxFjn
vcA1z/ROmTJDXqe2FeyVd9IZQMRkY5uytwnmzOWJsZZbawfzVbqWgptZMXPCDDlQ
yTDoKzDfboHGVcpwlyFUrQmsPokP6+1owx1TeuehxnZ2PSbG4tiA7/bFSdJeJuYB
Po+R7iIufHkeh/x7QCCgFLcdSL64h7mYkbWt+/j+nosFaWY6bEWQxG/H0mh+sl3r
5jqjxiRHX0fKSmG/DmUEKv98BEe+ODJDowTJddYvqbUVfUs3fzs4tdxBn2VSbMkO
AGkBVVJuXORmFFJ8aFr1xNajxodsT/a12OQe9Q9ctgSaI/IZr5qsS4981BbAXKqp
M/sKNt9S+tymYWATE3yeo6FMLfGF184rlxBwdylCbjlcAmiJK2kEEImdSG68eGZz
plhEcsjlD2FotAhUzYTM7eB5TchjldHJTNBirDqG7Ukyb7XRWg5IF1KfHYLqtdcM
Fp0+tjzFtJHo4xZO1HUUiPofOXmk6lhBNG6IQOlu6cEr186UlCbnbO+N2j37ub9s
zjB7Mt94qvmbgKTcsYSaJYv7PBMl3P1Q1PQJ+CA84XGkxt8KPObqt+vgWTthChl0
qMQ3MF8x5z+n+Ii5Qie/ON2ynFb+amuRoEl+Vnpj/SveYAU3FL6C71yzBFa24gjK
/Fvn8tmyADIH+5KtGrs6JJI4gz3Pwar0W2NVEhYk5m2pn0Z6URjmhMsYZ1WGTsUY
eZ4fLfDCA5kbh97/84coq6puRhDVERxilCZsqP/LTzT9BiILPawCqYijf9Kvt7OP
+m6mZMkgM0Ss+f3GxlLTErwML8DvxU+szYssLokGoBHStDxt31PP+UjgZXaPWyyt
sI05g6/JvN6FmmeWbk4bcvuoGGPY4z+WjWkkcz9r5fGpm0pNVEJUEpG9lCt5vV4P
9jBnArEQbJpSJ+b0XMKaR2RK+yBrURDxw3ihrDgutzRqQulWdBgzWEnMib/ILio0
iDKAgI9Zwx4KdDaG4vQo6szUBSFYqXEAQsW4hUH9f+MMSj0bLapV9hizM3Tkckld
OXzKApNtGwzQ6ecdiWCs70Lk/85UyIiysziEZzo3H+pQiNn0PrDUh0OKjW2G6dlE
vd3zGkTcEcGbdl7/GX4x6asDMTpUvKI16/bWle5LIVdp9ECO6b0U97ESdYIHog91
QBdf2PbTtzZzBFGgF4HKaEDzDcR6JIP/9gh2mg9B46Gq4KjA6GLPM6MzbXe4G2kX
/KTMRP0FtIt2wyl1JgsAp1ZMfak1ErEU/RgGpT/W+leMIXJ3EbHz2DeTGe4n3i9A
T0xK/gJv46zryo8FG8eMOIC+Z339LZQ6HWLndb7dt9OcXasHsv95WHJNi90Dy+cj
oHD63yfO+GPhRqBXNbufv5mQ0764mdcy+tBYxZDQ76AWxYB8EUROU822A5YXi5Zf
+jm4gisMlo9Kz4ZLMVMdXeA0LA5CRadwGBRCY+4w0oUfcvoC/NcN4yiY5kr50252
B4J9v+5iqW/xpWXux+lByyubNBG+j2mqRcRBTYlgbMGB7tGX5nWxdRM0RJ3mV9ki
koRQpo+tu/nVMVkr33YPVzINMmVTXhrFF1LJiyFkuwehconYV8ebMbfVpyFOM8DX
fX7V8nte+rPfu2r00gOPmbeeTU9P7znBNB0Gb+zqrSyp807Y8vc22F7Al1TicEbu
S9S2kS24XJiAlQFwryjRbljcVRAKv51V2ia3cngS8XakeWBTbg6OrOVp4AnHPH3i
AzZyku6CwFdmvu6uN+EXwsoeWvhkRwNw8HoLuRA/GGAvAnkesPFkkNHEVT9gUlaZ
BAyXdz61d17VGwKL/7LJjq35bvTUBlvw9TUApW12DeVxf8rPzz41Qr305I+iHg2D
aG3YXIP7m3TMCuduHSOAlp1lDaWtKX62MwTPTgUVtwgDUM+WQ7DvXKfdaHTP+3pj
DnE2hOhibpPtUY4eZkivYY9I3htwHLl0dT2Q2TNdJGDCn7F3X4G5NM4hispBvpJu
XokIP6Ud6eVTuiDOhMMzY4ei8X8TSrR84+Opy4dqvOlF/2eeaLu/T2Row1slhAdF
uGK+eqC7CWStGh7bEHE1L9YD4WHgELpN+NJ2tNuMpFciue+lo9t1qzJxrbuuwub8
GnWBIe8+gigHqrGIRAzWSzVzXPsAdDAkrFzCQRdhGRQ5D5WBNTc3EmDONeBwJHuh
2UDMqeIzhYSLdzI2x179bWbfgFWeB4Aw5J0MS9o0DIaGqa8GspOlS3Bme/ZWXhtB
wCVqE32xC3UDncNMxyXp3w7Go5wzwd47P/YqXoHge6L8omFyYzri+0kfif9hQauA
sRXJDS1/lznjGODl3+2uj0DZSs1ZvQqldACq9XnsEc3FqCx30DuukdPY2/LJAkrY
F1Y0uloGIUiikHyqlEvvrJ41ICJFrCuTLmfTSzF4uLIfH1tmcT5YSNMy27LPDyjJ
E+BBPt4y984cJeMmF/6iZGVGFV43vAtNvzhDzqB7eJ2rZgfPN/mk1RUXew6z3/FH
Yh7UFJx6boprdMT4DEF4b5TJse8kzQXooYmdquUmxyPsJ4ZoYFe6FmJgPpilH2Of
0QJCQ5JdZcFEG7RbQCb8wzkxnPkeXKmgknXyNyVH1lXtoRHVm68ONpX+/rATLRKQ
SYOghVt56QrRaFovSAPFaZicg+oidCVwsRlkpp1o2bD+6AiIcjF7FbtjRkv2AxKr
pkW3wSo2SZBzjUmdsohGo+hitDMyTuxHQ0XSBgeIMS8l3Lnw9bmKr7ONUQtkroDk
pzn9ozURx1nTLz0cqh12nrUYcmYGvXn/4z2pIAkauYf7Yj7VGVPuNRr5Z6A60MhD
BrR0W6/8zBprHKf/aFfb0J6BbhlYhR/CWylBeBS/me5ANNwO0gAE7VJAf0iEY3KB
pKtwO6cZrOvRZc9tF33UdSz/BcQ7JAh7BO1cE/dfgBffUvy3uOHMZUgx3yxP0DPf
F56JPMyqLkTJ3VfaNRgW7E8UWwHCHckH36WZlrMRbfUoAEVUEEujdtW4sUci5agZ
8HFrvHmsWB/2Q2S8KmYIlnFGCVIt0pnyHfnbkibTwCO/GLW3au4lcL6e0qfs/Tw8
O06750Hg3h2aXp492A5II0Gy0DDc/Ku7lWk9+SSrcpNR/aTsOvP230BNX+vYFZUo
2g6hlgOHhHjn5RcJPMtMyEkXQ8IOfRrjhAezbjy95B33IS4E1P2tksdMWoWG5Nqk
yWkj6weTuTBG2q30jzruG8xrDGIoRyLmsVhR7VOW+1GrZoDCyIt1PPSvPLalMObb
DSN3j09WVzcmOw3dA+uhqcZ71HtsyOP9QEaDbze3uw0hD+FMyHHsITnjJ/45AZqy
kUAvw6o0DHLclPNmYEIRR5AUSpO2B9BQ2IBFdJTviQuBweyy1foz6XVtYov+sFXR
j0hHJq6AcrcNChBAyb6Qaz9qmtfamIXk25/lYg5raoLwDmfcafU8yBrHXM3Bjqjj
uN9i6Dxw2WO11fkKanrH2/r8R69ug6nzWdFXw/6sNMdGnW0S34HdVorgMBeRKlQf
Iab/TnINYGgatJX/pySjFxJQ9ZGzqEMK5tptECPN53dpnjYv7KNZFxfR6yZ7nY+q
AJFn6rzCkuuNhFkwfVwOcrLlI95YRwJ8u5fn7Uz5geq4nEcxYINVMEir6qUXyiXW
AvHk+1avt5HxObkPnoTs5V5soQBiOs84413I4ysWOCYmwuqSZa4gt35B9+Nt111k
sgQIJSaU1M1G8vPu/iONFDCDCs1gGLt5SnXG2dGRAw+6X+TY7rMwEBUowHDlCaCT
g3pD5ru/OrGkAWT58Y1dKUWPDZ0xgLqJF5+jd1hOPGqxEJD69MPKyiBAZlPuSc53
oDxANNVUFeEDmN2CH1ho3onsQx5/TQaoNodi1ZxNrqZIO6xOuYX5HwO0UFsl9NWQ
8Om7w8uJKeK1GJNJT0H+vJEIg/WW8UOWKg49WXFtd1odbciIbcpPWtBx+gwW0OAd
NEliBf+g4o8/sbl/cpP09g4SOaErNJp5I6+pYwo0yitO9aa9vdDj9l8GFSUFH0qN
/QqsfFQKpdoQa+RvmeVohz76yJYkqQ/LqzSJFZNTn64oEGXtgOY0ssjxFE9lNLUm
dik/BeqJjL/KmS3tEVXud+VXoj58svhgwAnPACmFQFRNBeTB5vvn7CqiSib6tEA9
y/GRHaZtNLf6/v3prk/0SlBcPrhBt+bIMXFzPsrsiOD6EKrSJT2Wia3j16Zv2lMs
ih6NEx+iAr06W6ucEFBvNgLMVQogWYTma7nKghilv7TPsQdQ4rWGN1jWlAKMxdIK
Gpqkb/t8aCZWWsvLLISwNN4RRyLSGgT/lgqRk1BDsFRawxhwai8faVv/Vsdcku6n
9RVeRgzQNKS+/lped1/wIxrA73AF41Ai6Z9oQ/TPMOyadDAssxN72UI5wBI9dfq/
WTGI6uvLFXqLbdfxT5IB2vCcDUDuQPySrpt0AQAtQYhpSjAYajaopoi0WBSIeKC+
s9Vu0RUKd/mjO/oyKEOXNxxXG4fa9jMEBQrNmYBIlCD63+WxP8G/IR3oR6Wv/VbQ
B5SmQOndtT7wx22K4Oc/FC67ZGTff7A64zc5EmT+es5ERQX/E/B2M7Q6/IONPJk9
YegAsbSycGOv+Klq2IF6CfBairIdfuq9eXhyvUTbHCjpTHzFyBFPjMNt37e+dUaw
4KQT5yoxM8nZTz2AdiEYIGGgr9oq5HzOJv6BAfPs9pEvYSsTKbuCsQKgJIPqtAWZ
Q3GwEKCpWNw0Qzyv3/qxZbLBjPJr7VN3jtUXfx3qH4SZV2l1vUTCfV/noBzdmWxo
hcqMyWlT0v8y7Yp6RfqWZXlpaAstX3TCmCO8izpsUj2CMARqIG7Djy7v1iytQSAP
sYtHz1RhynUwUxQEraJC++e9aTqkjs2ZN9EdStWD/z+yWkrT5+Rub2ZOl5fB8zNO
5bae9AHWs00vj3qrekpcGLQHoayFPtTX6bwGzHM/6UPJBwcOVY2vrFrI4iZta4sq
DsdgekjsCWdwjPHs9HE1chQkTLSROZOOUv4Qone8ClbsyyovdNrBjjglKJZtCw5g
6xvnvDwxYt+aJhTJTsFLVR0/PpalPy3eVplwkMCG8upiGlhEMIwHLoYDhQK9PqHs
hSc7OqOdZLsfKj23UH8NH2AEiZ0zDhjwe7HDWWC39CJgDMInDk3Fx+nV8grbBigf
J7xZvA5h5e5jiw5bdvbtsK4O3EEpuc0+F+EjNxWK2IRePBAMvBtpGbHYuBv6YcTQ
7pVhQVBpBwutMdGfkReXG33m5C9n4boedsG1s/JFQKMCd3SYEAHYi3h5QKPY+8fE
Dm6eoeFyzZb4tYAYXYgip3jNCYTeDw+oyUhkSUyQMjoGQMpsbVxKoTlFn1ODgwP0
SC7ghIqQE6CZLXsZv/30+oAA1HsCR/uqvDeHTDbh5LcRPgC7edjE7viBDV56TVg6
LQixzn7zY4i07qr2/yR+9EG26KdOUt5L/OOD+kIolwg+SRBTp0WeLYHUH5H5eNZm
AELNEIxolRShwsroxRHbG7P991u5PQlF3MN6VIMZSOIq1ZppLOF99zai9R4oH8yG
/wR39NOtgy6rgHYT+Sz+p7LDwtFT5fkqIgdCkBKIjVd7JkeJ9hTqh/ldXsEhpGYK
yhyswW5XZXlfecCGoD5X81QW0JIRLt0sZe+fNXhA7MDcziy+WDpymmrj9PKBWJGr
Z8UFk7kt8CeGQQtDaZVseIhIIBeXhJKXqCvanF9klPo4HCKEDdzWkbQ3MFtBxKvT
uwioy8wdcUFdV70dQHuqmLsYV8E4ubXnm0Tk/2VgAjbUuIXJWXujR4tyCOzL8dlb
jZ8zGUlWLllX7CpW1CliMWMu+9btOB4uQjkaHTJwtDHknZ8TR7LvHoRQ+vPpLZVV
jekO6a5x1wu8EsjGMoulWvDRSVrchB74dm5sG0O5X87PtVFgl8Mov2aZy8VIrzId
yl0aeQBV2lUFGspCtde+P7yZgDv42K6ZMvWA2nwClYxzGjSx4iuBklr0pr4BgV4I
VXbB52o+4vQfnJbWVnOPNjuF+1unFWjhMJunU8AGvGXRoY5uShrzX4k3kcRabXaR
sJWVWcfZUbKGmVkJzVLCRvwkjVLnkbfUmokMKM8QQ3oVJ6FZTJeqDLZRXzZvc6uK
5sTmu4a8CTSntKXlC508mURFlZs6i4DYC83+0gEj+9oG4IHBzNmI/zjS2sW01wRf
`protect END_PROTECTED
