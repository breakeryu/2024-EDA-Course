`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TrsbQoWkadyQby1kpQ36SOYw5FPl6D+YEAQXnqGM3oFlRVExbe8M9bFD4/tvFl6c
jTy1XYxfRu0zfKMKNAZPHdaF6+uo88IQGI+q+lD1s46H7+gpz23qOf0lobe9KskJ
n34Kh0mPRVtlr/hcxinBAqWHbOYgyBb17Jjy0hLjKNjYqeJkTfDPqFq+HcQD/KNu
PpR1cbRT2cZgPxoF7VqJEiUSSmYC/cE2Wvfab6c7c/moGdj3Yno/ZS6QmoSR259M
bGH2NQREiXm7FAVPDg+9NrIxsYwOsWbg+LL8baZ3isKxIYnix7/f/N6AHODFfz9G
8lUvh3Q07r71J6L3KBAjA9ax53eEenRL697YsVjBLJQ4iimupITKQAOBpJ+4gOi7
xqlD25Suu7Tqjqs3wRaLqQbiKQPCnXpdM7duJ//BHYDUiovDiGr06/coR1Gf5YsE
KPe/7+yfycQzM6OIn6GiDciew5JA2ib1/Uo1ciTzQGB0k5lhnBAWtVtp2cM4S8GY
4GDvM2lfU3IfadrzqQlV633b6ZP0rzQMHgw0qEFZoveCEE5Wfw+AYjfvqORdM/g7
rSAoemoKcD/UkdrKVf8t5r6SmnA1KbxDq4YHspgEW7kK9vGlLRFbmRBFOT5WmYLa
wCCB8jSg+YVNsxqvwC4gxzoj/vLTZJYKB9S+ZEkV8wBvQdaxZidhkAFFcmr5IASb
5nuRDqZWjkHPZygeK5Wj1tIcWPiHS5EYnI0iOQqBu7MZmPfXmaJzLu0Bocsxga3D
PjP1Dh6JxqpeIBCKUmJekvEoj6hoB8aVLawlxEkezZBsXtddCYwMuoKimN2FmzJ5
7U4udmzoJE/qGgxxAQumazCD6KbPsg+OBiK2LFULL+lQXh0Jycve+zlwkk1L5E+g
5J72ZBpekZ/T7FULdyORi7U6URtij/8i+3NepOf17S3x0VEaB7cxmP37N68j61IW
bSo7Exp1xCPmp2Vj7bxf0DrZ0OP+rxjuZg6Gj5u2WVUMG0zxpG6jMu4WF6PSA3a7
ZwWgmR1okVvKFWB1jgwFS0IU0dxFqkfdsFQysglxDppUVxVO4XnUYdBkuUZCENz1
qkQBCp05VRpFz54rLgs4B/Qol1FLcSMKs0R0MMNnUObMpg2xbigFlqNyf/10Jwrw
C3LZcMfIadvmhXM1yN8c5pdVZsfnZ14zC/PDpcoBLX4mLS64nkPjeI1KpUtfohOd
Rw1rGchnKbtT17im/hHG/CnWCJfzDXS1A5DTBmncOm2Ig04g/sNPLJPgERkjsPjF
LZk+I9XSI5eQXt2J+uhLkQJVr5SpZ8dkEQqd2bJSp32czeGwv/ulmX/CrxeqiclJ
GEgvpfG7m3anrwjg/jY+j3SJadSdGEV6uSPofw8r+xn/YfDI3318Ljs4tfQEfU85
ZirIXseyfq/9iCEBZhWKfzWLhfEwYtSrBa0611dclPOp/19hsEz8UlTmGNrt7pCO
xIfZl7idGop+7XGLCwqkh5p4OadkRdtwpLV+4p4KJyEtn722Y/iR/VpeZkOOBR5U
i+voPjnywc8LJhcAq2BA13sEAJxSMCzHgHIq19CRKzT4OiPpLM2gytdcCE57FeR+
f7LxvAc7bRZfc3SrceGHMBXKjAEZb8EOSm9pAq0DrKVQRKCPpzFFw7OEOzfiiemr
I9PXXL8Ntjrj/mWBeXCzSDJlhY6l+4ruxlre+WYjhqCUwvyi++7OqSxTFjddfMLD
CvjTRKC8SB4WJxfgEBP5yAhgtVIpyEMADZY6w/C3BE7dCPFkhT7ryM03WSYk4ENf
wtkabCcJiHYCNf9W3CBAW0vJ9XwFd9EqoZSgotH8P7i4RdstM5JferboKQZgW0em
/Ruv5b8YCYhK7K3Er2AJYHNYQe+mX5qAeyJwY9BKPodDWjOJ8AIi/0P4PzXtztI2
glY0VpM9K6XScT8qTBH+2XVW1YMBN6A0DTqVav+3nk4kZMeBoPQi0cIw+f4MPYfZ
eDW6Kzf1iIt/ZULi+Q2x8J3GP4B0gL+m0LgjbKsWP+5hQCR2SPMyqpHeGMglla46
opasBMW2JsgFrZmFNG6S3gHUbA1ajBagBB1nEV3FwvWzKsVl/umAfpGekcAnZrCS
Xo2wiGqD7W4/+IhYHLMZfmDQtHJtPOZ1OSCl7aIyk/dc7JhzWhiWTcHEnV7TA3Lt
yr6anlzLERhfUFaFx4DIwu6KbqG8XV4J4KaA73Mj3JiYKRamYvULuzeWjIp+BA73
H1mSSyixPRUAvyzg40igsgF7+77dRLdwQbsYvZ+6K0Hh/U6rsZ6YmsaKmTTenpLi
5I4W2sI9O5odPzKGaBpnhurH2YgF/9DSozPZxnTBXE+TU39KViKxM89cBzeBDdT4
GYG1AamDkA8RcTp8NpWULWWMYaPuyQiKkcX4rF9IIuUZcXy4MCFashbgonCNbb8y
8Pssojl0hR0M9kEviMdEAmKkOb/1ZiTKuQon6ZIhw0WeKOBbtzAC+8VRccU8eGaG
/Mr6V6AR2Ld0yHTgwCV4RB8PK32QgPUuWAjm8FmLeYtQ57VKYFaYvUy3HLuIMIAN
Sul5Url65oAGbldt2PNLck2+MWiVEPRmWjBTw1UrymNMs+KodELiQHMiE0rddjAM
PBcw9mvHHyj7QQbB3Yp7PWpzCKPzexXbBlPnDTEKUI+XHRZdCc33fHxkbXZw1RtX
MRdVYQ3vs1REVAsQ7Tdtfubie7hBUeCPtzJeTCirQTSK/T3lGN5QYj3MGf/hNTdW
bcQCQ9zauSVia3dGAQgNpPhGAIzt4sOgvvbfb7EKMSgzUMjMk+gAALZ+4RskBwqQ
DxiiJuu6CaWamUCwFBe7HCaFr09PVbAsaOfCrDWSLxDnantxZBjd0VXDwyLoUIdA
nzslncFW6Qp4r24tIN9A1UFH7u0C5ZAGUE6xSWjcO04mzAaMd2maG7pnR1jX69fe
xbXUMJvSqnSA4amDyrh3tDfQ7mKaxcqahZ9Hevb5bIQaTApzbfFdJF6rMrZ0Kg6Q
Cts21BHnicVAkW083W6JAcFuywQw4+NU6BGd5v7BmqagXo5EKlaSM9+L5TxvTUbb
DoTFxgRE/pTY2PDCxKFhtRyqTlGQlPZLxfSBzRnkHoPxCcyoJ057wGMxLTVuEYxB
FDBbFuwF7ZZIk36qA4J4AroFg/ACpJeBP5QmgOzXhFv6ZXV+A+PtcWtrMB1zBzre
GME/IrEU3b2rjv20UJ9pO3fprsnQ/dvIooKFBvjcjeNJFj6ZP9lvqWaie4dCN9tC
Rz/xJkPSpewAl8JMfcWg5m1KRtZ/IPqvF30uhLJ8o0HxNov7uXG1mxASfE8WiYCp
akrVH1FRAx2c+j01JDmbDeIJ7IE5vC7sqB8Y4OgJq7U7n/zaFNbtgX8Pi7xmZ/jN
c60JWA5RJD7smXu6BfCNT6dlEfq4YTJW8z+qXKkqE5ueXHURt/Y1Kq4W7sXpG164
3QiYy9uCe5CgHcXWBNbYoXiR9q4G+siTplke660NpPwxV7fkWB96srj2CQ2hIxBL
2nQHlhpXUTjOTjyCcxEJjl5rWdOob/20sFIYudyHvHscSdSs5q3DnIjoc7TuMGBs
8PlJl/lrpV2FpTjW6Z9G/vVixuvb9A42Ks5tYnAJ8jTygp/slXC5vp29crQ2kkd7
33Y8xhjC3Ckiuqe+VHrIi8ljz71a5skiapNwVlHa6yxHsPjwwo4kz6QkV57/VQQp
CpRN6TbDaO0FegqeoZ8jWA==
`protect END_PROTECTED
