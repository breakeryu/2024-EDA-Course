`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/TE7DBrE3vVoy2jB9Aam2bltpoPPBd7viV0alfYiVPhXrLLpSBIGDV6wX+eOV03
zrLoJBvtM2W1XpkT1FGqhNiZZHVFLQyc1MBH06BXid+/JcRb8XFcq4YGugKfPoTJ
avkQcW2XY4EvmAy8i9HEu4ku6wgykGv9Q72tEE/vx3+CWmOoNsKE+0DlmhWuX1Jo
L1c6A6BpZo9e1zHYFPlyquzMLDYhfK6S4btLabdgBnEiJni6kxn6LTLqqyKev6yN
q7xrj+jqYMOoFzyUnSQHkBrctLUjZLpo9MEGJQ8M08ISLaLVothsPYEnjiJC8Dtw
7KwVfxpXSKaHj2+PszrJ/ZMf2oYTTxvoe81gAGGB8pRfzfMZJOvtQ/KlU0YOnRV6
20++RzPTrHVXFbj+Cwl7xrLN/Y+K7agFhn44WuvcJAjA6QDvKPcNaZlYPzY7zr+Z
U3y2LZ8K+uYAJqnYdelxk8egfwlCCPvoKf0o82Z3nMXxfbcZBQrFEJw93p/0j7QA
uWs/AWo0XA8ofs+TwOoWUCgh+KJsxjo8+aPabcJPFHaOTcMcKrELIHQG8G7UxUUe
SQYPdtG3+0frqP3vnjGWbe/QSV6Cx9sQIq8t3Hpfq8hBjtDEVNtMHvzB9wnh/dy3
/8L5boNwXm0eb8ZdAB1Z7AAJuWkGDj/ThITUYx8jTSxtRu3J5UlUT6qUWA0yd7P5
twgv5oeTZhtKXzfnQrNEQOEHocXiABHNtVG0rFC+gHAxlpNxGXJn6a1aWyL8IqfO
ePLaDpVThY9H62Fy6Uo3jeK0aGglQEQ2gt76A++xeWo96FHvLbLGYyidCv0EJYTJ
U3V5fZAlQHjM9jy5UfJcKy36kYgTvUwlZIMkg9W1AMxQ5REAQQ5IL2hE3MbaBI6H
nFaSvg63FFCytaXsMRckcH6maTV7SUqsaGufh2wzLXXjUGJa+E/7GfNAN4vuId4P
wAgV2maDNQpwynfV7nQeCzMPfBUivc+AvMr+RxId3mdRxqk9VKDNXpoBiqYiAOUf
4Tc3sVlrg7cNejsD6sJ+5kTOt/BgA6xmd35XTErwkYI6//+eGekhRI3cHXocSz+Y
QkLYczCw6Vc5jXazqjWpopvVzxPIc7U/xoqKjHkYbBIosk9rqIOK2WMpLzKH7vdf
vXCOlnKniAZ7CXMNJP101MpOzcRB+eE9mmBjpopaEk6v77EEe73wwtMrBZ1zQORy
k3t2wqIoZrdyEYEYbneAVTE4nkRZPpfeXM3ya8XXkyPV9Ix2FMR60SMjLGlnNaWT
7Y6kxh5cGn9iI5opk6Pp/93AUTPtxRC30SC0oeTyAbFQe4HFfL8AZKvBsP+WKUyQ
x+hJ5vA3tp54g44ArI9wn6zsAdgAVEm2M7k6nMcBgBkb/sFNGBeIcwSpjcP8IllW
wmUAdLaU5riyCwVIfP8bEUkznTLpeZeKYOUVfNfyxhzpGywCRhCzHZD38Nc+JOGa
VAOcrG9qC5QE6HyyA5lk0bbnw1jRuiirqrhIP9R/3dOS0esSXf/uZEnjv4JTV4RR
M9F0EOeD32GvZ5Me5BsCGm/JUuUSj454oIFqDnbPOOtOIH2tzXxuRqTV2owE7dkJ
y3JKlEz76Hgl/NJCaFHkvBX3YYkT5T40acgpGoBGONwsQfnJg4SVZqk5szjOzlTG
aM46Zo+eAGAaaybqJ8Ra0pOaWqp/s48vOSy0ykABbl9drAeDxCyfxMDnwTIEMCr7
DJonLstlAXBr2vDXu9yvhqkez9tuaKiqnQ2J3ZDrVr3FjPLQ0fazY/JRtKXeB3ya
IgPsZPxMpF70xS0q+urUaE/VITUFu08fg63+61zMezbrDIzWJQu+lexpMKZiWPof
XaMn9itdERuI4g18VDGYmHsEes2mWpEMsMLabmRwzBzGjJUfr4xOCwluL77zCzo8
NjcuRa/gcBIyLrDiRj3KfuTExOZlDegSk6AG/qkb4/3A+ncBVhYhMu8VLC020v1Q
DKRre7lMbguYKTKpd6xabSirvqH460CZ9/prp1jUyYVXhu/XV3QA3rogmjquPxlQ
3EtI/be5LksHnqtXIRKvg6ruUNt34XHIS6qQfNTFRHJGT8pziWqQiSu9uBBchJio
jtjLv5d9O+Sft4+xgYF7yKk2ZhTlpguvbcZa8bS6WqOc6o2WeTnhK5OjPntaqtpH
9YF2FeRuzJSofIwe2JHfDeJADOdOGO1oos9O9KnTBqkSVuIIqbORByvrCvZ0Pu9p
beAf3Gl+x31yjVgE+l4k6UFI+PKHzNVJ2s6Gd8aBHu2GHxvCqmzmmywqK/PGktzF
Y38RzFNZRYnk9WMBNvnKZ2XzUE3HpuCewnTJnQFH/D82W2aB1bXtLFE3mK/tfVoO
3M9XnftND9ZqSWOUvq8+m+nGyKiWLz0Rs8ImjjkdlHxM4T1Z+AkfDO8B89/pWQjK
95C13EWJUgIXmuGr+CTSOdOphMViSyPosP+obGmNxKTBOWfOM3/Iu7i2BCWyIoNL
fUV6tEt1ZUX6C7RUQtCpm0/pdak291CoT7jmHLAlwefuwsNuyVWxb6YdSgUTEd/G
4ci+4+g3Wb/QN0wflkujJuzTR/QmVdwHC25HEdg04DKSe/aIPeySTG6xDDDbULIe
KpvOAaOxg9ElGi2QtaNwV3lJYBl/iSxuVjdmyoW7DLPoByknxFhH1eVoEljVHemU
WpC9APTcyLMud3Lrd5AMDfqwJo+S5zvbE6BUh3zu1+57IgalGM48N2e6XNFB8CBy
a/v9e/jquCG+epa6Wbr0HfUWvW8pTI1aiadyucHXlmddiaeopzNp+2uKz8Kzbd/a
DB4Eh3DSCBegiFXXpOPg2Bo8Jwe4erERa31Ycl54zWD+NX709evBRuEox3I5Ljf7
AbpPnEC7bESI77meOztEJ/Mfu+V9mbzvQ7DQZw3kvsUdJ+a1MHYvfbBsMugws1nt
WTwe72xeSM+VBUd9AaNl7vkwmvVa9ps2579+6Fo/0La9wkM9sYAiBrME2m0LdOXU
thZygZhPzJL3qA0j3hlbNPNqo6B5/EBArWe43xcAqUKgoOyzsHGUw4CKE+XEyi6j
cIh6dS8OMaiJOOsvSoDvoKlUuNt0vL/Vh5duiVgOMkf0EP50lGDtX0In5Yqy3fnI
Ady3nn8sGF9cJq6/x02CURLfDdHmTcJ0aqfWjN/6/paDzuiwUnRsfSNc6E45kbCY
qt9NgaY7eghGLXuK9hWa+FthK8nGS/udriS7LMq5dO2ZNjbZiL8E9vXv97YlHuOV
ztHMUTo335j9cIZHvNxym5IwEy9BDwaSI+uiOBlGoSjbLUVn/mgiIF/inNqlQkGM
QxgS5HV5pcqGtsYBT44sXEJQU9SxnzMGyPDoOZDc8P+RdNGPqB86rBf7ydd9mLGJ
+PHsz8mIoV2DUBHjtVFBEyI9Nc26aMh/+kMNFRx8encrnSkVINq6R7Lw+gXzfRrQ
u3wsZqnwV+oBQ3IbpAkDuHGnTlG4ropo9ivpsL5fgVYhal1fDMIrQt1wcUC6xlSF
FMeCSY7qEn9kvVes4jKGbnOcFLDiRE1gzMftny6UKIlOn29g8aj+y1Pfv2SA6Jc5
ig0qLHT7cr9ff/Sgi+HfvzvgvAzYwYzvnEB6Ki43U+/69Qb+z/s+B7p/eV0l3v18
qyimYqMjOZctr66vGkUZv4auGIo8WyAXvRlx1rheX/fP5JTs+VRj9hvvA6Dw4HxJ
Xy7L03LCBTLGePz/cNtac+KDC6yhtqBaMgz+AUIsvPNfWD6QddJQDoGDqXkaN+mX
4Cs3dwNfKDi6/HStjShagoJQYXYw4swFHawRm/kCFnlQ8/6dEU9CIH1ccC/xfV1+
XoAB0Ah/CmVeQPqJAjn+uN34OcuR22KH3+oUBidKEN5Sv6Gf7P+SDitPR/RUfQhT
MkiIXRgm/WrCItmDt0nzplN89ZO34Ip4Yr2KZNAtKu2EJOouzb61PTbDwubYbz8E
YX5D0j+ueh0B7N5X6yC6PCXDzrebvpXu+P6nNTli+rmMgyTcmWd9ptpRrsnBo9EZ
YJRlPBue1AfzS8hHNl9w/fMIVLAE7JH790BtNIZ1iGIc1sllUiY0vE/cM5pJEMhy
vlBXDDMtbiJmhNnsAEsqwVeRgPM/hV/UwkqrKliFH9Es7yK8BXTPo3U9HhfHkQ06
ocxFFoWbSMjUBMETY+LSa4yC+rfkiaP1hQ2D+MnlN8eH3pKO+gMc5yRwynh7lZOw
v1Erd+TbbBclBgnYPiFtREUTKsM1qXOkzUdLrxQs79K1HePGVl0c0yYSi2XYh+OG
Y+A5qWt0/m1vuKByh0gUETEzpIcqyoB00qN3QxyJZVvQveGcPTsobre+8eUHU2Ex
b+gOHTgLsu/WC4P49W5yVn0FYzs4jpRy7+UkmL7/wtQIy6EulkasdNf/4ePZ30Vq
o4mOSHdyxoddIK4UBW3qmxghwHjhGqETyu2dTmjJL61VyEmOAL8sby6sGqX0i3bf
5uUod9dlZQrj+LFzyhVM7pBpkphTGy1G+VdxhoWb/RNXrG3K3vWJkE5lTlP1EEcj
Q7elIM+PLIcuNTsolYxVxRPaQxtCzHj/vPO5LeU5rIPEs+A9hczYJy2lYFyDoS2C
xSs74ukHJ7rVcyQrkMUgwET8SlUYWrU03aNw3Bdt/9V5bKy08rs5eZnoFzjDM2nC
97hdlDtgLd52Rpjo7oLn/iyFgrD30yCvS7oFSjMJ10oSnUtPwussIqcSE5mDbuC4
IkKtrfAIxjWNSLFY0Sjd5GkScIEBsDuPgDLfr+ce22qjzYSBl2UXoLbGLnBKmCju
6w7FJq+VxbP5K64t/MqpEo53hRgRmlDqN2ZTOScoLF19P4Dxre5AhlAsBOXN0r4T
jkSZ/HnyhMVGQMaRXduQ37FUqM9ikap2PxGFc2y9cT2+zH0zuJZEnh9En9kgQaST
7jXRvjswcoA8p3KSy+TBSEbzv69xHo+z/9sfgGLDfEtOtAtWlMIzLQh9T2BspHpO
SDA/hroEsE18gTxEqKTrJaAKZub1IQznKRh0lho09R9yEMbeIjfjbw8UnRYaRTpT
0E26oqUTA7jMQj/M24xsl2xj//w4+pmL6jL98BymIPWBrmjBAtVl2yAPyQ/IzF1L
d6dX9IQD+dM8eZjMTBj5ZZC+fw3FjspnU0FE3v2u21NjnEYStf+dOJbGWB4HkYJ0
Rgchw36t5WPU23Ibob6xaf6E69mZ3rskxPyq71/wqIBC6ETcVeA8yRgDst2fh1tY
pbnqscej+3AKRUj+6kM+TFtLtiDpFNzi8SXt0J3lgIFkK7koVGXB1X8DWsonfGvu
AqQZgjYkTtT9K6CMa8U3NR220/FqlAg4XC1aW6t9UhjqNfxrGtV2nEQ+9S+jFW+3
cSQYW0tVNd8Bha20dyPrjYrw7yiPkJ+WDOpSr6qnZIvvFKsXow6b4KoN96maQIVU
emtJIXSK/D4hn7FgUH9xOxWWj7dMgvrn06lqnM5noinztEktjnoJ4x9x1gWK2HK2
RIQLz/Lpv2cNmOBoP++7/LaVNx1GdRbcflbMRBJdHvsDsDKvAReanTa/1UxhExjJ
liR5vkWxIfsPYlI9LX+QuQWfRx4y8pXpbLrGml57zYw1teUi/eABaLZlRnp6x6XV
rkubTZ+AF798JfJa/nFrnEa2pMhjiA/4qtwrvf/YVY2BGb6W5zOZyFErbQt8yJUb
JGMMKkD0dYZ7fS+og0MhVZp+8ZNkTU2WDay3HF+aTIEF52kNQKLPW6YXh/dOJA9e
dR9gVAfSc5mEtYolU4VMRlTyONFoOESyA4uROSf6MP/Hpe8acr5WVKxHRjS+Oma5
mKw5+gv9eYi4Ri2S10x/nhwkYbso6u0h/VowMceShXLoSgI4tsnO4gGXoCDFgp/r
zD+qzYetXx9sQrrW3rvboMLmxOR4KEB6CySaIkk2hpxf1p4blAnOTfaC+cjXLEgo
dZNn6R/VZlLtX4O9rWbOdF/j3KK2WeshxsVA1GOXdSzLbQX+wnOCDEz/j+ZIr69I
4flEFyRvWOq9EXMsKs4JEyfOOgDb16musi4IgAVP3g3sTmDHOaH3moE8CAKmplRf
K22cTv+lKgw6dfA1F/S8MtWJ2U9FndXPYIDqsn6RXHbZt4dZLRRemrfdtACEhz04
EAi9xLVzwhidvE2tmC66wpQIbP2vS2NpZXBMkYi2vo7HUhlG4x85dbX9lph/4sTa
OdiDV/zL9yy47Idi3GfjhyJU/alGEJsHoihZGvVYXSVLGsToy7F5lBRPvFJ8Mp21
2W0rk4surn4xtlWeKbcTRbDYgbdVnQT0Yc/Zn72HasLGfVJWO/TVQI7b7ha6objR
Uhu7Ab4pNapr9zDDS7fHWuGTzQiVy96XbSL+su9+QGky3KmbsZ/h8RBzhS/NECMk
OwcEmaMZRXhbCA1BdXaWoeK6JJ6/ZXYG9IpCQYmkTVzPhm2lalbEEF9D5VakgCVl
GKaqArXzqLgSPBDaO4N6pZYN/fahH0MQ1lq5VF8jM+V/3OFXSMqPK5fIYn1Dxk9J
O1SkZqXhIoTDrn6JQD9J2SnFN24MinTZ21PFUbUY4j4iTIGlM+9cTDq3PO77D2pe
y72Zj9JoYf/XG0TKTw7CD8R7E87babvdpjoDxLexd9L6q1ijQoS9Mcjh5kk4o0vK
hAxhwneqs2X+4ZBx3WenMu60S+Z6F2qdhcmGBbHKPHGgOpwJNjlE+Sq14I+2v0mc
a2BXluvWjPPxNJZkrhLMTmPi+STOVVUlGKC2eTV7H9rHurnCEQmrqmb7p37nontm
ORlYatnxquXg5EF3Ni8rDDaLNmrW/erkns4w7t4qUUzMUwhnhzDM36Iaqu6NPPsy
LmsIYzSPBR9jo06ywgBrM/cKPuHtROJjPtJislJLMjgdAz5nkNA4tF12wkvZ8Gs2
S1WQqAhxsRKcs/2JHUuFscAJLmdvJD2lMRPCgtcMOWOggJag8NgD9POssdvP5LuV
iL0D2EM2Wi2sRO93bH/fdX54tsrWk0316iZiMpODeykE2o334eHTxyg5kDZk93D0
0SZfRml8vVP5lJI/olaTssT1rQF48HmpJvpzmkf7/yKwWY9zpwUDjaBOVV9eCg1s
GNsfJrrWhNFdwo4NTk75yYR1p5DGo2sFEXV2p9HBvOk1z3+PQkIf8IKjGRTc7RvB
6CgN+PbOLfTf6wTZSneQNLWbZ55SxbSGYDTTgEfPgXX9cs+l/TVnjp3l0oKfMASQ
P2R/cmnZO/j7GEZdZRiVz2b2hZXm/i6bEvWaN9lISn4LGSdAP6odP72Eivgvw95s
we/7IV8rQ8tCa4Icxd+TlDDtJgk8IDGzL7NjddR+0CsLRQPyEGsUwsjUGMb2BqKx
lWD6ZG/DeRpi0PFEVKTgZpee+NCt37WmBkrxvjsux03n2TsvkU85hD2OJS2gj8JL
ffVgrnou4+qiYibzn55gYwqfTTNu8dFJhAbiOi5IMvBtH3Xewbtt4X6nrkYzNvVT
kDj5g7YvogmguwX95vKiFrKSPuDE33UCmUaXDq7n/Moi2RO6jf+vyOy+K7U88TlB
cm5FUMZZqKGfYlHYe5NukeSqsMHMg2ov7zysPr5V0iEI9cflbvJQ2MhbEvsTLIF2
sBmMPdXdYee+K0v0U8LBSo9AhyV3rTyMIJIyYgYpKp8JFlYU/z1OYJ1rrmK8BnPX
eoRPcgzJvZ4yCBycbBA2lET0Kt4VjKv150UpT6CGv/M96KLO1rcwyZb3Z+EfDVEP
bUHg3M3035o5jb4pCm0fnOMBDsU+uJo69gtahuWt/ahdpVh9CCC7CjX3ULdqrD89
IGZv7Cg5H2ErsK3xI/9tE5Zc1wfAD3bP3cuHMzMzSzr8WQjWzS7si6T1aA0Uze6H
4kpVQ63ECCyyl/TtpVJ7/nmNaGjbFfY+USyKhC56NI+erGpy6YvZzm2MMLVeop7V
8UPdNORCJ1nP7MgJZ5ZrB/xfj3R4pZHPFtBYE5en1e0wyfMb3XMzfLhzhjAunaJU
0L/IiybzLvtpvT76nN/3HbN/HVHn6w4FQZdXnLv9kF2GDVoaVJ8wBhKFh+cTvVNj
dubAENKOelWeA7IwBjR+A9BejM7imdvc8lnaode6dM6r8mffTvMFz23u/1G9m37U
YepsN2eS5zaTZRMAalKwSGSqMOk/k004jEIjsLckmVbkHQZS2cOeGftuQtZshnKR
r/9ooKSWPqG+E4ijr5lk8WLH98NHCTYwQRQ1ZdFZqiYvv8AfUeaYOEEBGZRtNQSD
sRY/IAwMXW9aPmjcfEU9aM5JIEBd8wwxY44HWou9bfJ+z5VFLg5FA6fVGwVPaJfR
ofKaOtWpNtppeb4GkvMNAPY5o9rmSiVpJMHlleTeRHd3MGKgMOCxuwZZ6z5tAklE
WxAqeenikdenBunmZNnTbzAgP4whyxwtRDfMkNfaup37SybOuCC8DZxRD4fdwlqg
PSt1J/Fj+LRMEtAbdDtryFbzLmUIaGZ9xR1h9Sim3M4ygKBVzjSDPLsga6WRJvSm
oKAslW8U3IQzrAkNRiFjmbcLov3nYjYUMbyjJCAwvYvUuMCLTtaAFiQfm8XXMsIX
ofvFYsU0R+eXdeA0yEW7jiM/5kouQKEA8da4Ga5ol1F5Aa2OMMqYdnDymQgviGgG
6elNhlcZf4/6bfKjeMhXJnHtoBzThFrYlb4YLj41hOkt8JyPE28XgMTlcgPJCCsg
culJOBTSzIxnMt2ly8uRosSJT/QRHcufIKeV1ZKgof9RRw0/A4NTwn0G/5OU2UHP
gEDO05HtqdCBO8TlCYrES7WYk9aycQYKrXzxSevt5/UhNZ422qmMPlSkZXldW9xb
LOfcOR8TQbFk8Ckg3WVZ/OMTu6wJTiZ/99V6bnvOGfJ8KhSR3Z/txRJKWgDk1G/b
tuidr1twO8P5QnhNd4whqFDFbW66Ce63Wyqs11aEozwWzDszppijYJ7yOWTn/Bzj
3Er5Lmw9cZvcy5WXFP7YWWAcCqeNWqk70EboEKW2JI5CD1HhRFu2vAtygzNML5Qw
gcCle8bRrTDD4JDgwiByO8kHTjEL2V3ePzG87pQtuuT8wT65SSCiHxoKID1u3gnu
QWGKcbOUhwmMDo/xr7GyHW81CIBZlKC4z4DPEWcEk0pUtsKTMF7Nm2BPNynah3I2
zqKBrJy9vlO9R1odi1cqI6UKkuRngVka3os3JO1WfIsd1/dgWVIiap98amhSlbpK
0fEeDEA3Mr9FEQ/V7RCNFbTwlMYw20Va8RPbmla6VcLG6woeC8j8LjASb6E9y+tf
MQtX1c1Uk90Mo3XKpPTEbw/CXw/eevu5kCWT4ezp6Bc/YCnkDeaXfov0Ff5RBfYl
4JNggLwtG77OEAefbK5XHJrYikH93UQyxYt6zsxzrbsB+Poiogs4qZP79FE/azFl
D2ugmHruQS19i0kknRoI69ZMOudrxrxfvm5w86LBNEvMSitCxiucEQRWHc3ehIQ5
06Lsh6GnlsZxOjnE5wfhjyT1lcKIyr5xO35w7WuRdH4p5eoqf32XzGrjx9HrRtv5
kW4qhsO8LbInQRvfo7MeMbJ0avA/H9KhOpT3Uh2391koWy/ee1/+vmzLZI6vubf5
5Us/mLioYLbuFab7ScJ3aRSZUsdRip54/EQtCeKS1F467D/oES3kTq7oPKWZ5zrn
SAiCGjIxYjK2/oflQXSFoVyY9IKUNvaMa5tjdxO1onnih3nUq1atuXiAU67vdKtN
iX1UWqtFLlxbcEcXOD0wXgX1GxHgyRtdXEt/9tudT++ZccA7b0IhjR7s1tT9RjVj
IqGlI49apIhs4uRK5qZMw49hFA1Ahr+9BwYuqGKRng0I2XMFaqI+hMfvm0jTwFss
TRUX7CxE4r6C6nUSuCfzVfBK0MG0w14T/oCDzCuvqG7BHnGBbm15c6/b9AWi6Kn/
iagVrG1UKx50Z2w42J+jyLS6JcNI/m1iBBIXUqb054qDI2hSIbsPb4qGZ0wnoNYs
ZARYspx5MUNSd0z1ljccxg3wNYvwzz23p8xF3iUVZKdjsNfyVXGAsXZDYpqVvvm2
w99IT9PeiGUUscVZRCMm92f+n8Cc4RrTgD+ws8W7LRlVkTvJNLeEp3FuR73AWibr
p3megfeMUsDQR/xmEfMJsO/EYjtbmVlO582ZiP0yTq4/kUjfMC1OfbQbYIwnbVDH
svug2cBQO0VlkfSInkuJ5HCUnyWZq6l6XdrR9OFoOa3UMjQHUZnV+o0SPfGQ8izH
oFxBDW4dI2qGKrHxwsms+s1mINItJAK34u/wdr9rPmmFKKSnnfa09Yz9IYU2aYHy
lJww0qTvXCXMAfmp8BnseeVjw+G7EyfefWLk5A2nJLUh0aE4sA9OmI4YWPeuMgW+
6hHyIpTCmgiqCzNW3K8991iEvxZsIbq8K2G8BpziSCpOo6QSagkCSYTpDmoWeKsI
qps7HZA9UOFEoGiYuixm5Dj1jTpa/sgC4/j1dZf47YFPq0+OMXFQXnCk7+eQgpr0
+U6OJtSAOnqqq0k1oB0I+UxFhlahxKc+L56lQPlfzZP9JUBAg5JXbICrQZHl2tSl
rvJhkr+CeSUkokyvN6hZz74VjCW71m33WKlky7eRnFkhm4qu6zqJ5qAoe51uiRxp
56c9ZS2olpywFfWXYd8ifyEC7j4EOlz+aghjs1fV9/LsYlljeybLOctPFvgElBoF
pbvSfdSk3l6DHjgsOgL3dJ7m7yc3fSP505up8ZgrmLq+3C7sm3fujt2HwXsZYueI
YWuX7Ew1w1BP3zXkmuOvQiaBsV+hz0ZejUKSqLXsRBuu+4la1fX6PcNwT1g5KFr3
s9TKx+CqxFetjwILuNNQ4fw6XN5MsibyJqjUysY6YFq2iS/rHtiuFHIGbRIQmVUd
XOnwb4H6fAi35K1TofVGT7VDlswAMnKaz2zYJi98hkKhKeLzw8vNGiknXK4eqzfM
C63vHXia7RIu7/eRSzZ/m2bJbD2/DIlCLOBxwyTsItbPHTMe2Xbk/tBp2f/Inrlw
u9XclXyi9efv/uVJMVkBWiQbSC7ZCxdmXXQ4By+Yta+Z4wTNo+An+n7dAIBNhjYl
uj2z8dVpO2EIlhBm9c1addMES+YjUPbH4xEFtH8Asc9/+vAsUihR6l+9PPPThqKw
V//FAPq+slsIjj2W9r5br6wk40e5suPBXMPgZ62U8+s7KEbPlEGY/di4Ro9Ks8I1
zQpr+g9w9oJF9kXF9iqTZvpKXJElgVHqR+J4XDEvRLShNBcCDA1+U3MgJqZRe+4B
vJ0VN07zT5hLNJyuCbZZh8Ec1BzY+BLf8AoB3RZfSluTEOTQLVQmmKOMcrMSUgcY
mk2XHvnzjYMepJnRLaViDaNBn++VXK0xsDiBfSAL4ClkZFXqBK3fKx9LnhEzyQTL
egXN6YfSB4xxu/NW5WiY5FLl7EMyPVbtv/HnVwLdcQIX55xxjZJZnWH89WoHaYsF
yoCB+3PVdujBRhBIHH65F1oLT5xpF1nlkBN0yxEWhUKu+udaOkWZohsaaDMXnvQ6
YUKNusdHTFjIjKavEABgOBvwTHAF8BeanMtMf6WbmEJydhSwbYhOCsyFJ0YPu/HD
fR61YicKBDLDGDc1Z1/oyuaBXu75eLUlTU0QafunXnt+FFoS20J8iCTIRYmX4SVP
8zX51ekVtVwQnToUm0DDzBKYYjchDXps3UEQUz0MJE/zLsZc7vrAAi5rA5p/1ukr
wgEaXvPo+1tFXG8UG7Hx9I0Vs/ZIHBwJ2BZ26NpQJ1OuKtImTUtB0vp7WQ1az5xx
+XW1GgWSxtQ6cd38QMkV/VhhB0VM0+QhEF1XKsaIGlKolfuqbgP8iGSKFYx5W29u
VGhvU6h6ml1eKEOJqBV2yAocKLYJDX+d59RtqKAOOTG0ptn9y5aej2KVbqlDsw3k
pzwfhEPWpC4feEJFG/JyjFvt0WXopuLKNOqjMjZ6E7CP7GD8WD4B8Jtwu9n+/EkG
2YEzH99Wx+B//nM//SeWlHYASNBeiiiSNQkGsLFZuEexhUQDkgg2zijKo8o8wkI/
jta23gsu9I9YoLDAa8t5jPTDU46+uwU1aDYMnn+uq9DW/mS5gunLjmnT5kBztaOQ
Co1I8FKkNhnWjh6+HyvmKOAojS4gPmnsRkTTMfm9VgvCnlYfl3RF9BvTkETkD36w
mIbmmD79kfVzOV37zxDejRZR9NTP3rjbRPvRhRqIU4jJ88LBB5zHA3JRoUCwQd3s
x86J7Pi6woAPmlysYaG+4uEPH3yuOaXv0HoiS2BUgzBXUAqav2aeJHxJTJo3z5yP
2GDqCvv+GxnSzNu5p0EzqKemDW9X0N3VN+zEJfhbZZeRhIiSwLtNC5+H7+NZUCWV
rXtpzQcD22p3W+wagUVpWU51zsw6ODyl6hs1s4KE3bsL3g36C6M5uNIFXUwZrls0
iaX8m/pVuYOzuS6rMjOY7EQrDSJ0kSQuuFwaYjEhAgJovGRNXuU63K3hlhAtlPb8
M9pzgSnoViUpxPS+SHxfLVIbQinf0MtvTo51XRFq7QW280WoGWGCYapQUTaz8TDL
mFqezYzAYX3FQD28DrK+nVQ6Hde4tg5rD5z9KS4TW2s37X8Ez3J8QCZnhAZaT7i2
vt7kDFoZbCYy//igFjImhYv4HpWqojl4O9iHm0ntYgDIf3+rMTxcOlHnWVQ/0WyU
yhJicPXgLFVy4x9pm0BEh005v0Wt2JPYFKi/2fkiFVvXU2MDkZc1JUp8XErxvptn
dKBBTi/tDznZ2FPfBUUaAHolNCt4ZOW3bz3P8a4uZ23vw4S3CipJVYo2bVnuiZ2x
WUhnIYLl9+dvYvxl6295h0Gao1gBpu2SM0KL6kPstjVhQtq7e0ixevPfvrPIFjTY
z1tYj4mYDOwL50N4ybbZwvMTiAHLLH2A1xmUSQcS4UTjtn7I8IP8WOY+OS+I+6i7
aztmOL9lxTuANpttWKEu+hNACV8AJie8RpWb8lGL4MfVEe023xyZaXdrgrEH7/Lf
9YNKCreWZkT2nKTZ3ViZUXJZD9A5YhyyULSJYi0Nls/NOlH7btiEQxTestPp97TE
yp5EPtxCpSZPt0GWvtC68pcCZKzL3yrHVZDUGCuUzFmejKssb/osNTd8Ql9BC+d/
k8OseVcJQ3k+he/3Pnt5hSmLmWdxFjOpMiys7h0enq3naD5cskrU1EDPUzEoIsy2
pV2COqZWvHuv4NFUv4R5dPCJHRfwdOpTODxU8eWrKKx9MftEoQR1LM7Ph/5ngZ7e
GoQJFXLwvdJ3VFdbaEs/gv3YZc3DdxWiqzOtNI5pzMttAwBuVVbqz9wfaHpD7VGj
UWaOOy5H+SFFID7KjqoPS1gJNt+5pvByuPreDnZ07xKK5L6IWhI9y663A/0mRUSr
ytEG83SaP+L+qmg3icmKjgbm9ZRwQVTyfpUKL5xipag9yXhdwQx7d3DCxm+VBUvv
jUOFosdQEg//3Doz3KYvwB4pvJlNeyYyj5P4kZwVmtp7MdZhcMva9ZCrZv7LTiq0
BylU5cnEBbUydPxWmD7kJswYkh23GmWEFb9CXpCYbBorS+bLFJCbj7B7JTD7Pu6R
XvrfQUdi7VLovx5pHaAkcqiqp28pRgFGlPHi7rzStAH19wL8VIt44tphBR+4oqyK
ezCKijGESGNrVhApDPRsNSkvA3lqe/0w0Y28eknlcujmvUlw7e/6MfksxVwuKBxy
dTMzNJAYQZuVL0qi+3L4VIsfjjvXOeDZrTE2DBdunkX319n84xHII7EKQxOA8Wtn
BDrQgHS3q9fXDrqiUN+o2WbZMVey7z03HHT9k3qtajEbGol1TtFQdfMnnBDP7OBd
I5VX0vL/CtNNbHD+GfIyEKCPFUtdN7Wlxb7HVH6lENcj9E7KBj/XrAXTjd2iOB4m
uIQ77nDQLbZWUaKkX/vM3nv7QLtSfELLZqzk3156VfwfAVt5sXRtJTM0oCQECsuX
uZvwX9SJI2vsLeie4009PF4gDm802GEUvWDEAi969Pyw0PAbW77n9IwfxSbrHwDA
6MPBfUP6XO/hjfZwxOHku26MPvMAnQKIE0c2Obrx0xz00j/MH8IlHvYp78h1ldMP
wYyE4Jc/04qfPMR/2UspEDND6GrfD+wfa2omFtvOOlX0vXnDtE5kQBMXodHLsBOI
1clXP8oyOkMgxk4hYuqD0LHsxHLP/I/R4xHpUqvCExtP8cxqjPYeUCcUt0H7yrje
Uwelt7nxgabUCucRIFCP/EnnsxxtsevoGUJdVpsY5HVaX7Ei0Hy+HMbElY2ZlMBy
XCgYy1Tnnl8eeZ9HlGIAIAyVeWB9aLQQIF0OCRI0/XYdu6TvRuYH7FCkgMkvY3Oz
T1v+Cp1oglPbm+6GLw5GBlbJZzPnSzRVdOa6LOEHec7aT30FPVIFbW5SnaxYrK9N
v35D7DZsZJXQHVhQcv/9BoRjoYv5DtZ1/majpwH8jLIl6W7c589Zg1kEpwMRaF44
sZbqGkQ9Aeuak3qHUsH9KwaxEXtuFg1tYxWSuiMAVjjVHtdtCrmPNdkdZYesKaEe
F3UNcGfRmapef2KrSmdkQfOHOEZ3m/LdE6eCqU4GQWvE5GMFb17WNblmML709x4c
7mycOOOMWR0EkOyj8Rym99FIdB4QKYuEsk2Gied6hVGvSkC7W4bV6/J6ks+ZmHvb
1+QheAvyhPmIrKDOc/REgaCNTaVMll8JrIS2T9pk3FkAK8hSds7q9oYb7wBbOb6e
APC6sa9cXzSt5+2OC4NNktJm6YRNaxCW1DQvb+YABH2XBkymA6kPtpr5gIOCjcV1
dHh8KK72CFufGupyIotD79GueCEO//MN+9qCgvzL6+RFT7KdFl7N25hE0M6eK86v
Mz25xeIHc2gpM9DH0HSeSIDErppewfGZjaKouPxzjTabCT2jusGa7YrBsNIxs1Ny
TALrpRJ4x6mcoVyy0CtWK9Jcdadthrmq+W9L3TOFsy54fuUme+LPgteHzKJSGY5X
IDMf7wH942fv9E48rN4r5vv1zyyFSzpiygfempdPBxLVTT2xyyGa0y5pkfasxf6Y
pThrg9a1Xps5lvi5Ff1+/WPpp8XXMsVYLkbOjWhP7jzIPYiM0yhPPqKjIqgWsKYz
8WYlw/WoWDhawqaakUdPJcUjxhYVoyy4EyvVhhx5eBaahs1B1rIK26ZFoXTSTJNC
/9Ktj7MfzP+8tGq5xL4qELHs45fmSqJSyqcNRWGS4+szipTAMW6HD7J2fUE2MJCQ
o3vwMfbRcGJjDysROPUGkXF6VTHiBz7ZNtfpK45rlei3hGsprIEPJP5opQZU37OY
Xjg92YQWf95qn7D1Xooi+gW5OPuKknSpwRIEQIpxsLrW5gNMuNYpJqsrdNdb+iB7
Z2knKP6Uu1AulGRqDTlLCXHazd1MSuhDmT9ejgWP56Vjg0cS7fkB3qez7GBOynWZ
GsmRYXLbcN5QS0OlFwWXjbKx3f7MDfVC485w5KkxbXq7qoWyWDjgYA3oGxsNmooP
q4A2EvKicHjaEvaOCgirS7BcBW9fZFFNNzCfet1DIbtOc2+esfsRpRepLUYgswN5
72iyAcXVHFnsqCzF5jUF01oOUARH5HY+DlsxhfZ+Nvbz6R1zTGCVUoPoC6EuLyT7
AuJUuk3C2PqKxnGkuBEHVJ6tKGW+HcISRRcq4alJVuhOh1tDOE0LovefndE6o+49
hxU4zs3VS4AAVj7VooucZ2GE43nukjX6+XIGcu/T7wKG1QmWl6Vqwp5RnA3dbrcI
VyAGcEmwJBhqm+ueEqKHcqKAV3nMwK2b+sHq9TX1mC/XibsZnM6o/Rbth4ND8oY0
Hw43beOnExoiiajHfOhhff+Xtn5ixWthx/WFYAYcgHFlDcI63RbLk8eNLyZ/BRZy
JMWa/hamWuljTP/LXTppy66IBaSrSw2NEdndWOE85FKYOkK3PfTyQbczT081DALE
K1RDt9GlKCMbtdWZ0p9vhrhRXiiXXamjqYuGpJ4DMbR1oFFLIJiFK465gXqv8D1Q
1fgYkm+bJkZZCQeOtmq7LSZfBSAhbX1ABS9+79gq2zO4wPu0FJPcvQw92Wj8Vdih
PrT0GsRZ+e2/gMcJGu6Rdp1ATvP3Eb6oyoYwGTe8C7lgeRnv50H6P+9fs/iCCQxo
pAWB/JksgJqTHV5EJUfZyvgjPNY5M58rlo3vfV3J5fATa9Rqybe62OGz2hI5VjzH
Y+Lkl0/xk+nk/sVNoc9ds+CgtkJ2Wm3xHs/dmR0K3IWjhaNt90ZLVNekGzA5MaLz
SsVLjmdxh7PgF/xfdD7PFK2AQAhIHQTAkXivLFPdfaLuw/y7WjPvQ3zWWC+upEbn
iFiHhP5iWalQgOUcSKc5ZgRNXkzZ41bqYArErW54KYKu7wgjJVvAWTAVvthwq2g3
qscc1wa/B22Y3bQwpbvhR+6MkxFqatm2PX9UqDEPRSAaJrkCR5uXVXhEDIjpxsGj
fdUnrrwi4YvtTlOzyJXileGIPO6Wm7gc0xzj0K5sIZb99/qj8uhu1gCHWeE8z+6y
RX4KUU1ZKQqch083QMRqCUOfWZE92wbYEF0s/VuSTAc4GtQZXCrPZeYpjHiCpMEr
DrofwTsZ1rM1Nn5YLj56mTDepjgFJ1ld76bTLbZLquZSJSxeC39xEvaDpkPeUIbn
Ah80H0/FArSkAExXtPQbJ3DaHjWglumC/b6L6mHXRn+k8sK+rH02a80TizdFYhNn
LPKkZPRuefuyTjISklogjxoFzFhJANzR9AgCHJDiqHQfJR9giKSC/e1uUXsKt8kL
4/xBnteCT/2ysWOy+pjmN/F/yNScIt+k6+zSYuTF2SyZtxxSRa2fq4u1eI+ssBR4
VgZ/bI36DqxjUvK6SCmZII1TZomCmOGC0wxpeBhDq30qfNKYlIlXdg3Hj+S80/j1
uXDicmsg4UBWdbs+Imdz7Dwe0LdRxz+0jHgiYcBwcelcGlfdTNgsThCrMDrZ88ed
juPFuovf57l+IwkiFJEWdHkfzJq2H+c4/a+fFPJvLlrMeTYwJ5W6C37MAMNnrUbY
5IO6lmpACiMyLcvDP1A1RF5vgOHDja0jE/DUD4xx4tN1HE1BtDZQtXFocFGrCl1W
wOOdwlhQOCyxI6uucjDb0ZL7U8u9V/+HIbn9eFHXzQTQsgSa5G22O21lC5wOfDmv
pkP44u5HGduGNk2UI+pqE7p74rHHPr4xC9QLbAauBS9yCWpS/ty/bJSf9plQKlLu
woWBShPUEbnFX9uaCsRBA06xXtdSEJu+RFB6R2iLgLUVkvg06qxvMAsiSx7ZQoOk
wOWyFWtH5YNgAf/D/Jf0vI8QEvtEOaEmr6dq7SR/XyGgdfGAAYIDnbPlPN0d2QEn
izBPt41s9x4y4ImGAXBNSQqG+rgPm67gddUeMYxSm0/ttvZ325GMn9JrxA12Kvvx
iXeSHYTg7b2tmKVVBvInwoIgg0qnNzgLChTspSwuibKAguXLq5k8aZ84HXqtkb7p
HOn6EUmq5AxKEFrLtPPKlBP2/7+hY6by1o8iqFW1Y0XYHWUnEz0cKE5T2CUW8kUe
+FqdwSELX5EV/bF2woY7qxfqH2bngynoq/xhlsvn7a8ZCbDHt8XYWuJ51cfI3ZYq
0haBldNpQx9weMBL/el5kxUglmwTLNxUVyuLpscM/tjGuuPHW+/EZ+ghfb1N4CCI
yE+4TF7142PM4k/Gq5cpKLW4UHhreeHiUNkwbMQR/QX9BuqDP4AKarmST4pkIBLB
t6sIwgWQVfGsp7X30c9aKBwCMeOtCfwgBN952jAKFik0RI7aWjxcPYRS0GFLAD8T
24VOXwl4MfdzPdCxKk3H+dj16m919aAP42ik7qBS6Kg1N6bx2jcMF3QJT2BVrI1t
HniZX6SFELTJkApOrvCmCc52UXmpXSAyyEVUu69VSiMvZRUuyq+7cKOA7mHwrtqT
cP9x777iOnNQMDow12OKQEHrjUFd8gAwr3puUxHVJFSeqgz6pVOp3AyjYGj8nPK8
hHIvyqzdlCUr8hnCs/BOFLx/jRrqlJdpNbY8NAGeO3d7/L12XnSVh6H8JjTnyeZL
p2Q2L+TJY4yvdeKaLGzPOVqOyI4XW+d25pqqBZEadObW30ttoldRPBC8pG51AgCc
8wNBWri0hU9VmTPfzU/O9lZhiiX8drSwcEbjuu5kyuVsp35WADfvfLTLvqR+a2fH
kzIqWBtwGISSIpkTmGoTsE0vFdOYYAciob5Wcne/DTG1EAsUqE5AgJvcquh1b+jO
MjaKN9eCgR3HGk5XDbVtPGrpv5qWkFOU1KXMObkbfmMEiYW+1/Da4yGJtp42cB1j
5WiLr12puTts7GZ5w4cfphTp7+2kK1GuuzX3WfEu9q5vCE4ocIXjXjM/KyPgFyhw
4fDm0bxxdewrVhAEs+MHtFi/6bl7/CV/JGfK2aefpCSg8LWmCh4NgFNCB5QKjj2H
7FjFgPAyl3aXRDbuLIxUDFuddTAhgfmO/nKfxScN5zGuA8jMeWLPkVbk60Pcenmi
v+atiIvDptuDD+QakmpulJ7rdKWMZME2YwlPzBj2Q24upa7lxuAJUMi9ImdEiz3O
CVlRgP9JqVkCyVQqQJCGJEI6h6HNNk/KxnK8IJ6pdGIbTV6xKhwlt0JZi+ayAfmV
BVCyWlGi5RmFaraprbf3jcoIUJ+KaEOTKgOD2PVsMn6Xr0+RAGqNR+UmZpcdYLA3
FuIGLv+Y5vPisOObOkCNHMM2+u/Ho/FcTj/rzAfQkXWQSQpPGP7TCKt+FeVZUyWz
8x2LmSUnUPYl5NWkZyNBLrp/1qc/dZO0njcZ5dyCgRNWETJ4GMCAGLuXYNEXfnp5
pnFR200M+pkh7IhoohLMr6BWzikN7OF49NCu2hXqAszWpf8qMY1CQULrdacnCcrd
srkerLqc6MJCnzWFdEJY51iq/iV5WVgSsWtiHORQIxElHfnmo39ejIlLmb7CKCsJ
zNsXJcUwTzKXRrQXIhuwF7YOpENOJemDMGwhoHeAb18Yhg/qG/C4jO4eyP7eticL
q0b/6oZoqluwTyFhemBNItKXLR2dWexsUvVQFQI76tjOM9gQEsZjAw/4/oLl9ywC
vZqfzRgP3huKoJeB4xMHAsPY/3tyvWjigd+waBjFgzBbE0MhCWEHlVc2LuZ+UAyn
zKKyI3+tg/nOPodYlZ3iH5YddM6MJcAVR65thgj58f/Pzru8JdFVRqEXpj34Hlg1
NZaxHqB1DY+FwrBPZzUDuaI3s1W4VVSUtFAyXzkpiN5MFhDF4mOUYSOuXIjGRuYw
UUVnVJ+zhvIjLflljVDd7pt+gXUiOVvyWqSot3jfuo8frgjoHR6vF1I81XRvaNR/
JwjOS0aBz1FxKO8AZg/l2VV8wOn26ahkV+mhW4skJNzytcuLLQuYdFfKHUVJ+Boy
aYnWLuJLPKhRTyO6dPFVoHtTZ5eDKsemZMD0rcjmHtMDItoBiu45jhlncWNHyLEO
1sjoNLZWExatzw1KXojBEZznrpmD/S9hZ65MfvCW2DILu5a5DyfKWp6aVuqERDBA
zYGYwfwgc39nvJLTyCODd/a5z4B8G7PLqhyRCJqDWGNYr41goFDj6zBMof1sekE6
0eScmz5xTtkPkOjPWZRtGGbyeCNQmpYi51MkxhURSo+bueQMGIxCl92qr1nL+HTn
tJcVOD6eRMD8N2rsCf8g0yCdEdsW3UXviAFC10I8WBv+J9bs7WozCJ598qlBnfgS
K6C3U4m+Ut8WUh+GeNoEbXEjeWv82fZ8GMQC8cWVzEQZ4kC8mcUIi7TLTngaSPMo
XaKkbKIOjMgA+YfhKyS1NMFD5u9hhdUAtQfhVAPZCiKW0bLFT0u/LXdtVxAnRabV
2aveQMjjAQTHuLwdcXyPRsYxfBsRF7Lv3hvDq+HH5epBqHa4CvsiPVW6NmhI2ncp
mKDTPmQXlup+KyqUc/jp6RCHqGAHs3HIe+JEbwRpiZZs1caaC8TBD9iQcir2SZHr
6ElHGvUVrhfuXPfSs3c1z+FbkOOojRprh+t9Uh1CdN+steY/6Davnp6njdd4zHGr
E5N5ExwDwTpi++Z3dSfMSLjAkDtw4hp87NED5XJNy3wCPjcHOEs9Q0XiEaK9Di0t
nhxnUv8aY7rUMeCdS7L/kaStcfvjdHUg3O6nWvakEexp4ulJniTcsrDJrpdNfenI
escMhZkvgmJCkCbzlBmJclIUNcmFAxcpQ+WjZNbyst+kQB/7fUHS/7CrKPuOtT5n
2KnGDYI0YrSbEN9L1fehuh4ux3UUdeU7nLRm/x7XUnZRbKtktgGVSUD1/0A1rS6A
eGAKedM7ky54f1whBR+q54pcWcoI1Y3lsSbULo57uw4fYbHz47vZm8sCntZU3BHK
MIB+/PTjiUL94693pZfDAixugZaTWf6WMwI7dtlZ65pG+wROBpNEutZLMsETrnr9
Mp77xgmTxvRrgVXxx1HVJ7FZvxA8LC7VMN8gL55hMEXPQo8QKUAsh22L+2ZfdMRz
zIwuZxTYX9vtdeHNRBvWeuq3fDdO3cTYBszB6HKVClitPtg0Dd/lANENu8OziqOV
Ri2+WMomfOeG9fR91wdf9Sozw/5HwUycUbH0TiWi4+AGYIIOQ9SgXbrCeSvZEcm0
UGSk7utpyGOzldak2gcf6nRhywn7zta1mb4MzBZch1Vs/t56gsCNxHcf81ZVv7hO
WnnJGe31kwgnEYjK/aI99dxAwUDph8pMO5RrdibSUQ8A2aJi7o9fN1oEw41fpBkx
wAlXCl5vXNhZOHqgn+TJujvOi8CKDzyWtXPbqZ/nE6HKagd3GNUZd0DiXnvo+F8p
kRSiZpYK7SjdqSCZSIiHs0baX56ufXMR9EXKWYydi1nT/irNQ+Uyi11X+YMDBcvz
458IL08mX/NaUsekpqq9a1vfLJjngCxt9sFJu1wI2lJYkqK830+57nUmL7BcMf/9
Pv48HZi5AaPQI79NPZmkp/JQrUbnYDpqmHG5LUZrLdjDlJtDMcl4D2svZNCdUxMw
AyROynxX0FMe5kAtpvMejExtazEf0EpWDVfrH8W9T+x4MIyb/IhSo0l0H1AW/X5S
1yu2Gyp9WZHjFayKBAsaQPvtREhFPMCz3XtcEmPamcb4g5ByaShddT8P8u5CNs+5
pcdDFag9wujwfE1ohkOJRW7lk0pCcwJoJfNQVUPWFKE9vReBqjlI8M8LhfNTukE2
PwyNLDOA/nfWm9qaIO26gA2sgLmh2DI+zcMVOTjHWm++Fduce4UapCNGk9Gsrltj
YdC+Iil5peC/ipqyLxMiwx7/FznGQvtR7BRZ0RpJ5FLTqxVmSL0eBJTqScw742v4
Mu36hMhHEfICS9MNyDsw97Ck4StaW/Kro9rTIbGbasozUW3YCJTal3AlyQnpz1HH
ZS/2CwN/D6hBi072Rz/PucZnJPyVAuxYuDLWr+VNmnoWEyoVRhTMkRVeZVa7pe2E
dRRU6CufRz42a5h9OH0sB/SM3m1BNQiyK2cYb7+AGxQVbk8Vgu7cVQNHCQLKIyrj
Tw6n1Ahih7HbcIOwdF0gY6/5n3NANlDOFMUxXAxPDvEvdBmpcbV2z8WQs07dRlRf
soCyaSXrsr/0to9+kwvzNbr2Rp4tO1RlWhllVq/Y/rtunTqLgjGrJzHFSAbMz882
u1tisBlSyyYlxz9EFPBMKI2dLEWdvq4//UB+V6VnRjVu0rNE18YqA1F0ra/VllIr
r7ueCviyCcktGsvNgTVN8i7a/wGS1i1r0646of0iSreHK5BBevxS0XqgkZArkuSt
7nAbzV409W32wU51mRs+S8RLp/2rS8lbftqWecMK4ouDzb4dZO7quBBmsglirNxA
LE1bq9Zd9cgt2naoE/HrvMfqeQSzF0ViwPcLgJjxHq52i0B0cQcOV5IYBXMROELy
dbpmCao323zG626gYuQJfYgtj5bo4GsF2p1z0F6XZqZzNg8CLgFVhwyMvoo46ToB
R03cUDheO2R4CGrG5/JObVx28x9F/7dw5xLBn4EH2wZkLtqJakoHvoJ1cxLE883e
gk8Ux5w7ltAYrXoq1z9fB5ONHbVra1n+6UG7BpCAbJPKzbDvv8YXgTbwEke+HJJO
75TjmGd/uQBIycbjprbDoGnrFnBetuVtx1iNCOhR9XRlG72RrGUbN7X1othBeLIy
CsGEz8ePrY8rcDXOz5je2wVBYR1yDPDQp7AaeJwDQqGa0u/v+Dji/r28GenVpCmp
9oYmB/lfbiM9PyQTxtXUDqvlFwjoRmnl1zh9W5W6mr4nNueeloxYdBzYePU33cvU
khQryLLNEKnYlhqX5YRK+y0//unjOx6FBfy3QJgU2q+42xRgTd9Fh6gABgCMjT48
+W0PclzOsjUg9N/DEv0bpNU4v3VDXdODXkbKfqG5OxylsXmGlCwbV0MQM0qGHMPJ
11h2ZJSuQ71RaKuQtonSGWV2OifCWRHwhPf1g+FltWdEF8PrwY0uRAjCgls6qpzp
xWsjb2Pqe/SE3Y2q5iUIQ1/fhgYXs4MTgodBSLAGmoJ1C8IOdkFWJG650/xPG0U6
bBINkmLMe19YzIs+ZSa9yI3GYL0EI11DeJHmm0grgRwT5Kt3VqmjttMw7e7hAbF/
MzNuL7PG6Fr54r1xtPFHCX68Oh4SnQjB1zyV9Tuu0vg3gUzCxHnBBpDO+IxJYJyC
qOR7WYEmEowChVnP1aLhz4UMYn2EojhvF18gSKFzVKRUwTcunDp7udesFFVQybri
k8nTg6nj7MjywkC7v85k0MqMUAx8aD7O8vibGR5lGa128YkWRfwsxEhhgrRU5B9X
AMfm+ut2zsGx7rt4JlsZR5xNJeV7p/RJ/AfCZ9Be2r3X+9nC3+0jq6RCz7Qhyec+
yb/9huQi2ljUK9GrvcwU1c0AwkPeoAmJl2IDkHP+Acrcm26OXrDj0Y6VynjQLRUZ
9EE4d28XOGES7oXTXaHjFC6cWQNEewclxHt/CQNir5UXTcnQJYvYmtsfV7tp+WFm
OeBSvPZNQbEoUXdiMt7HFA9BCypAZ8CtNW/HHXOEDd8Jasvb1TxhZvvFuvOvyoMZ
Bh//MU0H/OaCeHvpPVNXk0mJdhjBD+0dgv5OTlTQSlWGuDYon7Gz0pPAjzXIDOe0
/1Ol0AScKx/xO7pnBZO/HP+ImTjH8s2GNkXZuknmlsBa3L36GLiiI39qX4P9bcvp
jSumXLw5j/AfogcQn55l9gWqV5/axgOPkxlMYlHxlKXbzG9HRDE7HZCoYEy1ggFH
LmSJx8CSy0+FhXx+qq6/I5rQkMNtwaSCJl3fR2USYx1vsKlEALjzZfdAREG80hwY
AK0kz+iJYD5PGZKBgp5ySQ5ZNZXIqE1bbdlmzdODl+hjAZIScTIVxMwp+avT26l1
u7hOjPrIYMj1LqZVUHy4tlathFMZSBHOLhYoFOyO25+DRC/WOrUBLQbkJMKbOldj
gEpnvzF9TvwlrgpsMMt5lsNjhmsaldAgQLH3UsQL81g9Apv/h2B7+usUMg8hDxbW
Xe2jmEOkNTNh+oLyxh/O69ujPEK0dbIqcZFGCMV4eEgnsexL/pz9faL7hPx0bkpM
mrqvFuwR+CQjyGQaP1NldO9Nh1o69XupLEiOfu/ZHIFHVITAis5xnMygPhyQU0z7
5VwD+SXDcC1U1hXQBlAXbT44hTWyqpcIeLw92EAuKaO9NnCdMCPa1z5UHManGKc1
o2+Ayq5ZvxHGUdKOkximCa7k97c0HKrB8ZmVcZWBhxTtg7zJ2hU4mqfrR8j/xblb
m+/lDe5Vgb70Sp9yjt8IB1D02TVfAft3SQKfLxD8uc6r5QPn6tCSEfJNLQsNPpF6
MzeAex4qJBwKI3eiGw+bIP4QiLsTTmA/DaK6FPzWIDwxPPgwiVvdb4QQMwbqbGfP
n4e26Z/Y5sl+bt0GEDE9XKY13wak0Ds7M3WitMBU72EWb2x2awJ40RZayjJpS+aA
GcLX6Jw8CVdyCBDYEfbgJpiZ2BIPDGM7cUo5KaDRBz+ACGpA9a7yuORSLoeSc7p0
Zxbog6xE/OXCa5NmUUOrtSzMG35J9CK45HLM+c7K4O9DTal2TEU30H1P6G2E9kQj
1rW9EOfRFlsC4wMvd+cFOyfmvLucNMoteVUwGynQG7D559jHS+a92g4/NHdUVhpv
AdOAR/ojwgjqg52R/LRS4X4HctJnmB/C4tZAXBYC+1boKve+yC0JohvaouLPB0So
RaT3HqFcmgO5DAihX61isohCCTMYY8nL4W5udabfCSt6C08Y+xWl48bxDhYuAqU4
HH5sVLeBpzm936vS1IaKcWPbi6tWHM4Sb5+7NOqIVz/6PWm9SlWkuXRfulRGysAV
odEyfCjb9De9Uwej02TdPDTqmLQsR23hme+GnHTxj0tF0wbDTIid5cZJPoC8UrIq
TtQdTKYCnu8cLPlrkyGLpY9ZHFwnZBlRTakJI6mMFthgXtoIEICh4x4LaTXs9seI
VhyYK6v6hXs6uLBPBJw7cOGqmrLTVj9EFJQmmsDMHI3ijXmlE9XolRQ0/hEFEF3/
sBUtdzEQoWetmGpBX2Juwui3z0RJF3pGq8EdX/KPCeS4H5VBGt0MDoEegs8GawTi
aakvveDrI8D9ZOKaL9YiMMl9wt+EWYkVy9w0Odmq2zyFGPtyyKm1OvYRXtMHFrnG
nXXbWN5YaGUz0HhdiodkmDmSpwWbfXO1sgOhAI+Y9AqzF15xIxw4fwoXpCtC2ED6
YAKS2VLBxBF7DeSxZQ8N1/xXmNWXcyshFKeyIhhT8Zcz8yx0OHA0WYLKHotv1yHO
AGRcXz2YdkOxELhFaLLJFpsZasnghqVbYogxh7auKGGShhuNdkoaf1LJTBHdG7EX
gRPeypbLC6E315X446Jkne6Ja0+y3gqKOuc205pulOQEjuCYQ0AWSMI7m/hAlyUc
FNcOAMPJLYf9SmyvbHzoM11RkFvpwNRe+jrWLhuTfKkuaVpRMB/YuheB45zx54Pq
T6SaDRbGBTVdfRrmvTx12UCn5L+5DONUe5XT/uTMLLTFLa7UzJhLC9k1Pm0RhQll
Zw83UqmaogBk/Hiz8Js8GGKHn4e+7bionn1k0ma+noZIC0l1N6KRZxp1+rMxhw+f
voJm/JYJNTJPcg57MM8n332/QRaqlTJe7HeR2Y07qVRbFHhA2sIid3XAdHcjyOWQ
EPKduEjGLeJVYoCM0SN4s1w7J87MZoQhHoMGqvGPy82fMjSspcNTMNmRALsVTcpi
LHVkNgBsqOGHLL/Cz3TqAFdrEI9kuvnWGPwnT8k7zCBmss3AL/YW2/+LiDs59RXq
yHzQ8psJiypHMez/AFViom64fuVRt+sz6U3gV9DFSjWsF0KPXgpwVRFYEzr0fSpv
6TtDSW24zvTYY+FRNXOnJKggSKCQN8oIIeP7Ty9C8N8Y2S06p049bK3CKy7/PVLK
0vvlhbtXDh3jixgXCUJFfNjROfEHDm8hNt+zyTZ7PDzM9ya2/kxOlHLg1N+zXBs1
jiB3rklAgmGr5acyJeGjpBmHgZE70kausWdU6QcaOfveuH9ikk3nJv0WDjGjYVGw
ic2JdLvi9lxYFA5kXxZrFENp7iYWabp8A5muriiubpx4Onp0vaMHsBVhHGa7Vn0J
8s+s4Ve9l2c8tc2ZXKeR1nM5b5vTWQOCaoLutyBdUC9AdnoTzd9zwU6Hvh0e9QFU
4Jqt4jZZhSyBePHbN7RlXG4W1ZULXGKG18qEQtCEPDvSrnXC9DQ2Er10+zGkyRHi
LYRQOELhmQP1CBhy85BKQWxjAP+ysM2vT2R4gA7jJeBM9a0RH0ODUZFv0mIbynQp
dBqluj2oNlcO3Pza0pP4QP57Ubjg+Cl2xszSMxrv3nlEiS68Ysp08mP6xfYy+apk
hrBens7/ITAgVL43ocoGMpTsUkKVukzVU3IEf5PQUcScsdWKJh+Jur92dyV8uAND
SdNe8rfVmBfmMgIJIyItntokEqEegHx2zaQ1+X322pA1y9oP9xPn1gsp70+CdohB
EFqMRTZmk33adgIMXjF5agAUEM8floFfWC6wFK2cWV6qmoR6PY8asgaMJ5tjHhd6
8pGV9IC+HEWZa4tTwjlVul1AYQBQ/0CxwJaUe98aZahM0os4YlNfvQYZqaALcqJP
nGhd2dVGgCkpvjcurHCo2wQvzhW4zW5Sz8GVsxbJZw5z3Es6Ns/Dj4iShd03jNur
PaukX4GGXLD/S81K7q/Ei9ZSwVWruENdUUNyridt5iwIAYQibYNLxehBz6ros+Gv
bHtriyyPSwVFUH3wmKmzvvZ7rcYHSOs5ToCFd/x4kKr6g4BsfHt1oCjKAe8qFt7s
AtKSzNtoPvcmQ1bjAZFjIZraSDc/O0H6ygfm1eqo1WRYOzLg1iiPcqS9ValZ5QoM
stcMhVIWS8wD9RnBEk1zWsvZJcVlpd+3y0GMx8F4E0OUkoXnAoGP47kSToCqEoC3
iz+4YYMyoW17ySY2PrYxW6FJ/LmBxwCmkhgmjh1Ec+cdQMawaCARQZfIt6Z1slxy
wVIbi5R27xUlKe5Tnx/xwbZwj+Hbodw5qSt8t7hEwvuvJh08DZ4N6HkPrHrWberc
zDSFxonty7NmyaZ+Na/V5uc+DTh8dC4roJbWY0MMmuzMjUEjcZ836iTYeEr28//9
9a9Xl0eKmCpSExqpRyPfuoQmEoV1uyKOu7zv/2G3tm0PZI/l4Bi2ZFu6DAL26ank
5Zzcq4EpSXicLrJU87vZ5lvdVh0Aqd+IKbbKTN1GC8cqf6OGadHubCvg4h0Y7r+z
5Gxz9xTBaOMjMRlW7bf8VLPePmiGvBIE7igyni44Urg74SXU5iHiCrgD1OBxXNhf
6tyoKl3288FAV/5VHHHWWmFmlofFnc90RgsLCnkCoqchNrCGSxLnLrUhyZricobC
Yn6nt8s1qzfBlsP2sq8lDPyR3LVc5Avzu/TB4TwL2OA2kZChLFc0zFtOeZj8JOcg
i3j+/libsx7dcCYUICKjRfjh5uGFnEcB644/QsNyF3tR2xvo/TG6s1CoqtpmkYju
QCAJsO13VOvQOcO7GGyEFX7IAIEbhTPEInehF0r5QJ+hrxBcGiako3FJKreuX00Y
TDh+ATgl1NDkCKtTni4dLwkBJK6bYK56/6nzg7D2XWjfzXC3Nj9fkSA0LUbP4Unw
fVZAZMlFPewQF2Rmh7ge2sfI/t5Ma+h5pfrg+tfXjqdEh4G9fq7HSP3mi6aGeGV4
HSMR6agsHEeKMLwovaBfuhJB+d3YIqERI0fTeED4fkBC/LKd3rAsO8q/AiCwC1nt
iyadDG+UNyTgUg2KxVbfWJAcoiTCfSGJD24vHvlfZGdaAkTu8Q0whxzWVCoAhIYi
eAvWhw8unECJLTkO1+utgQBhqQx3euucqFg6me5eVwPZ1Q1wl1QHRW1JNycWqdkt
oAbldI5BeThEhcP/d2UZ5sNfl1DNRDUhKput7I8n+AdJMfiyg7nHDvAV08BwXjzg
/T0K1foYhay1/cjmJpjazLMf+3c87NVCiU5cwUHJOO8BOGwU/2ZqqajiRT0aA3iB
eKhhTc6KGe9gfIo2JDEEYC4SIVykTUeRs55QcqPdU2ELR3A5yR0vlPGOmu9xJwoV
l6/RgJtfTSP3Z2m1ZL3mFaBr/PSZBrjMNvpEEungM1Ty/lX2JSMb3j8SbBapVY8e
mMFb4t1Hm12Ie8fWe/3UsUUYhwodKp7/HTriJtFgqn2XWxCQDUNNq+ptyV5NWUB8
OVNfL7ulNt6EJ6sBTXfGkdRWWDEG/AI/AU5SwMWEj9IH4A3X7+9YIm3nGEjUc8XN
dGAhHT+S1BYX5GeZIrn1dDr7I58BcFk0Za2NRrW0U2caxWZw2MirX0O/ymO4+YA7
f6x4O54gnbbEBvBhLiHSaFtYmRZ1bT7JXuLv6qKQXCC5fXh4C2uLci1l4m2xGsmS
W0QwzS+FZh9exwTUze62j7t9i4MsogzQw9cdde3dy+TA5NQTi0c+/1NRnOyBTeDk
ca8w3atSGPsAr5w7UYMKcplqKfTQQtEk1LtZv4LmvotgD4IDcPoNZaPPCEkn471y
1bwDsf3OdLYVqAdiJN8a2WA6/sbD7YKNa+Y4Ebrm7DwRWWR/jUAbk7Fpe+8LpF+c
Qkr9m84/xUmFem9Uzt7raFQJqbXP35CLANeZGrfH6XcLwqwAMsLH7cGD8/XnIXPf
74htj+9T/XLYLoJ3ObwXyQ8GMvsAGNK/t8s7q+Hdt6O5TENrvgQVfTBbgZUmWqzK
RC8a5yZ2Vzt5cUDsu0EDnTVFY3PHACu0U+h039RA4w6I9fZqvWdAQtrjxPESCn71
U0k9fARmTFKSqEgjnbh8FMwEJmLaTESi3znM/7l4hurWsYpedea6l0vsFuH2f62P
KZLEF6VZRFPutQtFIXVULiXljJJzhvxSSOzLviSYpX7LCjNXrHIanirLaQ46GSyq
TazGyEhmNJLTpi4uB7f25Umsr7K9bPkIrgrec4DPGd/f/SPvcmyCYSovsszZ4SaL
Ze5K2uCaWWUCBefpIycjsiB+9OnkAkIhbWnjd3yYp3jghG7W4zDFhDchjSrs1ilx
sXI2NIAf7jUSLrvA4XI/hR4K6AYgQhN10HZLVE3OMn7ZCEVvXUdYFDtv8OdzwCcj
1oC+4IYaC9hR7ywYp4E9TT/CvWqrBHdaOVFRQGX1i0Jn8sjqsO4cW8uGom+IFfCG
XikaTMMXSw9g97aHyy3GsDjKwVG2XEVIvCcFuJ01MmmjsMihtyBcoMiedsSHNYSi
3CDwt1VpPc2VkuISM+Br8Fn6k7VKHyPgougrkogxwpIMMwEIYYg3m9Voo5O+Xugd
Wbx0Z8Lyc623G2FlFwtiogklwGopXA6K1G2EX4ag2W1YvQZD5PdAxEjxvEyQNwrN
W5oDh1PvUTM1LGbSxEdl1IShpm12/GzSuYsfQr6t8EqaUPwvyLIj5hgIzFoESX01
CiKcPXgJLis+H5Z0v6ON3kWET28FKZXHwgjJKReACsK8IV6+EJbXTqnesjbUy0o8
Ri3GMJRzehC5BaEGhGkr+dhHU5AHyMsqBX9zWzP+bD1XFsXiGvSOAJBADcFpF032
yvSoaMSNWHPdYj9u9cSLVc47AugFH87lF2fYNo5Tuzoh6EexP/3qjqvEof5QIN8E
zXi9VFQgFZQ5YN39x9P7e/O7X6I1AA6jXMWkP8CIvjALZeAbtyplD8bS0agUNd3d
9lI4A61BjL8zNrruxA0NwoKPJJhJAF+KcFvll1qeW2tqzGJcvF8n+IBIfbcojL+S
qnHEsoGq9tleq6aGZwy6SoySyxTxugb3jJYCVrFYvWyTDbZEVV7PEg9/LGytTvFd
dR5AsTMCCb/2tIDGz0H+Ue5B6A5KSMe5rthH14VfvxGf5lVNadTLESUMjepQ0qeo
mB+Y4e2DfFHedneIHMMILobtd545ueR9vuw6C8+9o4CDY7SOMYTdz/KpScPArofB
8uX4xT/wyM6YBtMM1GirVPGVh7tOsqhYU0qFWiHHYquHFBDvB2v8VnsFxyhlGyEh
OevS9XWSKgdSfbJ1cs8IPxKB6K3HEnGuDP3+i6qGfKeiRntQURTsNlhkhXhgo2ER
Mvu7KBLcFf8qdQERyADYowozQg9XiyU9f5/Uc4YsxsTMqL4j/sM04BQdD2Ok/881
pIsQVIwtu2uBmc+fennPaeGUTmIFOGyGmWuc2qjUjoOQqov4IJNvDQDY/STdKL5H
4MiZ+vv1MqrlnpZx0SqLgAA4FJ3B2/RYsMH06cpTmeH/3k7tW4JaBwXpvs3q8ie+
nyxkkwJHcmrnH/zGQGvAKIx359tq/tbKCEiualIM0N5aveWWtNBAH3jDd4X6otM4
9AYU3Pgda0uorPFMsmo2ZgDQDaiXwLsE0eaJTnD4QV+ku1twZh8p+WVl6wr50HMU
9kdgD1DqJDRdzf+o6FM3cZMPztOLtQ6qj1Q5s5Fxv0tNR1p3IKoH7piB9PUoAeLa
QH//uLqk5XdRvW7DXBjYhtWVDdGyAfpVP1SK7SyFHXP+Gkd2C1Sljb/WWN8CQgur
UWhlFesb+jI24441TjRkoe1/m+AXKg5nI6oqsLEDIvDQvgzFTRaOMuqhpyqFcNFG
wcll9zvAnnKeKe9vYGFrmpVc6rydIIXzeLnVfJQn5EpEATA1XCUo1XTbcctkJ+Vk
Tr30eMvW98X3OWcNKZn8SdFTHfMr8cQyGkfCPIZJ+/97P1h8fjzrX/ToUTbkPURo
KLWLZyUqzM9w9UMcDONbiCb8ts80SaobXZs1UR4zHI12zx/wYHCbAgrBApls3eKJ
5lRMP1Fpac3B+yrMy6dN62DqcNR1RYNEn7QaBdHPJmFwYCxMHZYqxSHWPYHt8zvo
zW0JTkt7V3Q+nOGZbni1lO79+bMdZFD93CR/WeqKZZs4fEgXw7/VwOQyV6x9Yfkn
cOyT1r/9wJqW6SFHY9IT9+kJjXPACDvvgio9dUEAwrXo8OZiva9Ubulf/G2wEuaE
y+eOTtoi57JmNKfQ1KzzfEcK+/MTZeMUJ4rAbVJW384wWe1xm6lhskNHZBWUC+PH
D91+heTpUCuXX54Jeuap9I845qKz05oHlN4bEwzPycslB/ELVPzLTfYSEQ4tEvmY
Va0O00F//1K9kPeb6LOgXa2QvMcpzr8rEJB2jq4It9tRchGT0XjLeidvR55nfG3a
ElpZK3D2yZQTphOq6EQzjSuJDN3QVGxgOjSE/fCBWgf3WGJVL51THgGmFUhRkfxy
LGdaao91fXif9fcvNV4lTD/PwyF/EuwtKfFfVV+aY2Ua9AsaWGgLAg1MEei+oV4F
nQdnYHw7lN6X5isFZYpqsBBWmWbTIMMx1w7smg1M2q/BIO1tF0Jb0N7eDyhIaNzD
d/3OrWJHGWdqQpUnqykvNohevsxTL4C12C0yUvpakyaLNS999rMNn5k3N0rrpL8e
uXRkeC2jv86bySfds2YYQl9ev6ylb1yyuj4zblqXz5aDrhv6P2glsFkQ+6DVfHt+
NjG39Mb8n/deATXwmIfxxtrGxbC94pWULMf4lwLj11cEGNzP511O9nw37BibgMFd
l5Qe+yPFIjNOCTg3BEtmo8ICVKcwttjk93B1aoX3xGf2yfY6gsYZgPMBCP4nsozj
/Dun2bIgRCKac72Mx5VU44d/bkJVuTv7aYmqKjCRMeTCqcwf2jTTUhKnovVadqP6
DLxOOAQErG9bM6IJH8u1i87ZO8Duzmd7DYznMIqVTcqSSjiFoYmZilEhgZEvReqg
Qr0TGZKyUkRKRww6oJdWqvGnDAPcIE+PH8AJ5Bd893Ut8vQLrpff5LgNeZoRRRQ5
D52mBDLP8VYsoQQiZ91uMJxBaDVUnLhtgwmAkMuk3uaTF9fGfwMz6B+NK45DwUKD
250QWLGzE9vn70q6HAla2PZYqgQzZBZU0TX9unH7CF0u9J/i3W6VdFwseFKOx9pz
gJGctLAB991JdX4uEG74e8Lz3tywQ2+K3A4mp8iGAXZVhNukAwlnyyGP45DgaYTD
zzupZIj1d0AM4rhRg9tyLvOhgoJSngP7zeMIKIqIGBRk8LuMHKa4sw8U3xxWfVLy
utW3V3ymNVwCI+qD1YVoJqRQRjxI2//86LBTjm1f0kg+pv/pO1JuN2cp1zRRDmPW
IAAPxEsahBmOqHeiaKTCpTZ4aWmBwpfu6kuwYdp5Zc7hsCRsstEJAiLm9SJAQp07
ojhtayPHUkHL2suT3WGVNutYy9HCYE38BvWCeMG0xIE1F4MYOns4UJVXjaGDpoLx
yiIC16638EtdHbcZ7v6xk8VCu2ugqolt7cCZE8N8fpm8rKkpUuiQLtwKCPV3gt5m
uebzwFbObRpYtiP5mvFJbWo8siJSx+YKJL5DqM2ZDvuyzN3FQo51+YEICqUH+UA0
QE4ZaEp5Rsy/gqSFLx3MSp5LIJxtm4M1n+GPD6Jg2rhBOhsOjOobCO/KkFM7Yi0m
zWG2xvKkmmMOTAE9y7VV0XluxfQQJdRQy25mnficQSJJsocL1zmTqfzjF708W8FZ
8gCzPPfua+Ouas5iDyjutIGaK0PORpQ+Is/FYiR+Rt4nL0ZFlKNgzBpvIkPYIfKH
a39tGiPmeC33IvTELqkguESStQ9aIYNrmDefqnbyJ5mmg1jT/y+RcsUxnfOelJOA
kBCYTc//5gR+Lp8ATLg0tXZfGYZaH8rlTW0fN0Sqcf0UkfPL8/S5Ory6L4AwAPux
IVTcUgWnxkhqEiOD50peNJ5PnynO01QF/wRjBuaIR4Wt8LyZAD05+V6sFCWvJRFf
5vlfZrGivL4gpvw8ofBy8s5gqov236mK1vkSLi7IIwFceknwUCf8slbBd7EaQRNb
9i7F0++HrkMS0C0N88Ts0WCX7Lxs/MqyCXuF5A7jGJDcpmbh9IR9g6KhaIe7hD00
inMjMJ6f+X9J45MuKP+RLdril1LwVznfpcJofTX9ZzLBtnEmAAtWwerBQiUMQASk
b58j1A/JXVqnGssmENmOtwqoLDPWS2fP8/0dV4rEdmxbrknIk2KXp05GqUiMi607
En/PVAdGRKgoNiCU9sw7sG6vxqaisgkSKh7/1Iz88MCS++WeHeYuCdCAEJOkxTbx
vHP/5uCUJK1LvxpxaafTvOMW0K5Ha1I3lv3RKU/lZh7KcpNNgHSHQ4/rfQ1Ini0r
0sO/ov6l0YTrvjcC4u4T2M2ZGXyQyECKiljM8KNML31Q9skPBgRUV3N3P2PI3TPI
IKO3ULI0yl+1PZ3bteMbRgCfuPJqHlnrRmGZrGjUn6O4XuQmyKVaFyQ81ULyehXi
EQIhuGvOigukBT2I802DufJYAutkL44Itqsmr4sxlM2W3kr9yQVZPc6pEMPfxFGh
/jij5O4w3Ua4IE2+gtLV/c4ZRwGG0Jw9VvUGqbqPFhaADTOW9uqE5eiquXnlHwze
neoq5KfwgLPMGRBXVGpiweCVJVSnXDMcatZqDjeOangG4t4/2elvRipmq0QpkYeK
CZcWkvzovj1cxfxDEpB0T61R6buERepHvfGb8LL3FckA3cMzfCWUgecKE1eSGksK
hucsu37q9DpasPMebUf1Ku+X3G7McC6qBc1rUtYLsccuZk90vaibZ2qLLHJo8e7f
8mx9ObBOuvskE+hTkVkPzrkQ2TSknqwo/mJtCS9Jf8f5RthEjMYPsgMB6sHt2u+d
lMgVSxuSSuketnWSdrXX0YdWXagy8sHXxqFpe8vCjFkDRXTsZ+qCorB2+iqk2fU1
ks8yfuCfoNWpahry6dAS4cukxyfp5A8bKyqTucOJ9U3B+Vnev7tEdCg9wUHGVuB+
gasFinz8js+nz6z68t3JQ6NPipd/oklAp4M0BR2OfZlLyq2E837EZM5qv6GGXJ0S
nSoGo4VJNOcdfjYNpfn+VyrxBMDvmBvIBS9hjaBk8BXQjA9yMwAOuDjYEFY6JMLZ
sM/ok37n4lvftcrow3JUjvttafmcxDeUhuxfYbRaBXxpIIVNMa0aVoI74elZHyKe
UiJKvVeWzmF9c/alHIlyjUe2/c5JYR8kOVL8gbhHx5A80k1OwNH2IGMTLECnoHBR
mFL/WQ1sdOjnJD3IcCQb4XY9qxyelTnz7gtROfl1yUUoYus8HpTWrJDPs+mQAsUY
p8BJF+bug8NNDqShr74CoDAd2VG83u5GkJOfTZHePdqm5WWTSXD+xzTCdYtBcKfF
CGpP7SaohUmV9Drs5DcLuYMQ+IBPXdJKxpqDA1/N3uKQIkAx9hka6yB4SjYejuub
zkpgBMpP52nkGafQI7w243x8bIqnHVVACU+7JixFnCFFVBxK+K2LH5OnZ17wzYX6
tCJwC+wCF+DFx5xigzETjp7pzvFyjXxRPZOFC7oCFN5P1tsO3/F8+NBivixGpS9o
/nrvnf54CEltqm4zvZ8Opc+jlrv47cAgXjF6yp5J+jK9C2WNlQNTeoyfDcDvC9y1
SGO5v3rhOqDnQ0TgxnH4O+1QdU1Gt7YwqxL4JYKHobyZU2f2LZuu3IWhJdLptMTn
5VN9Vf9P7D5nVJBWLzS8CDDZZ5zkEDha8rIklJtWY64WWBjSDjcj8loBweMfTYKt
nEzEnflAPrjfhqjItet96zYvP2kqxa4PcnUpIZavDoc7lrqTS6qn3/GJ9lUCNY3d
K9BAaZ7qUU9qLrsErbkWWnuSpvKNBLYLvbtvwpIS7uCp1xULz6E9HmI7xR3rnxBu
atIP7epOSX6LiKsQIznoFCV9GqSzEeB0WbTI9q1kCgK/Y9TvtgKufYLF+/uivcH6
wU5C79gZgwoKJRZBOAclluQcyHy6LTp7ctnLA7jX6tvDMkc1zgil5td59hgZX20n
Mu8QkSupWJgzUBfJkMZSiAepXaGq5ac53pUocp3qYf6rYCzWdJCcYM6Y0JQWo3Je
w9k4eDj8c5BBePWX9ixXQsHw3jC3udnhBfe0PqDc6KlOzHHml+nEk4qiUNFTqXfe
ONneWhRzNDLpNSXF2nLqcZ9fTtJG5GddxB/FrMWOZYEQ8U/+3Vq7TY0prNSuXTmy
aOIE0sLabV5X0hETbd64DEjeaJmkggUawj2OtkUahDKSmdtbFwJcOzIMIIlmtRab
jAWuM3tZJcCyEbsQ8k5kRjNkzbLfdMlAsSZCrxlKJOw5Rc6hh/8riosEDnQ1Kfdt
KhXCG1K5+cIJiB42OdgvcaVQu9NoSnIctJV0HY+em/1n3giPjxUCPRnYmu1B4s/9
BRE0qPddQFFVS6bm+UGh44AePg2YAvapYSNvApF3F150ziuIxMzBMvFg2q7JJTTV
cHjwaLZNYbshP9oQ0s0EtC9q4+zB29M9iD3XipGFsoD++9Be/AdrUCOj/Lu3K3m4
5CcKsOBDzQsG7Dji2ZcjEOh4wIDaGKbji6ObwsOPnqebyqGKiey/cIuMJmnyqDt2
3m9MN8TIVuCOG/j/aBYyoCVShY8kH1dyHrEuzX4tI6Ual4vjfDgQFuq4N/URsdgR
8ll5XcaOaKf+CliwpykTVFk6I39EanyM6BbO+dPNWPmc0+QvkCVPxe6Kz3YZAW1h
GohG/K444ydg725F+pv0cQhiPkAT4n262JcbervvJiJjI+1pqumVD638/xxouvmW
4UC8QrOwuPy3YxkZUTCiCujqaSPeKvXlwduOS6xkWMjQI/K05DteO7X+wSSUyOdz
GU7yvb1cSQNN6tGgjA/F3P11IBP5783rC3nMnfVTF/4dbBLRLtc+mksIi7gaXniW
nd7YSbGxsIkwo6Ja2oYlDgyVCIFFOfQO7qtKSm67VczpIwsD6KfWJTk3aDhPoi0F
bU819V3NB93rkmg3bKG+yZ/QSd3eh2s/ShcD2263d481OuKX5Fn4SNoCtoe7obUF
Hun2gRYeg3m1nn2biv+dU3YuAqXYbC2YuG/QxfG5kGvgkvNTivwd0oezjO29JId3
JtIm0iVmwAZyOwEQ7lFWNkHT/VXHxVy0K60JhaFCg3a0GoOSeaA2m0ngYbEMt6nn
IAnX3llqVoc9fwcW+B86GmDlQktJnMd09GhrY8QG6swpRSSYjhgnz6ecGjSqVudu
bp3IBic4PRl19qtvryjgOGMCBWqpIswDYpN3o8P4eKyTcmeq5v+uHpT5G7KIIvnO
9A+FMPudRFfW/wJpCAqIuzlTYwjmdd9RFOe4ZAZIutJj9YqSmCEDMaLwozALSMMm
b6SuL2mdmYvvyFt59fqUv+dZk5H3+zy+oslt8Mpf79xnok6s+CzA8JgqrETNrx/P
/30jrAWtcLpvqPFQ01nZ+ddNGOgRJNxAQNS0F8kV6CVUuC2itFprW4g3xqk+z4jf
hu+Fa12zf+LhmQIXgiN8g/54fzoQvhI5/QCDkrSz7sI/ZPHeJWtL+mE6EZFTSCm3
4HAq0taD/O/rheuAbUikZ6B7e8L3NhAq5YJf7VTr1S1iERZH9gpluuZ83h6BjSxd
GgOQkd4h4Lbmze77/YgQT1Ss9QRadTIdAnLwTQXTnXWsDFVc2oLSChRjdRUlikGU
b+oZ213bb6jXR9hkhlyf7DJabDsmsxiyZPN9JJyNlt55HmZJgBQ5wVj212VYfIzh
QRVxYysgZNNertE2AKjkKxlLCWIreeggdIMdQbJV+Pfm4F01LcwUZUNohEs7qpzk
zD4Vfkf46u4WtT5uX5hWng3LTIHK8qnfQaOdTvbPtCdJxp9ftIrDdAq5w6D2mt48
buz2g998bSgqWwJDQxY/0q1gabdjwl9417z7/jaefeZHTrzOnyKAvyz1amtvQPbO
UuOIvZd5Ql4kQe21Gnjv7lfA7xdD/Qm2GedcRZN6EkrrbqQA9gY196SV6cC9eKmR
Kt2VHFGdksBKxj80RpdWpmAVeF2stEzXIIEl+Qs3o4BWLWTHCnQmH2el95subaOa
TXnwqzAexTPcIV9iHnwW3euZ5pFyo1cCr1pMkNZc3gBgJM5VKs5Ks5eoQeJtei4E
wW8vBsMkK7CZGYro6xpVv4s+xg1dhsftp+9mExOe0lggWuO5v8Hdp5Z/00xvPSTV
9NK2LuMH+IWKE0e3KeRVZ6fe0WSRhvmvLHghiOqoZwD4SyQvq0H+ajBscg05DKtC
m2Cuch0meBcIzocf3hvWHnoQIVta5t8sSjsmvwGzCuD7T7a6QB0datnAYAAR/auI
aSHPi90rCxSUqLZgV19l2bkW0n2Y+QW+wTOprMeLRJQB+mmpaX0YF3ewMsC6GszD
QuF9iAMt4MYIj75VRt1itgzkXhHgDjGxRCntF/rpHCL3wzgYlKnH4O/eZApPrfBq
kdk6fEQyze7TZ6w0o0CIp2kLBA4av09Lxs88ixsufEFFY+nTsbplAlPrqYIVZ2Gc
G3Nwggg+3C9Eti+GWZhxN3XYNn7wgB0a8czuqeFOP7HpWxErXdWLXT9Yea2b2MDP
fQ2QXQ7EsalkUC1PfeiR0R+x0WqLVdOOxMPJS/mTdnxyf4dbpk9SYKmQpY8RDBPU
WWFjPQ2kBDczPQBCRFey3slp1arBtTr7Eo7NGZrM35tqNKsDqvPlWCOK6a5bumwu
Dv0gDybMV0JcAu+3tePMdQXr9LcuT2viXgV4h3whfo3rDlXgzsg4qY/uahi5w0WN
svcbYhGgru3fY0VpaIclCty9Yu/INQr5HNzimVJvOgFn3hML9QE+/QdAzhmk92N3
+GdQXwjgNYrodfssIfX+JbnQwfRVS3jbGy5Fxt88LsiTdTBP9ZXuTVKqJVWY1HfD
DR46Zr0nstbjTOPnN/Do5qMYrAjpY30t71WiVhT1WiU1w2DzX5QjksJ5S2agKgSL
4Vihgeawy0TFD+4FuN07n6C4XrzP1BMVVoog4I/NzBBAP+7xMBJhbPOPqqYjhdiZ
tLeSJzAhmJBSMLEDgpfSISLVyGWZgTc61k9V3o7jCDrcZ80mcPQ9uFOKjehvdPGP
eX22K5Ak1ZVVzF3YozM088ingzouNUOrHibj5aV1iWeO9GizgOZKzErJ6NqcgUaa
9CY2zNnHj4NdqJ9Ep9MUAO1YKEYQ2WLY2n7/bpEX2+JqiH/a5ZT8HZPFeqOEhXyy
AeG7sqFSs8DBq4gsUycZnYZoCoGQhOwtCgD9FBO/3ZH7FB4niXLWajgE75q35/Nx
e1v7I8AF/OgXwDkrBUw3X7H919Sg2CDZRRIgP/Iu/9GQbllmBzK23Oqp93sxfrRE
6EM2feu2rq5JDbPAPaVZQmrTh8svZJy5QBVkSUit6busFoZp8nufKenpDQBkvV8t
a72Gh+fpwXkSpkU9ndL49GlO3fsWrcw9ha5iQqX/bjY/jUp7cbk7/8zrM+1pEcRs
ZdrdckyVTWrZAgBHet51MFSPjeFVsghCmsFwKcJEUj2qbHlDa5w0fMxl9SHSoELA
LfWwNx3FIgoPfgstRQlr7p4YpvuYxjc6nXsqWcj+sEQ1mbpPjQmh+iThX1UPXIHl
w6PkqFYA8fBcK65ic9ZyMkOh/oOqLoll6eMkr520N+ctTmiYZZhIuX1Vid3wXti+
Q35NcidnMQSpsfPvSfH6nRtmOJy/T8In4d44HSmOS96fgWMfG74KWgeM08k4H3gJ
vICKrI2Gz3NfIS7X+mIZ/AoUc5pal94th4w4iRDfx/RwT5wSH0PeMDCEn+IvicpW
JfrBkdTOhgibSKlq1OTi2E93dVP6/w2ztpOt5aHv5WVXM9YbSkrGS2jMIHZcMb6a
702fb2Xu5VPEs+W3IjBdkfmZXrkxxC2057PxblhAesJs+OzOvInsH0uoQdO8Y3np
H3yQyoHw1x7ULoA/BVU4eUuIv1Ft/foerRjmx8KBuSq9rpIikUo8cPPICCCx/6a0
oDB9WvctqhAhSkfXzR4W/kb65dSEDdfrzYabtZnGgK80qAdS0oXICknQ92ZmRZiu
CJeDM1/qV1iENs0+Rag8osX4uIZ77sjqTQ+SYJ8IhS/qXVDoIPWv+AL57LmH+WNw
A2L9iNwXJAFhQKvYlogC2psPw6wBTgACOiDRTHr+zuxOtxP5zUviEN07HS7oEuD7
9NRv8c2QARNhGfydTGoQUi1OOjo9LjSwhMYoq6EMcy5mP0iNr+eia1ScDDCPcvTB
FUJaffHXH6Bsyzg+vKKPwaM4KcolklF9f73FVTMMqZzW6jxoTE0mb/fSDZp1TSiI
BbkSbpws5xbCWoYlkOV9GaLc6a42d4oDO1PCFI1L+NLFKCDRNTbWp++ppkHm5NAI
mvVMQEsbLeT19SgJnAK25oSZsCBBB6IzUHIYFF9EFPeGRRivOk/BEf/fFHJK8Ygw
LmOtNYzU36QePRZPVzKJHlE1d2SmSBhqt3Bn+MFKudpgeMRl0rHdhDRg9vZ7+Pda
tyqGAfDTDcTiGraABJNOdRVWRIEWljNZZiTzKo63C0FXF3jEenEOZ7TOsippmmHI
aChlXYtDYwo4CGYlLO7ZzFZ3BsqSB3PtuhMPaIZTAIfXvPSUxs9RYjh1ClpGYkk5
ea9PpRFlDs8RpwchcVh09xbUftFcMG30Sv3McFYFzkkINXnkEpSyw2CcBiVpYpbc
/X62HlnNOJrkzY6wh+a8foRu6ajO+DuIMhBTfB14O7A8x7SA8y9rgnDieBInRYt2
MUakZw1NfrTXkXr+68iZfiYCwMu6tajQP1UNVDvSKNtVuFtG1icm6xeNf5UEgfIf
IA2Qv+afRTFN9oej6F8lrA3cDVdywmdom9Etzv1S/tOddQAzyxs2F1C7Es3M/JXG
dvqy9Abv47ZhZI9LjzXr/7m2z+eNSUK7JBxd5MM861JcYAHjMC47fWUC4xERnvVg
yCrppugbTi8SIjtKGRhN3j1RRjP2Gb26Py6vtVfsJn8lgYOe5qVmCCO6HVLy/bCT
6Gs7nDHTXeGddLlnvUqT7Q3ARGAacAMg9EfMvq2R131nyLgRoN2krTI0w+FQn/5n
+rARMIUWgHsy8VNWG6YTDqwX+ftQjk6ExeawhKfMllrqEed2eGy1XFicwodgQB4w
7rrWtjcLYxwvmezLx5WdWcosqlMWsapsCxSF93h7krqPjq4j65bML5Z3gxra/ZvL
5ZePdqYiTCmbxsFrTp85N8b/NNH7L9EOY7yZtYwynfF4/HFh4IWtNcAIvJmgl72T
aVnaRCdxao0e6GU3NForDpnGcbOZupxEeVYzOBRkrt5REP4TX+I266U5Fa6PMYPo
HYtVADKsMA4foT1IkdPsViQ0tqGnOblGRZ52Ii24FhEfDnK/6FoblJX22BaDS0fA
yDlPWqu2idOG5ASOqH/zGNUCWYawyqNxtRLl+R2snKnouLpl9hykFyVXTqQJchkl
bT0kl/0JSmXP3FZbIkiqR71lD7yavCIdm2ia9gBi6+sWOiYCtuTTxcpCXafsjecg
RBRfZGLdOyHbNxp6Goi8IiwjlCRvwyjiKfJiomCt1xzjIyYVY7nJUPZxWPIcoiM1
+x9XXwFLY27r64xUm1TYL4+3c7ZhZCIc8osufuJSC/NZn+tfkfDsb2k3H8fWMLnG
eBMX8Oh5Nl9bmN5hKkB30camYr18bvA6D/DRdp4HtzKCJ0E1rjq8HEXV4l0PoC5f
m8070GLLlBU3Ji2+Umnnd1N4osKgK9in1ThLZ7bd08nYLrBDHYGWF1PN/OnLYhPU
F2SJIjr84bdb1nemdDkoo7DWJiPp4GW1ZGvoT0q20no98sf5jP4bhkyyOks5s8W+
w1RfmkAzPNRoN1unerfpPV8KVOGlPr01IGuZYR5R6AUz0TyTVW9exAbs1Wan6fi8
jhKJtfyVyazuZRNLZ8Z0zBVRinXtVw2Tz7+La2MujjXnkfM1gU3371N7ZY0Wxsa1
FR3leRgE45K4NLmXkw1BClt9sRiSziFJPsmZ7PWjHWc9zt9EcliPoRoaupOgIP74
yMlcwx88oG+e+XWhWDtVTxjXFkUlbvts4bRNQUkVv+BvPg9AK3RStCWI7LeTpHCz
zccprgvrQf/izpJk3cd7KY6u2jvgNimO6KyvLcUyKl6u0X7zg4eA7bPmuUTWp7g+
RJC+MNBOyhL7jTtojLv7tRKEbxyG7qfhVa9phaWKrkr+UfS8YQZQ/7vXU+jmZiA4
sx2WbKw8HwpC5x7TyPtp5eYkaM+o3X0EjLqaoFfFUazRBAlcMS/TlIdmIZD/RAij
v0vhs/JwTtoT+SvST+d2GXOHHvbvNp40VSAXNrnapSDg15mP+CCYEbqJg1Ckzm69
zv9Lyg+PGf8xroel7vz9gJN7aC5EuQ+qSkNnxB2QSzSSaZ3WM8o8mbddMSjUJEDP
6CC2ASHOtB9j4FhrUdINGboY9QLajJdY395+oblq7Buwf7EuiK6Y9l2JkPO+cmyu
HIkQmm5W/GbRs8VdnoSpC6g+q98YXWr8yBsT4BpOhrbu+bex22uOxOn8Nx3iRPFk
HzxJ1AHXGYMveOGz2LoPYYv5eucbuMiH/X9gE9vcIceVcVJem6vBbf/NaCfH2yVM
Rd3+rcKcDsguDe3vuQgreTaTW7vtsIw/7Rz9bxNehugKOa/RNvc4cOxSbjjB54KY
MeHrkcHke+26/Wtxb88mG5F7Fq0zHux/Hgsp4xrJA4e59bqn62Ep1Jwzca7l2VO+
Myjcyk5AyenAqSzWbO9EfMVxwL2377x4Jd8VEtJ9vxQTsLECcu5Bi6dByUu4ojzf
Ntp1A++Bpqg9ZeQ0cCYo5MAB2FZGzYTSqEBIeN8sSL1DeNULMWYE+fyln/IQ3Z5w
pdHR0YiwQZDerHhvFl3PedtqhkVhzPz1U+0NcQr6AKLiBegM7ZYRcHSybo9h49r1
PPIV0lSEW5lcwAgwK1BvUByEoNA5cpD8syx3mNexzJMQfEIenP5NXQsKR0ZmQ/+t
ZEBAM9f8VvZX4lUPfmMyV0QRHkFF+llKhNTbkDU99N1TaZPzSOKeHoyTWTv+4ZI2
SCRqt6goaKJpQPI/E5XsUgHwFSlfalv8dcWkBPLeRDRotdobLYZ1dlfMx/zjHcC9
eXV+cfSwnJxpiW1Iu0PBvkcLQxfdglcvNjDa4gyp8d4JUaQ+EYyfak+302dxotyl
RmhoqmrqhSQBFwfswEOXVG4iHQGXu5BFbdsOe2Uk9G/53TIrq8ZaPBnKfofiuqP1
xf5hvPbAYDzgeyH2uvjaqc3AWsfQJQU8nSJevy6M7g3Vo8JxGKe6rQx84024x5cv
SMUeiIvDZCLlOkGznDUIPq2q1UwNd07Co5tC04N5PKkH5iXPh1QKVrG1B8R8O+V6
EI+XjdzOHtmQFTQzXxKEP3qNdLLIoPHeaWhM4pbpOVP7wHtSGwJO+Sz9ThM9EB8N
InuGC1K4aF5MgYn2GgTWVp1OBzNDQIANjOm2lZP9Qq3kx71v+hMtTu6CO2to6U4K
MK3rItOZeuuwFVkz/SgvzbhZ94nEfNueNRE6Atvx3eK24V08PG++ft24ihwZprGC
bzAQSrw1OXhx5jsf+zds2vuAGd3tO5NeNd09q5a028gxLaahIlV8k4IMcnwXaRi0
9tiJTnSioPwC/RL3vmXpB43HgXMKJNbJqeg6+d/+/F8+S0y7hNe1aJG1LpDZzV6T
MbKoSrVa9zcGKG/pS9DmRSE0hiG64UsNrl6bPSQ5DE5TUEDhcNiCHTDY581LPxVt
r6EPRfZ/BEcjE47MQx4co/mQpoPTKRp8RkBVZUmWcbSdclcsyk941wKD3QtK0bFU
qlBZ5VCovgOtQt2ajM4CHDR9ROkRQfvCsCu6hrSlzHxN4khgV5tHY6JZTJz42DPu
LuP+FRFjHGgUDomc++/784GJjgDg/N9MIcysjros7GTyHAcfEp+A6SQz/ESCBEMc
kEqoh+XQdINSe7ZsFDn6WaZk8AmcRDuKlOCSyr57mluB5DflrSsruNYrgsM6mJHn
G+ONPCDZHl3DVSUDsb4Bw5CNCdnvTPuI1QSMsKXUhCKdhsMuD3fwlFg3m4KT0qxz
zznfEFDR1Xt7ZlLoVeggp9k1p2/0PLobnPHWo3l0Q9pGgCNgWYlciN/BEfavdxh9
oYAgFy4KJamnadkewLERUX0etC0S2iqatbordwOe85IUTUNJOM07/fajcZ6Oj3H9
V26A8sEIvZkENTUFtvFxdPWs6ufAxIMlX3CeZZRINchf1vnZFiVVFXivQlTn1TPP
Um5fMYBff7B2dB0tE275PEScJxmAhrYQ4Bc+g/BsVzYYITJsJx3XUXG1X1NtmPPm
meS7hwP9N6ExejteuG31r9vKAjhrA7O0AiaUtNNHtScKDUj19x7fD3xqdN9540bm
MoGUnNUoOYq2EL4YI59zpkiCwg2fk0W1WpX9eJhtDeYROHhvsiWDs5qYuAKDBuh3
YCBkcfa6qK79YunQCjWQRRoEA0Ip/LOzpfvVOVRnXLF2JmP8WpT5i1I/GTl71QPg
jw1OkKKMZsHgMgR+MyXj/RbvYtaNSmBzK5Nds6E3CqU8Uo44c1btjDDkHty5KvS6
hE3BIAQJJqWhEhEEvzY6ytbGDCZBRnA1mvSSd9dTgwUFDSHLuLpFSD+u3txtbL/a
P8pHUYV9azU82c/X82Ul37ySzLMTnApXYYWTqVot1R0YERUK1k43cPlmaTgSY/Z3
vZcNRKlfzHYJz5V2fLWku9C3tORWSEAn0PWuB0x1ojnvr1VgZRs8+ddhEqz2SZm3
6dkGSPTDG1c61H1zd1Faq3O+buSjGRhr6zPhaz/xYWjUzhF6KmgN5UqKhfRO+bGm
COskVektU2bmgAlKPEWl0kwfJ3sNHm5ofICVcaTN4l4zlRwgNn9AuFWh8/7zLAPj
w5qrnVNkMBDZyZvWrSwLIhQWy/4gGNeDuXMwh1QfMtay3AMtuRJmJE5TECL1DxiI
RrI8Wrm2RDItDQQqryyoe18d8xJzgRyfX1zxL4XvKZZfEXVd9z+pgwgz9M3I+M8U
QLhVWdlT6ZH94DAfplTqZRR5W59NCpei0Lv3JpMUsWVZeqyLkdur2/X9eNwZNRR+
XZ0zpvrBgdg1+ablI6thh6QdVV9+okDGNGNMHCgoQ08eXP22Hlifc5UUSSf6Q0Z3
pLFI1v3NOoqCB/LwN4TAOMLghvMSoVHWOQ+3iQ/yChViYV+DFHKHK9oG0O9jwUSW
c90Fa+6s+TwsOgpa1b2Gx31HV35ggDDZPXaH5hlj6klaOnM7RSbKorEEfeN5eXXy
822nAvJTUYEzqcfeJCvXo2Tiwngq6OZNyMZPmislgrMInnhDiFpoFfdK4Dev27SF
IPoskFOznORfxFcZ2JGxR3eVckwvsKYE/Ywy+CJvZfW5ZTIX5Gbl1KyJIsmOyAg7
L9FdMaAztUf20SH+3iRKtsq9vo3PhJSgQn/Wh+HPpnyeJ5ooOzem0H8/Uuosd5LG
ccQX6mG9zcn8w1D18TMyBJtJfeC3VNO2LekaThUtJd2fKYbZ+p71VpWYrc0BnO2r
bcvsS4uGpR2Xslmu9yqT8kO0C1L24EklAOybBb5SyU0F8rq/U94hOoyvfsYjWNgK
64weYGb8TTnBHOw/xcoOPCJHpmC1OrRRAwjNfL55NtGoRNBsic+jWhXnbB3mXwHY
jeqphXBrz4Jyh1kjQfkqiLAz5iKDFACKTO1Mt/r0KZTFZXP7/7Q5He8hNkesPLDU
m+tL3AIGJZj0EVLPGzv5nIdU2n3+hp0ZMHGh+reki0vok97vXXtCR8zf19YU5Hp3
5scoh7vcVIwnENpZHBSUv49dO6AvVAIGKBD9dOQftyrTPooThMjUFB0W5m4iyQ3b
nceyBup5uwNY+ka9JoUEKtO2VvXM11VxCOo0zPmxP69Ocs2JKfeWz5SIVOuUlcoa
kfytQAJNTOxmvDnS2N6iGHPhqzOR8QhcrAnuwP+9IzejMY6RqUrmgDal8cniw8Oo
Y+z+NYtGzkBxinyHs6FPMlyKT7l2P5OJWbY+RvuVIHvLtnWoRWyCFteGcD3zNbAH
To80uZdpmKdnP/nFV2jaziHykKJrXZB70SsfxeahJib8ObqZN8pZgzvUCIdJQyXX
sYEU/7116Exx7TxnQI2+RNeiq14m4mnIzvFykIpmHkv2itWzuw8u4emQUF6UaePg
TQvcgL5+u6//T6rlzVXtCUqISZJN3JBGyROr8vsihsKouK21h+9RYZngpGP65S+L
E/h1u5vCr6nYPB0F4/i2sjBSZzTOaSs1QuZfBbOL0Uvvn2qNQyvZJ11Qt5EClNdC
6LYrqwTUL634wZDBJZX2Zhc2FcXdHpYw0evZrzOuArs2ARTA8vqGp4ySgm1mebfJ
9Rx9kISLmcQ/OLJJSUfSxLXtEFKhGJNWiz66iTefoZNU7egt9H5dXoB+rPIIrnCl
J4OZwhjxzpCCLst3Mgp+xC5MM9Ph8gC0h4QicTZZ8QEducVnWrWcXCyrrzPn9dKt
n7yj6zrvTHG8jbyyGNpcMZczBaFQhqanUrr8IdGycNVAQ7Ep640mzQLW1KLgZN+N
tIUHiPeH/zuy5Bs5LxDUc/FZOjIvr8gh3/yUgy2bvLAo4YPGigYwxvlpseE+M1ai
5OtBz35DQ5mDnfFnc6owaXJ5yrqouhUAxDRy6hUr3rFyPsZp3ysJ3YyGtgUYYV7n
QvUihXd78yMSWuP+QUaD8+c2+djV7Ey8Igx8TyGLUte6HFEE0fDEgqF43wu3LkMg
/sDYWjDvysNJzuUMfjKnXBrmkiYESV152Bg8Ooj18bS2Oii2ihPOT+OTNHfRtavu
zDfUrhl0k+CmME3HKp3o4vl7XJFVhBc0ab2fhKOnJhwgs5SpI5TcHY9uAD+BAEF/
xv1klhyLH8oOrOLwVnU/8ojSx5yTCdMOgcZ6pxF904wUBKHuLRLVQxQoNwRp/v95
Z6eBMqguZqVgTUgNqP8HsFsKl3b8VEhj8g2gxpJsBOktZGZaY9dMc6fGWdY0knQg
6i1UfI3Tu5tH/PRPdUe3S52ae7f8MM1dv+HNKPBmBRVuF0lBypV5lorFO20YsND6
KNSxWKdwXkro3yWRoBfOEDDb5PwW8+L6M6ugiZb+V2XECVXe0MHct9txwL/M1XUG
MYwfOEc8aumbtdSQq+Q/tINd5xn5SkPCkZ/afEGjr7xgDyNcNjxmHssT6yvU+0y1
OxE51u5E9pAHGKzwW00K/TydNd5mN063juk/27JMNvez+iYCmyeCIzTJd9AhPAOc
xLQUE1KVZDPabNGp9N76pkAsVEy3YIhVN0JloagWCCSCmZAu0Q9FAumuw615sg+H
VmwPgwkGvSH+L+DIjflGF/4Xa+HQumFe0Q+Sx09wOzvI6CJUjesV2bNDstg1chLK
gjEeiZ48bhE0EauvcgECCVlTSbn9vZdtz7nsOr+iMu90lPdpn5OAMDoPQ05LHAwk
BRN/vPSNYtsCTSaQjxZLNQqOsSqrrL2n5tDHUqj8ZTVIvQTY8LOEpYsavRmRy5oY
/DE4FgJF+AviEZiN+5cRVCBiLVF8VpU2thq7WFS+KQiukl2ROzYeffSr8r/tGQSD
/u6Dy/visI4sbWOs1CnUMuGoh/RlfX1+8aL8Fe01uz6SSA5kOtpvkazyVEh+oikT
ixTpPpakW4I3Ip/80mLaJa9JEyyPmj6sGrdKNP33VL9G4VqalMLDp1VYSep1rIJ9
g5nowzhurdI1jSN3Zwi/6jdPVdROpFdAWTasKsL75Jk8FZmyf7uLIW7B6Hqz9mFK
70JHkR6HXT5pwCTFlaVGXzJIkG9rYWD5phuBiMtdEPkcZW38CrbrI9N1ZbtrzUHi
uiI/tztyorWXEcsaJZQeN6gul3tlNeE62fDnT5XnAGWr7BfoDImZ2W3pwEZnAnqd
+jzjAUTyrldNmUrx8snMw4uptoUGA0AbsAmv92ifjlaT/3pJAWNCLyuWIL/iPnCp
F1LoWFREppkFyVdQmheL+RI9Ws/OO4e/fTs+toGcn6Q2K43biW/lEEe7jdQ1noWW
ls4sPQRXO+bCJF/4e8Kp38v6C+lujslys4F4KYOIBXeTXV/onL/NEMgPUA+4Yxe9
bkov9Nw1XNwlYtwwQRQcum76a6KVfAIbVVuLvaTEPoro93SlGkCHZsYsF2IN9Ssm
esB3B1fcrDjFKGQuljeMefOLjWzFyYy9FRe3W3d41xKt/KrefFBSjP+v1Sxux128
jcUQXWRaMVQeeksY+lJu7aryuV+beHodAq8Mcx/Dccs7ocoaAULL2lWcFjWXIrtZ
V86CzO2kiJVvop/gSejWNOxBtxb0xMGvFj/09rdtF/8S/5hUnFYIJmjI5uaW+yVs
AgR2x1qWMJiemrZPnaDOHYmIPBAbMEKtmS3xD19wWVU8MsONwVaP5QhY/OFCD8yO
MybWuLGRGuCKdIMk/nYHOxsaBwVNo2WTEP5afXm4munjd/8ZY5bNPP71D0IRTK/0
+vT/qRhhrv+9VhN4g5QKBtAmGUPZbIxRL0DvjlCxRft+PRfCFv+PRZXTLKWZKNzs
+m7j9X7as5ufdPJgb/Typr7s4a96M7k3e0lFLt+HGSbJuDn/Zggjr/HWfyIR/Q9L
8N8+IRSqCiESWYdhEynwTdNmyU5oX9iU4xTwd0KYEoRrfdrLsyXixAoCPK1jKarr
Ip7/YzwEKoC//lfAk3RQhlYPPKK2iP2y2paGNCJVsvILzhNGp4v3D2gTpvMgQKK2
WTAPfxbDQ7CpN5O48hxsI5ZZ68yLvtbjC8nh6pG9uce74PzouDYPzJnb6jfZ3AAf
15VdGOlqJriXxnpAWPIJsCHzhlStAwQ8yWdAeokYbmlxwFkhx7/zKZ19sdLnyJmi
Ck6dJIVGg20/F0UNtbV8bMvTOObgLGj4Wx8iibG09Lka2uKLMTq3M/CoGQh38oTx
CgSZhDNnCk5YAwEGNvgsIEbNUzqdsRgKcjzVW1aCwbEb7JqvpvqX3HSsloyqAbZ9
vLnlkfovmY5mCFkFWaA/hzicMCDdUZrft903KV/C9M/AXPga+G/aUUDQFAlzclzh
gUyaNlfbhA8fvTD+MLXSVhPtV+vpp8Bvf10N/m8ASWu8USvg4FRK+HYK2JDh4PlJ
ne971SQFoJ/TGf0BtejNKIxBIn7h1tX63qf+94IGgEg3jOOasqqgvvSZCAl7U/oh
bUecEcaFUUz5YiMLxmz7dRFx9A8ZGA4pV1/T/o8di1pyGNjwRUs+7OEtJhgFQz2v
9omRziT459++cPzuRu/VGeke6AEiBNGl4okAQ5LaIkbtuWmSlUmYwyGeVpexAk5t
OZC/hQa8dykKehPhiuubhaCfPzfNGOj4x80dgUjFJZiV9hw2r6DAY0le829oKzqx
D0wxk+/0dNgtDEJ7EnazDY8jytAIlkmNWsuCioD6cYqi5HWh7W6JguPLVLWG+Vlm
b9uBr8Kb/lqyWjCSWjdyava9Fz9V5jVEGf39CmV3Io6W/pCOGviY5Gcvx9yLXQRp
sIIRvQWoB+4n1mEh+7ozxjL256Isd8KnKHiC9om1zfjB7on0Zr6AEsPODBdOMrkQ
mUN/FDNNpUs4z5InMSGrfe/VmQasO3ySru9VAwrXnZMBIbQNDbin+Z4KBhDgS0c2
xO0qZgR3ZRckhG75Mo46Hb94dx2iSkjF0jNlCyPFqrLty9YEIBLo2b+e3HPiQKZZ
7nmHLVgbStOLQ1ickbaqr5YSQUrT9PXp7AOX6vGHesSMfYFLm61ALseZz7QqRVbj
6+ep8TKoSGGHJrp7wUkU5Ze6IyB25CmfPV0HVolcJOVSxQmj+DBVoE9o1vyLmId9
xub3AOoHGgCm4CGMcTSCswE/fMusGrNBd0ZraTx7JuXvIvPXMA5MkVfqZpM6Lwmc
plJ2XixVsBOjkJ4Bzw/c92Tpk19GTUIY+kx5UsQGD0MWcvgksglLWY8uuWGmsDS4
K3YxiJY9Is0Phdqjz9i9LcMBb/NRf1GN6j+5GJKHzwZrRbM222h6IJBP6axCnAbh
DBVM9rtxceHn1xwSwAJzGEAeg1dWEP+45Np6+QRmW4AC1uHWVDt77bBp/LGO2h1u
0jvlfm+MRz5Ijp9SdKVVje0V29j5hog3rQopBoOFPipuNNd3h5+R9qBmmvY5+DoI
vb1e3qAg17dapRnfmM83N2aOS9fF+1QiagPqg6oNTUERqdiXNsmyAy7ISA8acXNx
m5e3+FR9yA0NX7oryKkqrw2Kzz6o5rmB6V3EXptrUr0+vWjYbo/4gu97i/ejGJ2d
G/TGAXldDoGTLJq1lOhEhHeO68Vx0bj3yl3gLZqjvq4BCHZYpnZG2hs21D69CR5x
uLPf0WR90VccAAvZXmRM0Fe06H+ApaV5UOXA4MLMaICE7tTRanQBzdOHJrYQFCqs
xDfEN0Pj+yMXTi94KIk5DiEhScPNOZzCxTGkrtxqAsLrWdmhy4Zd+h17s7N3viol
KThs0VdrMChA2dyi6qVjVcBF7N1rpAIe2si0vyDg5+IxPzGLut0Zge/cBIAWBtHO
Brl8AR2GM8JN2ODFggwna0AQ8OqdjWFdrtpPmIyxCNKNprA4lV7C3Q8mZGY+hEDo
UCKPemqWmR+m2c8VcksHn+Fsbfq7zsh7R+wJj5f2dMS0mDVsvBSDHzylAlo8P83W
UAC7n5aIubAsXy5zS8G8CQweZbbPtaSXP4AJmG3XjjCn5GOCFGWZ8V+WrlCVQdzE
ziBLCzV9eknal4FRs9fc/yzoBTi7PW0g5BeE4/h0EOcRdOCdS6TsCzrzFkXbUFl4
ElTWSRD6YLT5rI5CRAzW4FavkHMXhd2FojLZklInq2+71zhDu0ivJTGy3ewIgaRm
SIGmdj+IosA4hN7Tpn+vpv0hLKbbfaz6VWe/4jw2cAgkwSzNt5vPOIEOg88PhYv6
lsziuUVvDJIK3m27FnpxoqAJrhT1nGmK7J9AWST1uldRcQoN6pZe+HDyrETF6+Ce
lNv/VNV8YMdIayuWDZ7v1wBJnu8O1usHrsLx/FEZbq2XpwLvEUqOsbsK6pTYhQMi
AM/U7Szx7tVKwPLNltubKViOwYv4k2mGNQpbFtp0w32JrIV7MO+PGt0Er15sWr+O
Oo9PMOja5LNQhvkjF4LzGKYfvhO2nm9DeJBHHY+0Ldv57a6O6D1ZSx1WwkTrszK9
EmM9w1MPyTI71Uxi2A9JIsXLGU8TCBo82cS+Y10Upz/mkBAO/NV3Nh2c+BQzWhXs
KTqiAFLL2LlmLiUHzYHqjyM7nBqkdbzv5pE9BMAnlnxUh7qumCfpMFgLOVO2jHq5
Lst7+DGT6qmTro/RV7r5oWQ0hB0em4hjBVpJvGzGAcKtfVGyD1kN8j3EOYRCWDPC
M804UFwiqh/W2/aCDwaJlU2p7p2Bq5Cxi+IVx2GGYycka2tV133dlgDtBrsJHJEF
9ygl5vinb+FKvGugX7bvEa0E32sJM7DBlufbz2cVAWMy3jKUbWIorJaM3ubolcBf
z7IiDEJxCmhxF2aDQ29Q5/Y1bK0Hc6UxK4CAI24J71L+qJKxZFjQtBy8Cu9rLzWW
69C4CETL23Xyd24LsvfHtuhY2a3Acc7QPdXTKoQZqXJcs/AMt5nbUsScED0yV9hb
tcl/RV69vkp5tuKqj3aCgKQpa8fTe5xVJ2M5hy3tDJ9CjCY/Sm7Dh1KCFpI9uL+Q
62GtojfUi+qsfukx6aMvucQPmrchTl58vPyi8JJMAkdnuIkaROAEVCH77U+wCnoh
rfQb/JpmwzrtTt5kxeISsT0YaM6dULYXSfljxxqztasH38+QNZoJWMSdpriKqo5j
Fs0bLieOrBqDsqMzuUXszdJEeg14p85+8X/wfXWh48h/MoFl00Bzu5rVeen8Mvpu
s7Q9tBPTlHGIcmRj1RBnIjz86MRvYWFP580ygdnL1kTtz4EWqzL7czhX2+rufoov
2JUpzrufVfCtWC471163Nl0BuXbMIHbMcnvzwXTX3vmUvnVWheYSw7ZKVVk4SNY3
qqVgtb1cHRIWz1ff6xUzyelBdCAFqRGkkLBlYy6uzRKxVtM9sLZh1n+uJKIFDP51
GRNGuViaMRTEh47syceITVWe64BJtDfdfJw/ZIEid7ecqrB3Gx282cd6Sq8UyeBG
H3gSyP/dv61E66xqn5/ugT9O2S4RaR/Ntk/HGrxV3YJq0gSVq1NzDr5dsUsReBtp
HgzpyfmcTrkpc6WU20YJsCd6As2/QE29sAzUblSCyultaVZdDa3vilSpkAqnl40x
MRLN6ILG/6iWWloz/UOz0HEJ7D3/rfJeHDiMp0kfiTfrCIPKJlDpcB0+YgN6ahM+
yk6S25D43Fz0AjwN8kBZx0GKJIdVy0sw8Q1gJ9Q7UsSY3MnQ/DwjyQCBSIDZFoq/
L7FCTSp0AvNFkoH7EpMwhtGgzZ3VKqA+UkOdzJ6XHsamWmz+BAwb7S61TEFx0r7Q
4vPqu8X4Lue2vTIOevATkJbZ2Mr51v26VlV5u8YARKMxVAmeW//A39mAOK4ZB9d1
R3WVvjVdQ2FXOM9T8vdnZxA14PEm3W+QHH1QmyK4FmBdVmSYUsc/lUV8RNjB47uk
aPqeNfhW24AUQgEsK+fdETXkWfQnJmMrYKygv/buU3uNTFpb7bqzQqnCA3sg1hYY
MrJoCXd1Za9IqUjkFDKQADkPa1buu9Jd6MbkdfiNGrC0huKPmo8pUrjvDIJ/eHBo
lJOaQn/ArVuVaZ7P4rSturX4duT+jQ5N8xQQMPATOccBCd0mGhMydxX+UnJ5mG2Q
4QB7oiIWcOsoOc1ZEd8N1C8Fs7a+yBN4XO4TJwMvcGPJy/774+2vB90DFFwhwq+/
92sn9zhIVZva+0SGYk/+gCuSsauXtZfJ53DxMhUbJJ29olp7D5gNCMVQx1GA0+Yi
Vr/kG+hka6DfUd/+7hKFqYnWs/rLPYtoM68O6L63xaoguaxRhM5slmpYC4C1kYeV
+yafq/fKb/fjzoprMwU0fQfXoIDb2n47kbe5GOOEKiIyGZTXBxLz8efxjgYvVjdm
r8iwva0o/FVDYAqzYFbHASraumUMcYQlY4ZsR1iNBAMcvqHdX/KsYlNZndKhgzMI
ElPBOYoC1VBJVIeA5iA1C5C5j+nmBZ8H57d0X+QgRHAiAVA1w4Y6I2XGMampIPrw
Fzwz/FNSzun+ZeqIROjAlSE+N3nt8y+FejpAqRhpVVdJEvq5yduMqidCt+rvUATH
JQgg4mzJkzyr0gVMOtvaa4uEqEEItPJN+VYsCjgJPfYSDJyQ9lTtQ67SvVpN9d/b
Z5EP0Q+aIeb1ipw1uk8rSYYawDGiKcLwYIQOUAschqXfyRdI7HmzL5VF+XAVKjRA
BjPHsBga/697MufPdjGNGkQSbLi8FMenytBYul7gGZRGv7Ff3gyA/F5eulosYlay
tvthj5pgYUC/KmNtehj7zzuZJ/k5nhrWpSsDGQYg4XXT5y48klVlSPVXbrwecZlI
lSUTTddTzHNLqIpCO3g5VXcu7fa9UhnWiAN4gXY8en9+zaN22TecgPd5BrFaNrkx
erFa3qzpGy4Ohb5/emHV5xkm4lHivFgDjgxVSnHx4oue6jKD7DNP43wiLmpOGOpa
9MNNqFIZkU0zzU4JZLsw6gdHynHNl9578BwGHVUoX+sDtmrTob+Zxe/UOB8EfIoI
Zqi/HdZIL4/tQ5YzHPWwHeySWc8wxw3ve7sbeflYRZ8N8cGDn2iFP5w3whQGzNYb
Ctp/J6+CNoYHIjBnwB6Ywc/2qasLJyw+LFVJRRqzB66TwuokNWmnXSg4F8i1R/YF
+RMdXD2hcgAvzA8Hn053B7u2bUSOhb48F3T3XSt8ELLNnRwZA8P+2tC4TeAW+10a
M1dg0hk5pQpvAabJYxGTWY5a76vMUmmoy5KrZXyhuzWGKEbniyoClfqajw8zmU+Q
DP1lxCr2mCKfIRMX8rXdrdVAlwkrKL69/JvMCXoeANxH9/cUXuK7RcGIfp6S+pF/
CzCWdy1dPZdLZgXGeydk88qEw5Pi3vcCW9UkyMIumIvB4qFZSrD6BmJUA8Fq99T9
zeLM502SebrM/4+sNzsiMpLX5nvS+SiwDrHsGOYT7myAS+LU+pFiD7smC65TvPtJ
PnrMOPM8WdEzbXgMmAyS0QlUw1XERpzf2/QjKRATvLnfN9QVuRmUDdmZIcRDkOXJ
lvMSU5A7DV/mFLapPBqNk4KXugG+pfPPastZQVEASrcEGH5OoW2N+f1ndYB8nsUq
l/MnCppTevL90npf5QN6ajK89w86Vafub990iizmQ3H+brl0FJOcwNV6loNtiEwA
ckO+82CWLAT0R62ifDKHS8UphMnT4qLrmDz8GSgqnqupKsvQaH99dyuB5v374Tjt
UjikHhJVk4BfkfX0SInssYHzUoWG+XfMFk8SpH37TuHi8tXgGup2blzOUy1Hiznd
EPXaosG262KUucPv+StQ3QG7JBWvgTLnMmYK7VrLQ6jlccDJMg6pKEOvGAbgnrXS
lDz7yzM6rfWg9b3MLkdLtNy+nsi5aobpKC/lFw/X+A0hztV05USwsnNtKnNv2/zC
e6KVR99D7e/AdYEv8pOmeyvX5Z2MpUt+St0iJCf7y37RSZdoZq/+XM4VoOKHB6Z9
G6XKZap3senU+QFiqPljVi4L2+4ZD6ezRSO4WCfUBmFzpsuLgWRy+IWSE7czyndf
AknvF7J+cvqXf+8VC5BpqcBU/FH0vKuJVOlnSUYthsTrqWqycqFe5xqqLlJuELAA
X0xxCZ3xCleBwRz+YQacp7jt9qMztm1eI0Bxjnt52ZziNSJIlLXeaeU2BX1/u9rF
5zalH5sRxFB0gjp+6Zcn8gRiTCBwmRgQeuFnt3X5rdZHH7Cq3kTW13YsdmdQcM4e
RUc4itI0cWaH9ZGxCclEA18DdIMp8P1BW4oN7CXr0vbShNfN58sBfRmGIaP0kh+L
3ojrsu449b45YjAe0nyCjxtZ/Gw0zDfWQ58t7uWDTPkVFHjVDkQbI+QZWOX7Zwjl
RSyRxeHJ8MDG8QPV9upIt5ERkoIDuiz5YbEG0acx9EOT1mXZWdFZsmh5fka5S2HC
uFDQBq5+vtiSlvCQvEGWSM/jGGMwF3ZrhcDkaMcXJR05+hcGQoINIFNLSm+/MH4s
dOASLiShVwmTQQmwhsmp2iObvKdhZFRSCrd5uk97+yKDekZEpEG2nPpmPyTv7mM9
UZHWUt35mmOJkUsDaeYl0QKPTyT3X2de0KlWE+p5YouhteFBXSJyzlNs+IA+7vK0
2q689nEQDqSzYcznVJjxar2QfcqqKio36v/BeGQQmz9NGombgYnKW7MMFB88M6F8
9KVb2Em20Vr18oMETq6MSm9JOYwaBmwtcRiw9T9IdB1jc7qJ9E/cjRHDlEjHh39d
A1PC7uKzW+dwJK25q1VgCl4Qxhrdvq02IMGYMEHyF3j0sGSl8MMrboltBvOF0ptP
4CNl4Vb3DSZ9N6qFHDSut4sdnGyMueaO7Yo2nKsjzXxQSZIwNMwGCu953SPAE1lp
hf4elyDlrSNA3IyUZFiFcLBDEcpV0XpXgcbK3Gb/+OzaQtA9++5kqB7DN0QLwvVm
NNKmL9+1NgfXPjZjOvfZZ05zEuCgESft63W3WHS46DYkgGdQqRy3UKRpi12KuQBH
6dHtWLqhvXdkvMGorYSgR0V06g1jComQ6u6YmXTWpvftvaTF6huzqzrkg9FFWWzP
7UnGMDnbmmywEOGVilf4cNKKbDdBAHBIJ99NSks53/l7scYElbrDnH5U36KRyvfF
ACIZTtTTKxeHe7ivfJ23vmhaIiUsuO765QwOLZC3An2pIILRN2Wr/aDKf8r4YvFY
pgVGi8P67Gr7eXwnj3aC9Dt3VShfHoNFqMQ7hvZe/SyPltw9xzz0m463Ukfw7uo/
5dxFKKQEBt/uiHGULO05ayntzemb4JZNDTHXPd+bhDy5g/Yor3r4FtajfZ4lPA4m
6RB6tkTdrDXL5NikIL/ktP1Ybn1/DN1k6si0cGxNkzlo6TVwsRtNZSPNHw4qXU7K
rmTJuM7WeGVE5Y8Ohh5BNzvdZT+LCBhqTQCTdlEyItJx+BPePIrFF7UZKOnU/8kq
PvLytxfpBqFCV3iIiPkEqGOxNuPWdDB+ENiaMNLFYGCM21LF0uhYT3ziTiCbVFk1
mHDLvNd+cDAqcjewyo0ofbzV0bJN6urAyv9PSWJLDrZ5/+1yxGWPr/n5wswJ3XHm
QyzFwFI3A1nDYQuPURo6qCkianuMyPl7bg1QVIgKE+PL9M1KSmAoLyOFZg0rAN64
gG7Y4+HVHxV5MRvuj4N4c40myB484++e8dMe5rhBI5Ux5PqVC32RQ8fveKMo9nf0
VK62GVI55rqs+mggVKLcbIssX99kLqOkhSLE2aZ4xOIR4zGV86dK/zWNKzr418Ir
H2ad3/y/oNoVzt18QfTVx2tY+qabh2cwULb2py7bf6vpBKu4Umj5iORrd2Q5/b4H
mWAP3wZA6fQHt47fDeICUC1QBXRxEWsxqwTnVoqRqov+bwKbm+gQjMSrA0CyBzkZ
nchk1KArJr/JQlFGiqaJVn6J3Nim/RDG2Q+UxwUGYHuq76kELMWXreV7Bve66SgT
Reiisx1TER+vqZ1zN0J3iGxLhe24EXhA5dK4TtgLCncHcnx1G3RiuKigC2fZvufx
q3fAZ3GkCgqS07tnq0anmy+aamokTcG31tFrlXZLHjZaRoPYBkVtOroE00eOtZvp
XNo8RvFbFiS79ouW9Nh6DZs0H8uGl/XPNSggkzc98AEaNwOL5sR/F1LPh7ClXRz7
ZhM4MrBVwhvZ5AXYFPmddc0GMm1ef7FYQJDogEfbOkdP+sx1+dpSWz3S+gkluZDN
EW28rcG6g3Im7easjHuyR1TYqQktNe9YKhVkCjD5thOCKgD+NWd8LQ0VomjeuiEY
SrGla1Wfq0H6lb2VZcs27j11oL5hBUbZXIxQx0j3nPf321sS0vYip+oMAxB4lHsV
O7OCC400h7mtwLYA5dhJ/YAkhJhHWhyLdPGpAbCRfzlxbtjVX0pj2yJUGwJ6BjUz
JOSw1tSAZHDF66igI3cuuqWtuRqMVm1G7Q0X5oPO4KPKA0eyslGMX4YiwKCt2b6J
laGkGomRiVpwj/Vtl3D6LXqJ1CWZ4R33DEvUPHHN4i3IY5B6AIokx/kW0yWqXlS8
L5Gv6bB4Vic08rqSbFBxipbYZi17EN78Q2t1evoTHEapc4dgtjwE/dKgDffrrkPr
Oq+9DOEo3i0ukS8GVnG3159bZaYMkC80vSAJwiml1f+8HdUaTiLF7lhGICbLjfqE
mKTlME3uh/Z/NSz26Ly9PHp23d3M/8mMVzHM1E33Ak46qZHc7LZ+IZVacdXmRBOd
HraA9Iz/sQ0/E+3w8/wtWjHAWFH1YZ3gCBnAyMspXPQAdXbdR3x93IGCTV/xnC76
N0AEF7cwx7lc12C2UurULCOVu9xlhxM2WtazLC0JR60a/RSygKTzhanpFPu0UnFu
CusqSppKzmwDw3SxbZ5fmfmPBk8eba6u6ambK3EsoNqBzZIIBmh0sFq2H6Un+WS5
VpyCVkJ+TujwRcqFDtIaq1o26NMzAV17bFu5SEgcXKjpUfssf5ZrjSOvci5H0p7T
CKHOB20CLpZhxatP4fCrKkVkGGyGIHM8QRwjMCJL10QQYRgAAzA08YINeznopisR
A0KKIkAclXCKgWERVb0um0rFc0hzVv9rPSdzj5Uy7SHceBKXw2rPCfsoesH0UG/X
NagssIqmzHmcTEmvwLTc/n+MC0ouac1Rfk063pMOUk1CBWzGnfemPEd0X69SpUZi
N6SNrp/Y/3FTK+falA8h2kMmXFVsci331JGg156Y+3wrluWQjEZhoLdwZHnfiKHY
GHpKDmIXxhTLs9viuaJxFpfe1G3bjlCuLbpkCFqa/eItlL3CHiGYwsxLhybNS2ME
i9WxjK2P7V5H6ykcQViBQWVdEQA8zRV9gRvbRjWu1NmEiGXmgQI/nv7NW3ltJ9us
HtUKvCB9VYFQaAIM4Hl93k9NSHdya3siVtlWCHLLhWVhja2jkBLqPtI9+CF9RhsK
SMoEBKjpij2sVdFyTDAILdWt0gckplNcy5iiQRXtqVCgjgV7edLys+NYPqthH7Te
YZACvjdpSd2IZ1YiPUPAI11qxVyNuiXFGeLuGC51RXYc4O7IijSgKyEdRF0/PUK3
p7FlUZeBeQUX+ZUsFzWnc8NxHpaxPQAuIM8GZVw8cPVbpMjwp7Hc1R1SEhLu43xn
fb6Fh2zP04X4kVBoZiFW1HzeUGWvMzE853AfxcuZJySmzglLehRdQCl8TsJy7YjW
uPLGXz1/kjtgIxAd1UGiRxEliJJ7VfwPnwDqMOcWUD/T91PeJpIYfkRppJk785GG
eiJOJ0hHILG6qIKYEqsSmg58tySHvTQjoR4ezh1nq62QrfozoDA9CR7SN1Yuhdua
lLMHMUUQL1kiZDFbYppfQ4JV63Or60VOcSrtlMbADxNZyMKNQXhb7v4XtX04166Q
FWM2Ev+/0pNfwOR5Ef0EJ2jrAU3qDJoDKOonP0GELaMZ5qt9Yco9U0mxU7XA7nP/
35//A6tPz8pCDMAbV5nVNP0ydU1P3seGi4CGRqu4hxToCnsedsSGy+kRjzlSVD8p
3ESvRP/No8jwtePQ3syzQiBABMCJ+o5judFYUPgJFuqrAKDI7QBqU8yoKRPNl/oC
XOuQaeBXbJKYhYZTZmYBWarav1chSkjtrMAb86t6LcnehAS2wSxSPtX/GZNcBLhc
9EfVp6QR7VDrNbN4BBtCMUxJVc6qlXisKEhMmEpEL4B2eQXNwzBhXIVu1vfA+5ST
CrhZ+Al+fAFRTmdv7mAT5YLeIT71RtkO5fw/eQxdYSQm5Km8ozL33lIvOObDryX3
wmYxuWxjDfr2ZQlYp3vRgyjDrS5XdywMTARewLGH4Q7S9w9j2mjQCdTqMpKJTrgd
gs2gXbkF+ObtbTMKhtUetUzgwQJvmuxnMoZ2SoXN1i/yLZVlN421MlV/O4dXbnxl
9nRQqVyWAxgXpzxAXhNWau2mByoFvEDsjsgzsmDh47yhHVKzLEwRtZuQnZUWgp6G
e91kXKU/OUP5OiGtSBb9XrelGkrIIuRiC1t+Xfz981OaaVi45YCM9uXbT7tVdigR
/5makZJwl9J08C0b0tMvseOkT0Q84jRez8flyJyJpwp5d2KJTan1+HYjGC3qhw4k
seIiJT1PNei9R9+a4eC4R84tbtwbeSQ+T17ieY2+D7VaQHNvO3q+nJ0x+5D7Enyq
mxLV9at0eEMyAROBFB2ezzyQI3BvJ07+M92KEMSjGk6ofe4Yx0aSIXjvwXyayrvH
KsVHxl/8sudqvxI5VQasxkPC5oSTEEIOeXzvHdP8Ch73uGrIVrRElvn+h2LQSJ0Y
IN1MnZ+TaQLPG4mZwE0eXMSCLgZoVvXGGg8Uz2/IpzMIPAaHV1EXAQjkDXnT80Nn
SUTo4M0htaDQXAZR+FtlR5y2T7Ett9xq7hkEi3mwoEzAOJ05zBaCGAwZjXpwsTjk
5bLWRwDiMe37TCFmcaiN/OWYXgh99u+aaYriMHXHnxZ+qD0fxR5SrP1FqS9oKzjY
xSom3XsMuhT7UG+Mm6tjF2ybnihBOPn/WC2Kbqltc0bo3N9nD5/U4awUc3EAbPRK
iP6DGkYQhKw2V79p1ceRWkQgKWcRq5IECUKwK51nQPgUIkDx+pglcnlChOqaWJqx
Dcl9QP1Pk8jZUrBbdgcHWx3wS/0ZdaIN3m87HedmfEtqmJ+YlWUn/ZLUAb/NHxOC
OboYWvcR2fFDWxiqHMED29HjrFT5Z9Zq7kvREvesNXtZfw8CHIb31nlmmQoMoNdy
odDd3X0hrAxoeCq7XM/XXMfBoGAKjoNOoZE0HiW+DryyIVD6tMI1PTCyWMjLFBXK
oEU/j0AeJiRUGAEUFNzhMD1OApMIxDQmpPsneb9FOnLkT+uvYKIn3aDFYLjJTEFX
Ge9zgOWWXy+5VCnEzYI0L1GK7SckeqFNhGXVIT+qDgMxeFnYBz9EhODD/UmyaS/6
R/R2Q3l0gJOAwjok8QXvtNF1Csrs4J9AeiI2hJYKC+zC4gkyP/fhnF8wfu9DTcNX
EXHzY5Kq+B1K883QsdZOYKFhpg9zdYwc3hoXHIL99cFyplFzR9mIrXpXlOaXm+9H
bfFC3BftXwY18HDE2Rh8kOnvDUVwuAeMe5nAWNIYAjLXJnA/BlJNKDLbTEAHhC2H
Lm0MiE96a4RDjZTq6t3D44OPPeD0Cz3FEsWjl+P6EISVScJW6//2//TTTfnviN8E
BJdSBFKPz2/JFvGxs4eVdWD1509zlIbrrxCZE+08Xr4/n5Pc/6vzfMBdYrhlfX71
kKgr5AxqZFZ8Xv+RlNVGnmTR69mR26zttEeKMeFGOB/1G/k1Gi/DxXS30343Spkh
hx5vAAt/exmkg8pasrKCq6/miYddOFCa9WK1W9aVXSjUwQWirXwcoCWgyS+fPnzn
XzmfLbnLs4ODRlBEvdipalodlg8AFL0XkspQ4p6qW8YsWQRZp1oEUjGSdxrDykX+
m98aG+tVVNqEULXLo/2HwCqKpgYPSu8TFFNaDm78b+cTbM7YVE4idBfOEP5k+eRP
SzdNBjydjo2Y27tylx22T0sbErnRiS0SDS4y1umHMfZRUaEvGnIi2Dp+NZkT++6j
cXqn+WuolopJZGTZNFK/+jaP5bJRDz2m4QHRTJ7Im+np5KAlgYzh35IMZ0nsgG57
N4Lb/9gAesjskdZKassl1acaBreM18aTLkQRUtfN1btUOq+EEBcH8a6V3kZaqDpR
u8xZn7fCoKtDZQPeqw9FUcjkNHVlqlAxQOGqiBB5R7amFGqGtm1oCcjIFiYe3gBA
g1j0BksLPy0j4qKiBMutKDgAkWpxo0sXTomojgLHXhFYIg1cdtff/L8CO+a2rMKH
/nhtMeKoHzeKbnfRUeA8/i53C8k112L78vwQbvgdUaD3WEXyffEvuTTmfP9VlCux
Y2FZddmJCKCtajS42zyT7ssJZ2rQIUlgRtoM+jhNicGEiiu+xewIGZVn5NoJJM2u
Mnl3ZLSQua87QrT9NPBr89eBQBYF/nbqyXEr9L43akrnS+JcsTxTnEuO7QwtVtxM
u0wCzaIR16cdwZTjqMPo93RMH25ZKEYlZxGJl1PL9iJYXypgV/uBL4W5WXeWpDAD
TE0gJ2I6Ww+1UupIuJHR/poR2sbEZODvbfmP+w7pHRC94bw8qxqE32KPw1oEBfeL
ARtzNHARMhJJnvpZFtAxuwn4LNkqEYIsf3ukJsd4G17+0pZBIjG80KrXzH30xvSy
KOn/5aRAC5X5wXeJbNGJt9rPjwr2F8bYpXkNPVZ6AsXswO8JI9JHJS8S7rmo/Ona
dJ/VpsM1Hl1rqB0Thb739C3bqBzUf8jwIj0pDaKmnkqbwBJaVgu4hRoV4jPohd8B
DUIDwEQiY9JotVU4KA4yQFECx4hu4o8TPqSMZxFvymUgZGud7tOHqhXGM7Ml7RXa
0/Zqd5Q0iuy+8umPRcY+Ew2AzXULftvuqJCdlOJN2D1xQ74CjhDC+Tg+mafZrLHv
Q3ijcwQn46pgCsRF8AsshY68DaNY+uvyKx4qkRz02VQUM1B9Vsa3LxJnQ/A0WSZm
5isjdvNOURVapC5ir9guT3F6ffiPqzRqSQurutgqbLS1E/w8MifMglGlDS/1EJU9
v5DwS6qvhhumb9EWkdi1XvY/QkRAcAL8STyIGC9g6iR9mxRJoxAial6BfBeQNUly
h5mXupAhAz8mS1Iux85IInd9v1fLZDOWQ3Gdpyj4vbTNq68Smh+XGqLqaTs8nvQl
CmtNZaw2LSy61Gu113HyWiiSPY+ZjsYhgM2wi7JSkT56UHEN6n5Mge4RA5as3Thi
22idRGWknU+1jqhSwiTCFdiGXCJENKNum4KaxXNs6Plkn+zj9uSIakkeIG22k6Ic
trKZQxK9IBZUAUO55db9Y9fcBOJYMH5Et25V1TVsg+KSzwf3cbse4cnA17CUSin4
erhgxA2HnWApRqH8yKerfWCrvQK1v5Yva6p7IpNZoIWC1a7ionbSp1wQi1VksVdT
eI1PCMffS2kJu5rUZIfqc0++bhX8cFGqD3EnXh1kzGQn+hgRqGkFxypOytxXRrjK
hvR34m3YU+NVHyZp8OiY/iQgsNSpQrKCCjKa/DxkYc1k05a3X2OWvUiauGGEvRf2
/gmWt06M1jE/UsgX+QGhjeJ3oRrSG2QO17FRk0i6DjVcjBp7TIboOu+QuNUe3mqI
yWOUR0SBwf320wziDXiWeeOnaO2uXKr5pYkYUlvsCMFqtTXRVprL4859K/wnwdT3
AsZFzPAX+bDOuwC72zb6onCD1mH9qWLm6R9pitEJtobDT+NvwJQLJdNiJdBnKJiy
BCYCkalZQPwJCbGLJuismIBUuoAHqMCa7dMlDn3FfWPG0EhdbDZnyNb5KkTmBtoN
zg9dfO3zMM7JxyhA3jjbLcIkNJlXpXQTAQOcRlYudgqohjC5fXJvYzbcHxCsmEAH
ZqAtWFuzES7IxBjbF6LVgUq0iXXD4Et8hdqMEcjAut6nZEwSbPpnpFuxg8+hGNgf
BWDCIubjr+HPeDTEqndH8AJyL0N5j48G3SSDsv1udjpYKnJtg8k51+LzKozD7U5S
IP4AXy0gLIiI0J5ZW6ZY3x/aXRgWOdfsW1YwMIIAb9eFL815BWuBGsve3EIEOc5W
Bi0U+F5nf8kxgCfZ2yCoEETc7+br4/MdD1q3BCg6DDxpSS/F2mCtyfy9E/ivSF6L
c7YFCNb4bGFKUznllJJHOVw3AZiuw9VkXCKERaYQzlatwi/qyZA4fifeFUQUQ6L6
7FdGGe24MT5HCeS26j5SG0O4cK6sgDNgnCNHBPtxc4ivbp2fpOG9QMHMgTWuuNzb
LHJiJTfOiGMKE3EaByg4RMiir9ghMvArZNNTJ6mVU3AbuZwuQ8viGY12qpHb/NVq
ZZfPYtVmvGoSk0/WuPcPWETzTMaHVKrcx2bVrDMg446BzZes5BcuodpcPyB+uKzg
uoMuc9t9J0tjhscO5duc5eVvESsyINy2DA7A8udpc3g3bU5VRZeee6Z4v5TzXgvK
SRGgff/R7mWIry0rQs07qFVovEpdVpTUUa/99zttRKl689P9FLWO2RuLJd0GwV1X
OnI26MWly+AbE9evnk/UH5XgeXcmmGdOyzW+bPSmPED/i7usrb411uFA6rwe36/G
tsbkJo7xm7OeNb3oqMKpqlvbWjguiFYVqr5oBb0wesXZzmKit4A9+FViZbIMOtCc
6Ln+A526ldhVy3+zDA9gmQnhgK3sOKelhjfBQi2PmX8Lk2wcwqwi4/MSAEWFy9Uz
UmMJ9lX/FCxR540aIlCYUIa/a67/ZeeF73UtpUk/tzbyVgpT7gz1LcWRdo1NmSSN
7cv+5u2iDBtQ959hHMXnY/pRl3wpavzJaTXbITq8pw16Y7OJ+8yukA8BEGdtUD0x
bGjpalVFPb3dwvdv5HMquPe1aniIoPKH0MucobXweavpk+7+SFRCvMZLIKECS6pL
LLQsKLSUJBM1xeK+OL7ZvrV7E+U0bkljhf5QmhvwegRo7yFvVMHtnnvnxYX1wDLs
vqMe/5+D0hZtmZpRM4KNCGbJjzGHE+QjvhWURFNmYHLChQWirGKjki8CxP1EBuSw
h2aq1+uaRSMgkkGcaTjHkQ2rHFCB1BFRPOsCkXgiKed1WdllGn8dnt2Mu3TM5pxN
sOHxEwocLdRvwr705Hv69YJWmCUG9AQ/eP1EudUxagrPRoDzLb5bm7RVBhZtZuYS
Ou+V2M/WF7ZgfjTeyO/M1WUmbTLqAQpKH3aL+88cZRS8O4+Wmg0QKH9YoP7qnbZh
l2IpKBbLs7zLxXmb3o6BTKFfvLqO9n/A/Mjfzxv9azxqLMFrFdkI2cto9ZXHnvbv
RWY1mQkbXDtGJdHG30Ij9MfY0tc1OB2X28PDJzSSCoaMaa5nPMp/9AXb0N8EtKz0
gvuyVWNKgvgqRThkxQZANZnxB1eqQIDs9OsodKWshmYxz3/JxpnHVBNf4R2qu51d
Q0AQCW2upmlmPTTt2pOufjxoVm1+pEVY7PGbn6c6sXUJdEPNYAJinNuUtjB0Q6nk
1OzIU6ojV6IRMIRcHuJk4Uw8sRgmzIrbQ7to80+QCuoK9VPcPI0ij0EcLt7Uc5Vs
4Hbzdv52o2AXaw5aow+ZXM/v77VDTx7wdZjCCZq961kw035FBFwFs0AHdNfguAon
AXXzM8N5xXZ8PR+a+JQquY1xzpHvZ4YJJnlQ/3FYg8NP45VT76B7xtBCDwJzeb1U
zTUXtWNmDxsFEnygIFuKh0fjELb0B/LMxRxzosS8NgIxvy0JnC2V02AmEvQGMF2z
P+oQktLBKKuoW6l/hA3oPJpdZBFyzstjJG7bVPb2U63v3Hb4MQQxlFGUdHmwNh4R
Yi7ClOehI6SPsi9Hg+fjTaL01YOudK3esmH7wpgoY7ZSRemv0d8nrOv0CLbym2aq
orBeAe3V1z3BQ20dabJSi/73esMxmkcUfv0467/7gCP0qNgadNDs7ULutMXWj+KM
L4KK9mMVmZe8Jnjbu6rCr9hchgGj+ZfyML9AWNcz51OhYiibjK1JBkX21i1oBB0m
frz10d7LsNI713bfwbBNSyfjfa3DLsYD8YoUyi2Z+5BtHGelbd1I6NtzY++7K0D2
jpNWO5Wi80equmC2JxQSTGey4OmIHuCb9idoCsi0lZ4KLgl2EJde9oQEVGwrJqyS
4IeimmBENAMx6jlvK5/VhtB0VOMVfRZNJ8ULuzckyAJ5buXFS9Or+7vI23VhzTnK
PfXgObHHdVdWqH3VMs7OOzdDhFyeec7Y05BrOT9olNYj9zd5qmNfhoL+kplwo/jD
kTZKXN7RfLmb+pA4mbMZNZQSgxwp5TwU7z710KBRIgwpdstck8UU5kO1UKvXx0Xm
bE28DWuWbt2LzTCqS1Jg6K+9Jckzqzjn1Rvt3+kEtbOKqZLS0U1BpVFK9xV4B0CW
TbbVYbrNTqMD6Dq9UPna4FRjMHaBRpy3Hu5M6iu5klGmnKhe6gCxEGHmu0NW8xbK
Y6ixfJHcPEKep+chGlew9pKs2WtLAnY3VH8T4kqeYGHv5lvicpM8QTCygxumhbeW
DwL90uoBvDzUN1tjYsJOK7Nt8s7ldCNV5Jei9bid5FuCuqz0ohfPVDikNNbNqmfA
vtzWY0vAZcsd30Z1XVVBwKZxNg4KViQaO9lyfpgqfLv63rTCt7PA4JYbYY0BioHO
TDLW913hqtGljTeSS3YWyRpDssDkTDiOCmIFY64GS3c+ELebOyJtfgnbJg57RJQ6
qrhDLBY7vuy839qeDuQCjoCmM5hHpvHvvu9+gpHbr/JTBJEIDmp8Ym9rjHArNcWU
R3ah0dB5m3rGvPWWZsJVOHHn/7ESQrxKLBu+n2o8euKzy1RO4iaaksDqax0j16JD
ylIgtROl7ChnDSuZhrPGMODnq0osfaQ3bSDJ4xAOunpZeWqdyQjKIqCV/c5wvy1+
u7UtmOY9rOtEgQV4YcZxc8ORbzG7hLhFjA9e7ORyzaj/w9xRzcsNZyIPNFsUrcDd
clUZfi7lU9z0CPdhGZ9kea3bQt/EzjVRgqqekY/7gPxzcdFNUtdTUYTBHe0RmutI
mn6eJ06QUDt0axvO0HVSaIBAzSSigl2EiT1bHzosyj4Veme1GX5l/+IVrY7wbDoh
9WjaYSXTg056JODY6z1KIX/UYnVRd4f7mDVc9rD8Clbu8RSf2Ss79lZROfXuqb40
nF+HKnasS2UD4J9cAmvWIjl8X5pG5tJOPbf2hu1w00AQtnhoxgWZd71dDPIz9PDP
N0OMid43f0wACyTYCJ93NJ7ymS/JizEFyJTXXDZjdH4AmuO0NQYjNaJ17gwB7JMB
2EAyq8HJhwT7W1/utlJ6SPy6uzcsiwzTUgg+GPjC8rZaPosD9RT0gfRxYVYcBuaE
670xpWlC1hMIa3v9vkYZDlqc4L79MqVD1JskqMsrdo/nPdJAhRMAueDyKxYk3tbi
acgHKfZ8dGfWLlK0AYKiX1ptQHz5w71+7Akkec8AJTitsBr88bcFqcMG78rmzWG6
dFq9EJeLKk9sZTafVzBuzLAT3Zqx4bgHbqylx7nHUTaWPVRbiHZkRiYWlpyc/l3C
/dEqdrTjArJ/f0Lf4wwJGcAAAdmfu449qHt+WhgDvltiBzGkKyN9n7gR9m611tCX
2MGW54ewTiCq8fZ/DZfJAoiLloaHiyGwGL1CgNTE9k9/NANWy+C3ef8oEWPHsjhg
OvI0bsbiUNk3WbAHXeJJIEJEdVr6oGaAhr9T9wsThu4er27GvWqvxdqBxziQOry7
7vQ1Nh0tMijlgRK4Lnwtr7EeMxfuVjHA75JWaBDDd8S79X/xmmB9TqqrE4vq16fF
Z0TXrzDUGJfQ0+l/uEGo6AOwDYQC97ydnFqWNBa0dJDDUOxBnJ9XeQjOS54Yvqrc
KKZkVRjQcEGCtann/QfQA4C/TlT8m5H7UeeuPyKz0xdwyaNtKr23sY1ENLOThLAG
u2pX/vmeP+03c34w4cMfl4sI+MxhxL5T9xSIt9n5tHfgew2/4GbIgkOwV2XcM32K
kEx77KGo7apFeqlsipclYpUrfjfzA/g+QwbXlZrKtWCsg3OoHuKR1ksx8XdZyL8n
CHVTszmZ5706N+BjTcw2AFrWDaVBCV1NCMx4/1x23BR+maqD9fCAUzRVUrw3hWfF
/GGNuYTvxgzZZJ/SGs9FJ9uvAG06MKsnpHjAw4V+DK2RAUfCWmKtCrSxAe/X3gq+
DxZ8IH1FjnmHH8ZKb+JOT+7J5+Cw2vguvL4KWPQDgsWalhQis0N98etw6BaMhVX8
5aRaA0SqD7i8Uc4Jf59YhTeD3fuDDx30+9XDbXsKU05GL5BCIqr6AzARkNjFHkD9
SYcj2YX5pTvkq3uzywki5W235PH1ks4H6lDPS0Kp7a1/ITOvPIqbdX6ww2hQ0aph
ClnLyTCG39ccz0JHCJgD89TGdwunLsOQwrJLTbveR3UOp9LF0+rMw4IB3awJtY6K
rS912QAalOXhPSi4IIU3vroqo2lCdsXYb+inZqv2n6p4FHnwVQfSaJrE4u/OOxRl
JFOZGR/hvk9E3/S1fRpMVjhg7IOhNFzTnfqTzC7P26Jx1f8rEtwjY9lHpepQSeNd
1imXwQyY4nB8vuslNBbt062dPMdbmqwahQr+bNEFw3lTvFCSh6QcZ81kgXR8+CKe
GU0/ux4IUsKS47aqNgcauuV7rY9eZUGQ+AmM63JAcFXvUfAoMn5Pwn+rmd6IMJck
pRL35722qqO4fMUPenTZO1cIxVt2QBgjdZearfj0QESLn71O4pSd2qvm2GAoWKlw
bAlYwU9O7WO4CMMPsSpZlvQvqCM2rxnsHtdZg76+cSLPXWrRyWO3IfmsG2YZ0PHR
hM6Ilvs1HkMVb1pUp3JRlqZYaTUYhNhao8tbAcmIKC9m5lC6qFwq67bygzveYjuj
9MfLCla6XamLCaaaUI1Jk7ZKFu50gGoKZVA035Okhr6aG08QaiH1Nx7gVs1rxzm+
n7erbz+ylFBXpHu8lCOZZ6X4u4VnDaLClCMBweec1BJXqrT5sDI/gGdoBDl72ofF
qGNtwcCFAprJ7uaPmaDwqeuKzv+iTGrA+ZdaRoJBEBogMYOPYM2FXN1YDOsTt6Zm
zR2KffUlpAUbEQKXHLkSiKI1xAlAY/ip4AsFSV3rAldhgVTkZh037dMq7A92ZehM
Lp24luLFu/R2nSByaublfymttgJXpVK+eYoygCCcSpbLhVuY8HD3goPribrQH7MI
q+j/gBACPe/3RVA7YNEHR8LrBqSbdRwWFNW63QxmC2gRa1/08zNTEGZ8H5OAOxJk
A4JbkaDRBc8hI96Wis9AGBEEMFKFs7c7hKzNgNrd/n1w3qGfY+YZ/85yIOCsrprf
0KxSa2AMmjPXInLShs0Fnzr/eEDiyaIE5FxwpvxzP2wuRMgspkAhlspGpq4YFL8p
SYE8pLB1/Kb4rSfbiiV8yWXdgxoE1OvaZGoIC+j7oYUbS1rMzDQhvMSVZtyxHFTh
J+o/LmaifKAXG+FhkP6jY1obyAwHwjloRz1GjB67U3/Wzk2sXBIlsfaj/EFvleqd
yPMRHwxGb6NJj3L+fnQHGYguofG7+TYla3qbAhQlwZImVc6GTu6KWMo1fRbwkQUh
fghouNfD0UX+ZqOUpV9BX2NdYxXPrlmhoFjZwl+mZT57cjLyRYDZXFbXfz7364ik
KoTjSaycEyQzEOQdkLI/cYmFH1MV0z+cxDUSwgrUbfaUQCRwwjHhYuBf0rLgFNnD
ht8Y1tLF2Pw+1GSe5CVUP+XZxGFYjWCtpDyLFXog1STPl0tr2AdmU25w8yltAdvD
qoDXfhWYop1hZRQqsDF2oGgiO7GYiZiWKMAN4fZSqAxiIF2M3422bF9LyTGsXoaD
19E00Tlph6NLL6a9Fq5DJFF3xVqta8Pk1n9UsycsOhDIuh9ewaR/2DmZFjngi5hs
0+vKaipGUGbxgnU/iV1YfshA9VnNiv7vLB7xZaigaQnODafnGDHIsCy0xkBFWfsO
wCNUbOoEMjIj1KlpeuYMPlAgZS0tadmIMtUGM2G5Ojgvg1A5rZajeQS2epmCHfkQ
YQoRXMyi3m1jS8oXAG9M4RQ2jje7OT4OF/rGllC32ojO13FDX2UgYb4yzIN2Czwg
MKnLatbE/m2jCMOddu2EF21PSz9M8FaXc3ZRDY1NCcmk1PKS3l5BRfNMM2vKXvR0
tkRiToYL+IUkMXF67cs2/wag0W1Qh9OxpyJPqetOs9vhRH8CVmhBFfweg2UTydHE
M/Gn7S48XG4PBORKE6n3BMj1YT8a9kFNE/IV2t2qlff1IkjJlUq/yt8z/0TeZWWX
PQspPgVrsWJZMNCvXq15l1JzSOaxij5bvJkeq2pez30iOoko2IB14W+R3dZJ51jT
2wd3iej9+/vOULYRUPZvtVFN18vRmpnLXzqS03rD5nYsLl5OhwKKu2/YYWVecBTa
2X3yw+udJvWNldpcUmKCgblMUW2FHJ9REAre6Z75YB71C4/nO7rt776jw6Rnj12g
xhZ8gHp5WeykJOfEWBgCAZIFctbp3op/28mdM39nznts6UdcfTIo+4MAX0l+bcNU
xU2ESKswjBMOkknIOaGhIvIE6O2cPbbmlsNRazotCCpmo7uHkQHL0Q6cvpUEtbkc
CuArH5rRxXfDZDqvULaNsTqevBC2c85KFIDW9fOmztH9T5mIt+U7amOZU4s9pj0T
CQvQNH98RpRLouX+J6Eaa6lQao+U+GmjJnxs0rtGHL7usHSaReJ1stYgEV0HMc7N
JASr9ICV3emV4CLa5FVx8FPAVFp6JU2slF8UtavViMGXd4SetsRUyQrF4gac8S+7
0fdJixaRIrLmF0RaGRUyHYg8ZZkFsVIbYpWWcHQi3Ty8Vp7R59Z/qMQRWrQPJj19
tix4icTpsPqZHmmpG50lqb8uqWv/O3i2+G3pAh2PbO6uW6u99ezaoWM6zQ6F9Sdv
TDbqsv7OxZ0x/TIbvCOjffZI1s+6+jTanu7oQRxb0rr5fRDM0gN1v7s/gFZ1YaiG
SN1BC4FqZ7NLpyOsXZO/s7/vkdQA4fK3371q/fynPtHrK+QnqJLo1JRAvmoPygcU
3v9P5ocOvwnDquDp0E0H6aqr7Y9w2L1A7XvSIRTDCOLGTxpgJObUqXLelwSJPRId
lfZSBOc6b/t8gn+Wivtj4Xm08mVeD1jnlc58+e/4hwDdIWOK5OFv+PdIVHCL9nh2
AEUKUA22Iuxdz4gr3r+Ssj4lPCa/DfGUOIMk4C2JL1QkQ7EGQOqKmOOxS5FM3CPs
9ijO43lMXl64kb354aXvnBBE+lMVAO3aFculneFZYidFdfx2gzkEVgfmZOg2nisv
BdpeAPDlmo9z9370ZY0fOuzjR66wWrR4aSQNL3+I4EBSdV8INoqM/m9I1cKR2p4U
dv8I1JvjfjmrjWU5Xp21UK7oueCQ2UE5LXepYDEj+X0CvtjmWlIuE/Jb+MJeTO9j
7A/1jMSXrwzARZw2wYz4r1YmCq/cYYcJhconzWNOyMLWr4EEL8HyM7PP9IV/d0ow
JyRdHZa6r6ga+MeEDqtK5JbmNcHnl4KWUBbUQ3jrfEGkzXKT6MvAy+YoXPjrVeez
o/XRlAjwAapXFhK11FuHlYaEdh40DNo3I1WdSO3VanDbKBjqMNXrLTtNwL7u219T
5o5+dr9RqfYfZc7L+5lK78YTPU/q0WTpMuVTxYKKPoC8mOfzFwa0J62BLr1JGpB9
po3P46N1xrIC7cXQ6OCAt5fhusJKOCgJfEywRKrQ6JvouKH403lsaIebREPcgSfN
bDRtJ2Uohnb69CkyLgbGWAIy4Wdv42HhwXP63X6SzpleN8eFhwuEKwIDtUihV8CO
W0K0pqNaCzv8uBMUZlVi5W94kKI8LG22w13s5CbMsGu2K3+7g6qORyxclL5VQBDV
hVjAxWhyOxHpxeET3posOzNhgiV2yU77s7W56msLP7xHWdYTbjRquHjbsXMpv0Mx
ThGY5eOkrOLJ905E4Vn0O+KK9Q6lAmi5/8Q6UpLLyzd55Fk7ohohhtZe44UtSeFr
ImyR1iCZ8tX1f9ylM6wquAzxcrcMhaGdhZgAqfHCrCD40ZonpY+Xltgu8obVSNgm
k5a2H1dhBA7j9/Fye3m0JcqCjBwUxEZJI4YF576ysXm6HopKwjhrlwioAwWN+eY6
BWHTqCl92tZVRaUgkZtLEDe+8MxD+esvMsL0YXa0LhqR6qVBBb3syDr5GUEpgeDW
/v/y417Lq2NgWA7NRZ6dE9KbXYatwkmlR35+EBB5HYLXhfvNpTAxYIwF2uFdx5Iw
KRYUd74JghgkTZLMFkk6MB6cqcM0tQWq0ydLnpw3ZaXcGaN3R2A9x5loQrfQG1Kn
B2MLNP2kuTNMX/UtPIb8NAls2teqPZvLzm+7a4hioXhjH3iGMDvyzNed3Zz0dKsF
YmxyW5XgjMymeNjgJdEGZ815WSury3X36o7F74YCG9hZl8uVUQSkTkJMLEoCH4mP
ghqhkAPZbmzlC9mS3deBFcP7/dHs+Mmu9tT8/WVF0DHesutDmG1c87PK+WdVRX9E
YBn8FhMp7NW8J40ITu0q3ZeidOPaxZXJfkmUAI0uU5tKsrue5dr9RFrOtKLn5kJv
B0ESC2Xe8haN3XkdEapQ55azlIauoCTLD0M+/idCAaLIflWlsS7J2y91XPkNjaXx
wwR+18FmwZ8XPhwKisleDbRVG7T4BnzdTNjXpswoxj0TsNYBVZA866owhRYuppVQ
o/lLoKnLKUKypkrpaKuR8LBCnPFmWrPn24TOP7RM7zz0XT39FpM3FuUblgeAiWSp
FOdUwf/AS9JkGq9e6UIMT5P6ppCtascjOVj6Nt7WwgmW5wWELjxjf4EUbs5zzyjw
lU443066mfG9/WG6wPN1LMvXYdgiMB0IcnX3J4Iku+Jwhn1buLxAxyzqp3NggHpp
46M9QFmhnM/+YlbLiGciO1sZfR2OMLltq0IJOBkb1eVx8/ZkrXK9n8mbIe0v2gH8
8YRH3Fmm6qTASpCkktxY+wuMnAyZmLDU0qf4j7CLsy1lniJ+cGLoMQcsrCWo47Dr
ApCnXnfYtWujTBZDE3XKDPI5rh3g0/VHkE9NAs3WhkDAmnqifQsCINTmzDA55Y8L
f5tqNKYsGkw9GuKfTVFlP2cZ6MWisyGn4zQIn0S50Cgdt7ouPNeB7e/cIqGnAGjd
5tz6XG7g2zeaigxlSXZI1t/ok3rXe+rtoRsRIEvTmXStQW6xlBsEPz48cq0YQ3Ka
scQU7hSwfx1n1BPpA7pt3vTJvsA02qjK+nb3AuwqTYkDgo9gO5YSpyeCiEJ+CfRc
UoPe6WrLrrkeSFTkF02tz8xESEX+nYliMg3yygPtln7juJnQ2Ykzk4pgTzznIb5a
zfkPLX8+Q05J/esYsh9BNRW8fuLfecv+Dqixt6fV16CQaA+gab5f/mNYYP0W9xd1
OculEPXlIvdCpQozydT0ghv1d0Hv45LypEBbZK7kQc0RQ/wk6Q6De+tHbuA1C139
iam0DCkTGd2J7yVqPv9A61pPrn2aiWQf5OkFkUl2fAWOBJPt6tB6hxFdxwBnWd3h
mO0asGNFb8gdDI/VgFNYZTVLM+PIaZT7nIR5z5UZYi5hdzUSEsTm4+RtWJKMxkzt
OGAf5l46eigljO78oGzt18DE5UmAV7KMPk+bKTP1tFmcv7KpMYshHbmvopmbKh7f
BVd6Pt5Lf6ekIThPUZFToKQ2CSIodT9qaG7e2dnDzG01NbT7qu3g9m5ZQdANYqNd
BJnGVifU/ppHU854NG4360SYNTM+LxJ5jWZiR0IFIT7P5xk3V5+aWHgx2EGm+Wty
aGuPr4eXVN5pv/9Zfr58qXHhJwBJlnfqo0IJOwUj/j3ixYfehoW37u0l61JFHCsJ
AjszuyPBlGEeajt7KmR777Bn2dowaLFNSACl6tAkjV4Y/BS8AmRs3MDhdpFbrwcW
xZEh6I6YUzTBa7x33eEd2yeKyX1/NZBrDx5prM2RsTCrIaZICddSZc/0dJUnDHy3
hMJvPZw3oNIBGVSyMl8xB7yXumVHFrgrDls4Wsb8bWAcUT9W0FQggzoVDK7RV9No
QYDswUM8Ze2+H6t7fv9eLUQEBdYeYejjRNQUcdSV9ObdpcBigwWnV+lVebnLHpYU
QqV8u2Lv3/ym84lNWpiKsKcAFJK2xGgCvPLOXFgX4NYk8lkXRsFVASxWt1Klg6GS
/WKBZ14nqeDS6/siFO7eoQFlkY40T6QUABm7acVR9G1xmC7rMqN+7wbL4Ti74iO5
lMC9ttHa/RTenD9PwzmM1UGicZ/WyNXuKoFHki30wP49GkbvV0Rqx8ak1A9NbejY
hcXFlKxwcrLRm5tPY9sYLP0bSKSj/WuEFjm7QlQeVMNLBfSk6IImYP8UzW8NidiN
yz+Ke3tWpHgUoxE17Tbo65kfUdvoYOOdwqAAzC2oQqo5qF7KbDy+IZ4UTWPG/7b+
uJTa6lk5WqnqNkozvTHCoGUEnR3woKyay2bGErJK+9aRg7AXE0BIvDbf56HJdEnL
Ie3p5GJX9uZM2rSw3GOC1DZXn9mqxmMYHWZ3rznbD2l5vZ1gE8EGxWVA2Kc1bQki
YyA4ovKj3lz8OklhXFuRgWoNv+VYq+HegLBe9ZG6tyKyQxeaTh1PNtssL7/QgAeH
8FzMzReY2+k2XyZeTxNqYiseD/GJ+VMt9bmiKHpG2t+DB+Pn+RbiXFCt2BRhf292
HQJdP2Gj2cwqXGDFQytBt1TdZppI0A2X/70McgltSm/N/Lwqu6VQUKq4qNgKF9CD
jVuva7zJFo5up9bWZbDmd6pIIqvFW9GajwBPIKo4QU3UDE4YlCSXDmMNp6vnXg2F
wSF76JFFpCqX4dVxunTGnLAaf4dtBQWM0s9rIpJ13/pFRQUw19AC/Ro7YLfSRSg9
ypMn06smUGDLPKaAk7WQhNMU8E6k3+xGRpFIbuBx23Q9pvKkJ9bnwh7IGqRNra4J
VP4Tf56fqqD8Imkvxf0+bo9KYiWYDqJPq/h/2NUwICFK/2HB/+LANCvYSoPdkJCu
HXEfXgepkI/kyzp8+7mddzdAk+FXGRhjMdvGbvIZZHausbD0JdVBBYTknU+HAhxY
yu4J0sfxVTMTbsp3RX8IV8tJWP1qiwuHYIRFTy96GpN9uvXjrv8TjGibU+FF4UG+
Vuh8lCmPB+f6rfpymW6rsmGiijBFfIp2HDRT6QwsAmTQ7xQrrzSNrHDn5LVb5qVv
fBm0ifjyjyPX4EmEXJZmFbfdHpLDAwDf50Ym22OprFg327ARTg4M1GFX0Oi6moF9
0tKiCozU5quWYORhd6trz/btFYqH6i2Iq+iGjIVGPhcdX3rcZ4FKZ/dI8mGmRwy8
iIiyRvrhWh1wHiRQkhQ6NOUul40zyZAiEbXGrXKfIrDmecHfVHdBLC8Odof8GkCb
zlOBhZGG0NsYufEMZ2JAzxNUTEIJFNnlfZuwlTIQNROBQToVX1wWNTt82z+Jmzv6
cy/NLQHbonRxPYL2d2d5CnuMZwuGqyd7lVs7oLuoYQFuayzlY8EUovArqBhx/HUf
iqfoikiZCExwzXkEQ6/KnDmHVfL3aEXWCfBA1fSWth6GG5rl1YXEm+i6554PVteT
CIcS5lKzugjVaRDZfC6gSJZwQH5LlFpek9iwEmjB+QvLIRxM2946dk6ozddvhXOz
7+57v6s2nCB+N3nfQupXKgoh8TOmWan8qMQ7d+qNTIomRuC4qA2If/Jqe4H/+yer
SkshqAzBC8LTJ3I+U9Rt6HPdLIQnLJiWCO7V/QW9/3DfD+ehXrpG2qtOVbw7yWVf
/3v6TPaEV2y9LXIjigxkNiBkb0Ik8trqDdJhid7oRBwbQesM5HSxafhoKytDwRwr
UHvlM08xfuE5kYpiAlqh2L2BTXwTu2jSl5XbEuiWOpDyhE9GzAkzNfP+Y0lT39cp
wUhtrPaI038A7RMAsb5IWxTbqOOJfrXiQ74KyysbXPWVoUMawCl7+yto4d7sR9dd
ZMczNAexZMAGKRee1EGisPzxeubIhvLmSop11BhVBclZbX/ksBZwaaSMo9TKE3Ca
2imtvhc8ooHAjhCXmTOnlNnq1gGW5igs74urq6eHPoNBKO7GYOBmGQypGRsvlXzS
6UpmlmIFnDpbnLMsS+b/THa0Er+H7oEQoRKVsTFETWauouRqyEpFpN1fHKz0nOS/
jnkn0598swnxhiQmoq5/bWt0RQbBRpg9vXm5/8YhOsLFmJ8Ha18ArrWEEnFODr06
41N8ejjQcIcjmuwpUKkUIkbzv1o5dlsCl2atS4R1OAF99WU0Z1Tc75ftA57J14vX
jO9QiItQgkf7e6x0O5jPm4GYGmYoXjxPWKrAmRKhrsRytmcpWqyk5NpeO0OiDLUk
JCSETJXB0vU1umN0WoiJH43lSWSsTxsXJtrbu1yvIwqKcZJIJeYMgeBsF7u/kmKQ
io4ZF7v5wgA0hhO6z5SbT6UZK8ARRsaVJ2hMEavysH0hA5jjNUdC7aZnXZpd5pvU
0268Y7nZPzmX3ic6QDKKq2amFzOnJ54E0zGggY+2ru8=
`protect END_PROTECTED
