`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gtN55eM3eOwXGYG0qU8qyx9iCBf+ziasNjD67GpCgxYYfZ0AE4DzRN4qBSgGHe1r
pAohhXppXPIGsQbb6iFG5FMEKNW9V4RzA6TNO32x8WM9mRlUshkzRwvhlNNCuZAl
z5pnaLIIT/cadp060mGmmuRkY7jz4NJdWs+vWwqkeUCV0jihz+Y0oS294HieEEe9
fiQug/BcfiEI3ZxxoM8eV1XGttuyFEris+l5hSNvY/YeG6uRo5i7g7Qu9enOE1DE
jRxey97OT9C+NHqbJARkAxCheDoo00gPSdTmQTO8ufZUwXKIJdr5ocOccNT+97lS
daKgsXcrVIJQQeQ9GSsvE5ESqFAeNMWDP6WEAXWi0eCJdF84KUML0+V1XxMwZRTA
WbfRsOeoq+1sicAWMuie96DKU7xgIDnN52PO1CoHGKSThpQRnWNIyZhFOh8auq5E
w1kCGGbMlyRPEw8LeaX7ov+QXV910WpWAeNw1HIyFoKVEJbMYg+rvvCu2/IeBo1S
G5RWFRVvWLQtu+cB4Jj8bHMH9OE9IuF7HLXeqf2ZUqpJGcJ6H9Wz7NCCndFMlD5D
xSK6YzveT4bbOHvksKomrIRlHPWMh7boR9RIFyg2AtPQs/2HTTUlfx4g91DljOfu
BaNrAwHmV+H3sULEZrSoNRzeZw0I9zXaEkZC3JFepSq52VBe9KPQ4FIZvO6nWwhD
`protect END_PROTECTED
