`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lu8xL/vFTFNgaAeLuUwefvz493S+7cAYgCqNconwOf6syg0Ei23CT0WDPKTN8kVN
h/8tciY10Lvuco85aJTTtCLFo8/g08wdF8XH65F77JvbXyPDoNlEl9d7P0rRkd5B
l/IPWadsae6ilD/sJP82OED6c2BTh4NFg5ajSX82E3RNrHWWzfiTaIgv0kbYSE/j
VxuWHDaomIHlzPNVrYsGD+XWtOHpc3BtlIK7vMtAxHjgsitTJEIJyxyBPopfuyvh
MYExJaexdZroRwJgrtdVopBatLPZNOkzj38FIcV4EcyHyAx08cS88f6wrnBSKt+q
VF69IQFQ1v54f7X1+QfnlDbqBi/3sZmM1oACU+rcREee2tX4gTcjQT1Uom0Q+Zvx
xYaxDPS8KiSoH2oLNxrFaaTLD2faet0xvjGOzDb5kE2IYoGthcaRdWZnX/PI/7mo
nB0ReyK76JYg5l+JSVtemDma1d0xg9cPKA7irfvjVg1dhYGWdcshO/VSq9wdsDrA
7OzPIZgiYRtUR/O66CLAhfPpeJvRUR1EZR/Li7CJwz5yOmvkG489Zjt0Xeu8P1p4
kUregjFR3LxK8YuaKDLAhdnGFZdq0QITX6QxNL2l9Q9rfwAIcoyjuobhpJWEaw8X
zO+hi/YzhUN4EElhbWPKDqq0lOzM1JhyDRBLgeBJJARXbN2pjQxJoTK0Unw5DAqu
3FpF1PqesNgudxP/L+u7jI/ZGotTF5Ka7DFQxjU9VcJ7Hzpd7LSy/73yctS99e5R
Uuph8PJ5Sknl/fbUQMRjDjisA5jXssXMbVw+Qq6S4xTytKIxY3amAXF7rNRPOa2a
RkeilNJHEBluekseNKJXlFU83HbMQ+jtIms3GykoBGhGsbk6IBdbJ53j8O82aUM+
/lBVakXNn82GYdDO/JzKxz6esqZ7CatWmWqyOyBRFcPhxPvxtpuWyXchXikTB1F1
5YmRa/+Adh66PUyNqpIGw/hNx+16ZX/FpBWF9iZq2MgpVMpKtt9RECIBO+HEAbbJ
lOU5mnZVLOUDoJlavjwZiqFpVZu7A9vBMxswxB49/A6zE2pnE+/dnIpJ0WRtxksI
BXD9bPwqNoc+kZ2JBE77klvHhnp5BLSlccFxDmKrk9m/JHvd7EyNr6i4L6yBiMHZ
mle3N9dJwjTuF0noEO1xOny8sbEFrLaUYFaAb5lehNlbgMY8zvBJc+vzI/DYqlje
DjtvRCaz4cR25d+b81AD22tUlnqmkivuwgS0wMn3S0H4LnYV4fiDDIf7HCtpsfyi
IR0B2Z0ddJspu03Sr+I3jdD51smzJdsbFTBBVdyxWYWyxAcqvzQYhLRF9mQWGK5J
yhWzBLCUfeOaUzTQykgqrisPcBt+7caaCa7BOf+XzQgYCRhOC8QPeQCfME/VJHAA
3JaLu2kbDJPgS7to0oaWJq6TKOBmZ9Wuc+1WNqvI3lc0Ey0j1kpzgAXy6rH5rXwF
/OVpMwXpaBOKE649QwZXeQdhGFXIoSymZrYDHrt+swbh+dZeKIRfzwBFZ+AS70gW
ENcbuzag71gjtk/0kmCHsX0Thm5+vOnQ1NuFaSn/NS427mOcptrs7llCJgZDjR5u
eq1hVHTE4lca/Tle+nyQd6oTzul9CexqdjzelA0IEn+9VCSx9lximktm5v+eDyxM
28wazP3fbOABaPBJ3ZVNp2nPm7sVcpA7iglNmlNx/aO6RRf8V09GAW0vV7YqdpTK
c829L7z6qaXWJhJcLbtvBb1TFB2CR9sbNbCiandFHA9dACce6YTgMIdlReZqyGYy
rX0pIoomCjwaL97NKh75IUi8iBAKjFsrUn4lppxks0WrrO0xJQyUtkOL7ZVtma3i
OlzbwqhK5fekwXnUVlP/z5v0nNXDd+nqSWPGw79u1EFbq13LG9bSUrrsqzBNdyxm
/OPXmXtnwDDuma5UkCCKG4kPO3qBtMC3QXrHi0KZJSXxpAdLHokqKLreUHNoZc0P
8MsTYHpkjrNx+w3fbaF4dqwyKz+03e9nTEJ2NyqBQd8FYKVfLqRcAcJJgg1FY9wC
z+d/v90RUpe9RRAtj4pA155LsLqsX9TzMLoWNrSaJaKGgePP6jA6PqpjiKZVIpuG
5rLoYvraD4gcKM62uc4q7JvRkWlgHumpDv7PMn/YVIszIxolZOLkVqD+SxPZG38E
+/BvBq75HBa1Qjmz0vv/+0jDAeSzpH4ErQ1MtYjeAbhe3v+1WQ3ktkIoSJGU0IPa
jYWyRx6Fs+8aYFsrW+IrcjzwSS5B5Uw6DKW+mmiOsjm02/8eI3Jr97FBIV5ATGgJ
qpsCbKlL1gPzjHTwv2B5uByhfliPdcd1uXamXPawYRSPURWvJtCbQNkqludGrUTp
fFw1fKva0pFsE23SYFW/3e9q2YmJ1VuOKi9TwrW0S0FKb+Gk5sUNlAmKc4EDCWAE
GBa226AZ5yrcfkDelbp44wM/ux56wMvO3z4Rdt2g1lThFO8hlIY5lRT9DDpNi3vx
oCp+5jdxgIDZBY2DucdOp1TBkRzW8qhRwKuYV6r/qC4a8hHgIuU0Kqr8li6xD8Ox
+oPzvnIqB/71PKv19lJUt22HFCIHd5GSdg8WGD48aYefjBzNEpUHIzopkIMTI8M5
bV/GlWWUtOi0yWhtGitUbhdai66N2bTcC69Rjfl71aCitmVJ50oGyA5x0Moi6qn5
Z0mfR693i4198g2ZpSYv3SQR9zwhqaZ64iBRXEuxJKrz+ztN9szWhyUIYKYwZVTO
oRUAHc2g/AZLItffFzVKrfqvYIeT+XxIasiasEy/rrs0369iygDNRVWxcnbY3wa8
cgUbEj4lASgsYSo4k9kTVlm9KGoBgYFezN2WfGFjfhoTVb447v8J3M2bYguX593Z
NHZBP7/nSGIfY1ssg7QdautSbQi+uwB0381gOvZJNagQtZ1d3MK3tqwvZM3YHbPA
1TRLMq6mJF080ij742JPLoAmdWdFfxFh8fbJMBMiEp4lDRg82O9NcNOIl+s/5IGx
P1OePogKxYrJn7U8tTrlQ0k5U56r9dHF71ouTZGHLiV7GrhGWpv1wqvlQEYg1yd0
UGA05jF49210kRgPUV03wTAUl8XG5tYDoELYz8g0Xav4yJygqRdXoU5eCIpDhbfA
mQIQteV2Zao16ctAQAkkjx8baUJxxeyfq6gvRpVoJ8Bv/amdepbDAgec8qfCvuBb
1rjTVM2TdqLXFqGuVlinkSC/tcgwl10Xwi3aKb6TCH2SaQ0M1/A88ejKBdR3/qzW
ZnM4drmYrA6lVMKF5vo07Oo3WxBOhj6QafP4xvM32b1607quCoHkaD0XY0IrmRO6
LeoPbGDvqtwR2bOjQSBE6WhcyFpZEs2yRMLyvNPMipmAhCIB7+80ivEn+RpI3xvl
gPl3jMDRNjIkTR9vWZqxgoaDB3ZQUBdsgUIzktj6m9VfWz7y0hEDoo7hsYORYmrg
1pW0cPnI4yyGN/MnTLIVsD0wLsSy8FDG719QT031xYO7E20Z7iHpQtVK5k8ETCpr
pU9mDXpsorn/NV4vI5E9zq8bpnW1CehRw9qLnzLv3BAn2VM3rPsALyp0zWVmxU4h
T9rGsIKtVFEsebvX3dO11/oHnvlseoeGo7vI7WNcQNVjv6IeqNZ1dwMVidpHbk31
MVXKvGUS+lB5oAAl44p1wA3KEzM1aM0QYAyi153HPjduVzuiGVwXlFR0AcanrrfR
sGhC5TbNxLGMRNoryXsVgGsdRXiy9kBkHM8HYCHnDHl0pyPLyRHq/IQkRU2O2fVc
0YXIebowddvM4Tm2F3CWmeoPu1JvHyq7QUYUKWoSrjB6RsME8fT8qoMUJWH6um/c
nGIm+C57tZnWzoLJCa6BPs8i796JiFm4Qi3tHUqYLQHdd0AUkroPIaOWSBRD2o8B
LIunQIZP/Xhqrm46yJK3lANphiu4VT3MEDT9rc/WzhyegAwZM81ug9ped0NLJlEe
UXOTPKd5IaiKMJLcuY/36QaaOgvzk747TKsY+2bfyBiUNuJ/ae/pA3qaL/16GjtU
ywqrEk9JzsnWODmuvOhREerDEBYfc47steoEgyzd9gP9qTVA8IsTLfGzLffn1h3/
4+mBmGsAXiQSB9Rma69NI7wPudN/8uLPHaGJe7Sug2umEuvuK8sibR7P+hXlWnd9
xyyUAPCz/ejQL6kn5Pz37lZyINRr4fRHpldhalG3BgmrwvMFJCRdzDC8vHllOUjM
LPBV3rtIWk8zdtKtagHwKayJOsjQ+YiSG4QE+fq04vs1WVYuI0t/t/NILJs1BGA0
fdCpyolRnDjksadc9h4FZWdQfbZ6pFazJZSCr5VGKVevKeOX09jUsOH3QZGdY98E
vBeQv85TyuWhRIpIAGTosCnLzlJbWG1sctqKfhpO893ZBmxzarf544IriMRni+8Z
UiXDwm62jMlit3ZHOA3IRfLYu5IdCTLikDxpTpAHyrrKrSBVKZGyZ3lOLa3OuCCT
c0rYoyL6EDo+C4NfkQ0wtgMmdSSgnyDKQUcQbjZqch+RmUjL9cgQUOnXHqmBefp4
Kg426zimx9TIsMYMOkxD3JXms4OKPDsa/gB8IZYI+QNT+vIzgIDlijyrkrEzNx9g
AvMwadZvfDkdWYPT9E1GOW2vy2CexQV6ia1gEK+wBkYqGw3xi0knCVqh/ONlrULW
2xjmIQWOkms0vh34iz9z/6gehUzYwskRBl7kuNRF8sXSO2spqN7gNVhWcg/oo2im
a86176nCzswtGNpru+pTA+yLHjYfoDlF6l313Fii/GVYkwVeA4KC4hqRLpXtcy6B
pqGgA0Jbcf3pLXsswtTGrxnaiYoRlch56gZdUMbYKetnLOCEuM88uIWgzqdJT5pm
+XA8V6hFyB1pcw4vAftBvEABlcCTOisb/0o4J93hf8RxXQWI7b9HOtn5cJ0GliSo
e5onmiEVDxR8MSfo858oxogghRmLrNqOf2xjd6F932VcMaLfyncK0yER/OvNd1WP
1djcdTF1uc1IqeJJU/nZwh3pieSLsoYk80PlJNw16wcbZVDeDQYCtJFDCDaoQ7lN
7KAL78kWo+jEA8U//ydZUkjLVI2Gpu42nrXRirsUer/UHbQcygautvP+7rM16JXF
BGA94poofuyybBxcpTqiPfFNL6xX35wDPP1ZJGTasVKtV7DXZzeye6JhtQAmwrte
7xkKhGQWF+mM+n+3zf2F7R0y7580A4nSc4jaaQd9cQ5kFWYxkem0Xrrhc7/Kulvo
vjEGUoIKvhzpU/8cXzuZVOlds6xb4IAzp821jqN7yRgKEby0DeIhrFgyigedKWFU
fUClzgAMjVs4paCm5cVhFDOkYDka6eH0TvhPl+67ZBx+02Cvji6QeMaKofeH4xB+
yrSBT2l/nvuQXQU2K0P4SE3Z6EPHH1Z0GOVGSYpVpcKKsuw9RAgNtHCOHjJNeMZ6
9J8a2dp8+Ma1/BBukvKmjxJZ3nI1/DTcBeqQFRKPMKuswQE7AROXx2WU88cfAoed
Cu+5lV5iaH/CwKvsKoSG8LipzU7TugHqKSPc788TfSAUyMh3CX7JzR0+dpBGJ6vr
q8nfk7oJNDjD4/M+WudAuaq9JWph+RPiByByQ9RsVl4yOAgf/YSluBCrh49r/8l5
G723LNMVnHiZvWv6TdLu8Xfancv43tSQgm/CgdbDfGNZu6Zh9YH4cPLc23JKxGIh
ogcu5Omc1t1wJyNNur7z6z5o6pBgOd+QQT3tpp658owf3a+fTmnzGJHARw6PV7gm
9swHPHqPcecoG2lKjZkOPEjEC8+20fHn+YVJpsPlwuqodEGobnPXxztR2GP+qrok
hH6a+N0dsilbBqAxqfmE8aNAy70YeNRCTMf97K4FCOcW+knOk1MH1LTfEpiaCIU6
/ho1Kx8pkpaAwPcySr4kYlnK/iul6huT79gG7VNqkKTcb22tppCge38nQkh/hvln
QW9vs/z/UmeyJ+0hAa6xMYNUOWpQXT6F4SAFN7CV53500bCC7goFSMZWW7V1BH/X
2rsO2lOm7dK1KIOHxq9Tx82ud75Ezt66a3rREPzwVYH6OqgmLC8Rq7aull/PjNkm
k9NK1HX92sUmJhAML9MbYmahC+NENALgzsesClzbEXc98a3lXFd++Pnn7jQim+eW
m1y+wfSWl/3pftLNP9CwpvJI3SwjQ9VpP8F25EtCwD/slDTgOch8L4mFBv0TOS+o
gp7kXTpl+Wzq8n7DqEuAs8h+BrM7YtX8ynEHPsKUlb5cmFqw68I1mdywtXaRfjhu
3yn5nqnW861cypCpmmvxuOyhVY3d/Ke1+9AHZztQiNjQOlWZP/bmW5GilFxe9nl8
6UwmM3yWuTHRZF3CFWkSZDUd5FOaK6tA+mS42JzwJofE3RIiOISiAcmdB2szSdWF
KjgmlDPoBO2h5NxPQmql/Z8vp1xEb6RXzJJAyLONqpohGV4ylTqew9dCkw1BfqKY
UnMRMkbMQL3rRewEBf9cfCVhJ+ZMGUiUvwYSqOdJyC6qMBdh2RuAeozTStTPtTaW
k8UyyEa6LlmyK8Vmd0YVvXDG39+/sbTy7Fu7NuUTLu+LhNsGc2JJLywZYhZ4+0D8
p3OL7QWuBrsGE2up/JH124dPgNWzIWQt6hQ6hwUqXWos0j6insldN1pF9SJgQpYl
mLhLBdDqFEvbFpeGMexjwQ7e5EeW4mcilMIbZd+uMd60sdESk738Jrxe2xxEIkxl
Dw1Fq0IlrFDTvO2QFC8RezsoBJ9mvayZtc9FZ4zdH0vlnI7B2AyUAR0GoQWFgY9/
RNkcmHjzuOrGyhDy29pj6hL9ATgbrjJCbCHsHmIK29FbLtyRORA8qLdUEpi8baY5
3prPKaZOOC5qC8EKwaThpMmGasTQz9TEbr8+F3T3YfNfVrUogygv/EscplETD8QX
3KYeQW4LkBsvCvkXqsZq+7UZQNyVmCUoJtn6oK6CD5C5RtTP7JlPakjfg8W26L0O
G0FPfA4oXMFvOb5iCbPILG10phvP6nyggRHpukczv1QR0HGJoeBUxe+atM46+WA6
24JWm2UgF/gxlNhmoTSd8MMtkLjooTlpqyPamB5UVySpmkZi1bLSs4W7gf3++WsL
P1Ve7ErptXJub2/pWjdH/AY6pOmXha5ALpkY+K+VJpOalTOv0DxiL+yfWwxJn0cE
aUgRlQfZUlypcjm3J0ASMKVTCEd4VWPKMFcsugv77gg71Hmkll4axHumE4fBY16Y
AfNZrKMhIs5aoreTNXjQzwnuxWrVIMQLzZfBLn8X6mr/26eEhv0pHqu3EiRqil5j
azlCPrD45/BZQGyZ2BDAByYEXOZsJCBa9WN+C8dISvtvlz0/CfNXWYQ5YSCHTPgP
kRSoudZRRgKiMSXkInd3mYQXCtYyKyYkGOVMIInyXR7zONZZCvlCcK7SlJjcbApm
rqHwJ1D1UWg0YrGEL1YlqW6fMCw5eq1zP90c98io4J+IO5Ir3KFkDTs4zEQ6eejX
CyHO07oNm/oC9OEu7OYPunwIuTr1sx8vj6xG2JYmSwy9LaOch44Mob5jYwpI57fv
S5iDtOllJ4uJlb2CQZ8wgAgW2U42Uks0jrRu8YZcRqUwm6J4euMwwsHeFBvyDFaS
V4cpDfw10VZ3zdOkQqC7lzMME+ES/A2ros0JXusBoMaMWFt8ZP9+tbedESxuzPB3
HBvvlJQFIUd5G0F8jwziLZcjb5E/A9Ja5X/xAYduwmyV/XEiriJud6MxEVaQ49X8
xoMRF/g09FHJXkD+n37jkxfdJA/5gMLFQfbsVtI8m4nKnZh72mqrV9XuN7WOIWCX
/e1Z4YaStMKno43Lfrcwh9O2UOudKnmDx+N+IUMRB6CQYU8Y209pwDo4KqYmnRf3
Ed5889JTU4efBRgHKWfkGYJuU+FcnqsG4M7ZzFolwqdlyIP+XAeYnHngX1Akt616
D8m8IuMqvWN7Gum+xnGCeuiAPyRNTzpxeRjWEdqqZd0NYWfllAH8iN2bS71PGkwa
9skG6LcEalAjJxnmhIeMXh2l+KOc5ngEiD7Xv4hmsScud3NkdcrweXyxkw9InsTH
dMf3g3TZBuJPlPKSV80QiQ1zeW7BprC1TXapEjcBzFvJMNGIQ2vBcV5Qlt/KkukX
gAS1efqp3N5AoviJQJsd5y2hqEq+dBnniiFAzkSDSdf6aEhIHb8vyURMnQYvs7Bn
KNVrMqIy380D2T92j5CHzErb1v/YznSN/TtgoxpZpjZy1uTtGFdK1Q+JwCfeyZLw
5+LbwV++5UijFyDkgoKCdvdZ7U8/r5X4dWt9bmqymSzr0DbW3+oAjvRTXWgrz/gK
E/Ixxkvk5nkxoHw5L8WXLL1eRPOt/keUvCFg5ViDwdrJrfDxqd7tWapseCQu8W8P
tSRE1lTJ6v20and3ifVtkpJ6tpN9GW/khHLT8FbD9g3wTxFaGRn9sGbXCB/T8Mmd
y91RABP3SeVmQxr66Lb9Ri6u6CCZpYNzR/Zlu7LL1yvTK1IfW8ojTZ1AejViPQMn
400+itwBciWeDs5YVHlGb4kbfDLGIDbvOQzX9IcXXWh4Q9mbs+i18rBOsc+G2I0t
kgoD+NzJt87akWl2/XIM44ugpapHl2Ed/dgz0RtJF3uFHuci9y6zkQ+XT/H4OPDC
LEQIbEKl8EGaPz1CG3dlGk0Qv7jQ+bqBMTy7izCzLt6+1vivScYGSe4DY24lYlKq
zT8uecKS+zN2C9t0J9CKSSMWv1wcHZoSeCwaj+Zq8EyU6BYwEuOTSevhBmt2q8H7
oyLeHgqbhvc4FzwrEbr7iFC0sfGVYfpqfBwF89OKQl8nEVykx+HXvtIqDVoGT8nN
RcYnrt4uAcRA8LVIAIplxpISH47yFET8BDx/Dx8zp/rgZrirT0cmU5dYDAabC1B6
/+Fg86XD/TEXN3Z+hwxOXFrEadgwvtvvMbLqVL70CL+USli2i6ZdFfZoMwl0NsEG
y74PR5F3qqaKdERu9K4b1BRHcKR3VhfC7n3KpmUQbbXIyCgH8aOTnh+woa1M5pzd
9ZslDp/4Yv3xkWhxCXY5WECCiCooky7HPzz3Ju6HEubGcduJRkh2lPesjYLr07+E
wwP69aJQOfbszEki1Zp4uvkSsAO+HYSjhresI/prMGkUDAISixr14707mqBMHaj5
ZMuoXh2LxXifyqUm5ZILKgWogLk9Q30qhp4HTr13t5f5+mLHUsiyu75/LcdCPVNE
kmQsUx0Pe9mZTC2me++BBFrbOE2omv7ASR/4dlACytuT7kMPcbvWDI85a+qggNDk
Z168Aatea7crWbL2H882dW73yvlO0utegm8JYZb8h5g7jD0c4H1vcysKER7kr0n/
Ng/xEYkYLFHTBVOnj/vcHDgCT/3prK1ivCIEGnAp7wFkzc4DUUzyezie5WfQeaAi
3vFbTtof/KBfS11+wzbgWASEWoHTdHa7ys+fkJA39aqs2bdVvJBLyoPRwln31V4k
GK8NY1CqW4fDFsI7HetK28ziDfSdYNSPDfh3LiCmLlTbXMa0ofgJvqETfBP1GXu7
+Q1s6iyzl1diEpal4D29YU2XjuJPw/x0dH2h9LWBxDksQpU72OWPEg2Mgdk1V+bB
OvqwxD4c7rp7fUlzIqgGhszn0Gc/pQEwHswmNjLjUQP3Fzby+lX/tKDB5Gx2+Wtq
2k32cC6x9kmiSyZ1ly8LuSigraxNzycox4v+Ii6vxm9JJajskfQgEy4/kbTHWfq9
3UTf0smGl6BHG1+jm70PE2wEi/xHkH06pnsNDt2c42fRtmuPSbxOKHxX1E+3fSMD
8PCSWpkOXcA+A6rqTReFFercgeNnYXDkxUtMe3rlDk7QTXUpycto/D4VK9xIfx0v
Je4oOhxRMNUs50mShoe6dQAiSXDYpapgznXRBkaZSlcwzaf7hd6vtSf4iIenFjC7
Qgt+rGr9qp32Bvl5dLvQONtgdeJYhfr1SjNQhX7JmAcAju4c4bbKnBQQwv+Vm64V
QG+oFxeSgTUcppMWlMQwSCjjDjZtPHh0nwG/vuE2kl1ZDaWCZhQfeBaJz9frUlt6
ESYqnHMmroXQ8KnSZeWuaB32nhM6QusdUSyBBa+Hd7xP46QIvMg1ugW5pvWpHw+P
HSQUMEWozMp2F/hsdRj9zcdPyL0oLhHtKGbBaDTvtxWoEByrPjZu376Cl8Km7CyK
sSfDrFBS9dKvmUfq1LlS9cL7+z6LhMqey3Q3GagI3BVAdzLMafq4V/8iJ2kCnEBP
bpBNgCCUF5aW4z05KJfN7ROTZMx7j1AMPGZawoJoElajXvfWIdjYdXRh6BMK4N15
Tae0g98ayV3xSkrWmR9IyzQlQbNOuIDZAI5zljq3utZwmS53rxpMdDDeAewMhj30
4naAUim/6rbHNRkjkLw5nh259+OOiLpBZLEYvHEqC4Bh4y7cynlfOJMKdVyK3nL8
OK9zUP7MpV2KqNbnzJU7WWB9OC1+A3DXUh5TFmRGHPHALOO/lyqQzFCIfLBH95dY
CRr1Al8qOXE7OZbEqkopPtEjncQGZbSdI5A/lQuEl2iNt+usqd20QS7bm+zaKNY5
Huam6op9G8REm7As4AVJljdWz98E2WIU6wUzX8FE3JKi/4x6uleNUNX6y9c6DAVr
ueBX9SsJW7LVwuSw6fqbaFbPqlSCQ40LaYUs/gHa2TUZ/sdsxww08x4JnsIB/XoJ
N9XlRlLmxihc+gSMJTiu1MdCUjKPtrCHnbilsxtLKclkg3Z0vZXRU+w8TS5FQIfc
TfEd8o5FyPGar26d+v3Pvo2Xk/8ooCYkQGdoUKMt4hXWJiNmQMSpiZCf9ik7b0kY
uHL6HJ9654mVDnYbIcc5Lp5HwFbNr7/CyaPC0WItRfdEsuuRMpS1/lomhCOkgvxh
Clusrj48vhFNBfi4Gkl5Q2KkfqRBrdPPsXnLSullQrCFNA462XjYlDyUYNz0tD1B
EcjUgHClOi+HEAUVT6hRJVCxG8COdhKe0Bl7g3H1wsn/SWREyQaOunzqGFHPBhY0
ckbT3Pj5WtXGiUSJH18gANQZkfE+hg+sDf7LVgrqVzgtuxamcZ+OE6CDYRaxHu0D
QJ8GwfgdbJcmpxXCNNrDmxA2dQs4Fw72chFZ9+fLqQfM9mLfGzN63LC9RvTFrGHW
hTrWQ9zBbV7HU2iPnItTck2CAYcbJH17U177BOAs7UFDqfKj94tNkV9drJPXcyfl
k+wRLmsbq76GVrTY+qiVCTG/xuIGmq97052/JJZXwKqYwmkCVxSnba9xuseOf6tS
kGZ5eEAtCmYFKj7FnvsAdZxADjrw4mWdNWJ7m3EYaDsWvay+3899zVQLTUuLs8e8
vHPCEDUkF4a7XsMenXLv71vBbXiD7kVf7TiR3miKpcvTv5PoBlFmlN0rQMij54rn
7/QY1zE9+9QPzSNa5xOsfWx/oJiEj3JNiW1vB0Bu3K1m1Iocy2AEhsiMCaGC4AZB
fpVMRk+OE/T7bOE+9l3ZTZjwyjowczoCVLTlcp5IXp9tX3gfotxzQZLYZUi5KEdW
kZOJqhHSz5Wc/RSrZWRNIMMedAHIbrMHHyi/v9McdABkPG3BkPPO131oAXhkBPT0
8iVGaccl2kWMQ8xArpSW+iDpvS1q0+0nRCd7Vd464LDkwenuhxfM7X2sbtH7vBsc
AEGKoKepuTE0NKEWI0Y3ZXAtMh5zjUh5262Gz6aaM418++ER4588L6KWZgp5PJow
ZO+YI8fyD0YjosFkXmUYegcDJ/faxnKB4md0YK9rFa2BKBAGAp9l2lyZ/uwqz40s
3URxylqo0s0TgK4kiGIcm9B1JTLTLa4C1rZM+eXnpxIAaNM1qL+pzby6Y6P5tJ0M
D6arIvRtSuvfhyVSwaren6Vz0SMONbVXBlkx7dMMfguAjYmUC9aG6mddd4z5lrhw
vSL3hLMw09BE8gWu12ApSUGhXAcL9R2pXYBObVt2QrAQIrFehiLQTVXb6EyFzd6p
/+sdnOtopX4cMWiP7GjdLUI8i3dQjFbO9n5JO0Z6Rx4mw4vGI9+q+j3kYud7T0E9
aglgXHLR8rOPjvTZOeKiCa8iNhUx0R3VihmIuSoMvAzJ0+rTo8I395OqIokZ6eTf
Hbld9B51a6Y2nX2F06NoT4gFm3usVB90ltWnjtR67wqRaaHEn7m8GbvxbBggQ2F4
gh7KWCSUta40ftHTNzaniBWr54sP1Lf7vJeXWjh060t3dCHbC7JfpV3SXfCEy/fk
HVSHL+49tNZw13yZJmihgTF8HritI76Xt6Iik5hOrQvbpYu1FNjKTQYHlbXJRD7e
FdXTf530OGa31a6c5dALxT6zyDxSk377WE1sPzYDJI4159sYBtNrZEfChP+jhdaP
oFqB5Stdlv/zOhP3SIW21/KvSDHr4v9bAtJeUyCUAAW8ZlzbEwxfDDhdfL+6F49m
d67qj5zhDp8BTEHcrecAN6DChw2CE5g5B7Pjap8E9HIq7EDTIHckP5fYKY642i77
53jBLzoYX5HlHG8jBS5ZxaGiIO/bcdTuuhFHIjLOmcBWPwdiGYM3uqt9XAsNOdAb
NivU0ceW8tKD/IJ0Dvn1PZWFwJWC1qP37PUkza1kbpRKlkWGwUN0nTvUCo/qWQEi
oJJkXNhRCGyKZpVfTycwienYO5/W/i1Ob4HDrQkxbCu2whds76vPfygu0NSL6Zqw
Yb/pfN77yPYccOH7z7goqfBnmbGgbsBOiau1dKOmOTp1uYt981Dy49kEdov5SBn8
/3kG+36wEPQuW83sqj/2EI6+tdwIoEp8ogUPZTY8FrdEErJziHU4lBw59fl45X0u
gYjsp/+z9TrYF2BT3F+roJSwICHFT0yA0/oRksSDgZStiv2yfGSI+4/bOWbLuiBb
tk7WxSXUSGdRTPNyu+x06hlNij3dx9CIN/kNiGXdPwcSmerpKNAJg2DyFshgfg50
k6KlCHdSNiAbG5yvbXlr+1NExYBZFBRYvDIogVWNLFNqFvCLP65cnVrHRD89k21s
H1TYuDeTgx4VCDcUAn7RAPvxze5wpRA47AbaNTI54mpexq/lEVqpbW7pKR0laRFK
gTw0bMF1zrJqYx4iRSSXTUfeYvqCl6j0QKAQgdk2sZdikzMhA69P69pkEjDuL4T9
22+erJq+9uiWvfrZD423h9rYc/6+EvTLJvft2y/59LLOU/fzqfgO/nSKR+BcYZgu
XoWC7C2GoE6GKUVaYHBE4+KVSRejAJUxGxGgJW5rgGSXfUPKOZ+3EOLLBTBf4mjQ
KJbFksXm3ejlThG9+vWMxNGgVWPoZES6Vo7MzJq8SAyxG8kFWxXq674imFUIokBo
B0v7kAMQNG32bFYb/t2cMudrN41FenoR3VgpQiWa5ScWsJFerDeWyyIxNodIH8Q7
itchODgdNufMKzmQ9qL11+HnjEk9x//OOplUDH6b5xA/H38qJBJDoegTdEsSKMM2
wgxm7DrAVLb9IfARIJH2JP/OYbZTx5y7N64X/ddNkWgSoeSKRzM1ErCcsgBTyJWA
rvJLpVS/4O85GYnShP4iWE5Y1NoL9KKT0HzAhzTmsKotvSsMAxj/FEDNWFcvPkCH
8bvyYgEZoyvxavsBGjJ6h22pNPAmmKXSAQxPUCOwhtfz+dQnVvKxygMllOz83DYe
lnAwzNBsUMLP/ubewhgFYFGl7JwLPuWT5Q3XEMrUhEYuH/drNL82AfHXaVy5IfzV
QOY/Zus+5lGIwQjF9GeHVOEgsgBgz2MTAzbJ/T3yI75HAqZDM7c0LLKa4/JTBFdk
xqAj8aSSZwC6os7R5RrI3kS3RcA70gtDS1ejWH1GOqBspK+j/3AcBffWjOTRsyIg
bOkjvcRDNGSVE6XFK1vfz2lqOe0x44R1P6uDYtAZ2pOYUISlcyM/YjDJ+hlMKIei
9Y2tf3p6lUvTTSgrjmTbnkfSEd3LrkM4016UUgqvukcZMm99jquX6SmrlLHxvG4P
cSN2RgINSIotAUNIO3AANvpQTy5BX0IHiqi+WpIj9ap9asVwHC9/qCiMdaAIKB96
6pMUj6CU5LvOt4+vmWyycHoAUgYG/UN5rR9fbRBzjzEeDTCvOV/FN9rcNQCZbzOI
RzFFNRE2hPjJ3wDMOWyNTQzC4Jk935yHlqyC41fd8KkTs7S289reKHioZ1U/tCeK
BP+RQ+G6yeCyCLWKo2gbXOs+fV6VwkEJGdnrRMQWcg8hEZjuBn/Edyfl8bWONvzC
lxKIHJiCenvoc0pSd5TTBFKVT33DxasbWdpL97xis5SRlH2rzSPrcANdvj5G2dik
XJoMhecykhzf/LLOI3XR4HI2Q9TS0S+vwgll0wba1kaTHGyj9NseMJr2E9VflwFX
z0mIXfWqWEYDWplhfD/P9kVJea9foT8mxqGyyCS60X/p2L5a0kLllgVQBou5F+oO
DDy65sLRvh+pbu0oTWAS33jw4AKRXIvf0W2DjOa+mZC+cJb+RF8ksh8w2IJE7QFr
9J66JTPe7etZA9tyvtnIFISTUkl48I8pJwvYnkcVNf0oktMT+DjF1lTy7S8uaa5H
hHkK7ch/kHrsr3hLjyKxBNfmA0LILTjg1n9+3fRLXI5HuHd7Xm8YA1AhBxj3NaHs
85wuCrXxZdQrF/Z7gfA38Zt0PgKyLh1DAhJy3IMRsv9+i6IWmVpsVJPu3mzaWfSU
i9IAC9zIfJqClW/MSNZGH+Im7brIUdmcfsd+FezmCPp+vTzURcvd6HK90DgUUxYE
MAcSwKyLKeXkQxX145XBs52NeuVRiAUULb6IV+LX9TDCxM+s+ViFolg2nm9uu4pI
uv0eHgtZaalGy32p9MyJOEKvYG+IWjPbjN6K3ooJ+bs37GMne+e78HpPxD3d+YBN
akkWIL4DDevHXaCeHqnQs99axBxvogkev6bu7yydsN6sznqocDSKvIi7etkmLV1J
eSJbkab6AyWyQCTFRsMEWJqRqYEQ13iShkVaSqjY0k5orqxtKmh4D85R+keltIRZ
8mpziB8AR8klSSJq2TVwDosTvUzTTcI5j47yp348YA9Zy/cQvMt81ZLgPNMjo1gA
+hM6eikLfuGGBbbeYmGbXoAfkwSJFlVRcXTnIgR6TqaUt81zVVRS9PfPT2OKhveF
PD/cAFZVP82dVCJA7JXd85Hn67yUmDPwPbRoLzmNd7xHXeOdps7HfsjViKU8eEpN
aar9Y/SoaAX+2Nu4QQXVujPbsf96BECvizzbD+2lWvzUWPpgqzUcfNqBpjwbC15k
juA8TfPQYuKiOdexnYP0KpjQdD/mQl840XmTJEDe73nT6B5qGCWJAIz91/+x/78U
fug6ZE+Nn/aNn0bjdXJnwb5AEI1730O8U96U8OvQdUEdoc8CzYaayGgGi4UQxwGO
3SmgDWJsqrWgEhgn9Zjj9nXzv/Qm5hUo5ETLnXfkQKHE5QHIo0Dxu103+gd/rw+B
o4BqIDOYUnB0tp607YQlH0X3eAhgKYECpe7TlT92WzDUsEuGaJU4uLe1xi/hOHE2
6Yz4Hf3TFuZdSfc5QdjAS0CPggzAbnP4eOpbnEb8U875fAFLAJwOGtrqGGdZvnju
YX/xClDU+EDVSSePCwLRyMJ7JYZzin/miEemb8vXlrbPHulyIAnfbigbdXXIr9yO
NgV+l4mnJsicwfo14vnWanZ/9bqmlxshY3lwCrsOIz2nLdBAyX4rrbkmZXrEGjLr
tBAjopMg8XjQy5uOq5n3e9sg2fNdo9lgi40McGkRMktygoImwrhsb28DxDm8MDiw
Rajq68Q23yy5tATUp6qac5vNOzEbc37rR6JbZVEtqCEhK8rV2Nb3REhhICCcjzDx
9Vy1nLxjPvYs38ADBsHO/PLa+M7Fo/uLrLeevL9ytRWhMrqwbsOjX2oTKIz2gRL9
hFzyuIyCAn7ARw4JlFSbzMTCVPW1wRbw8OV8OCFRQoXsnE3UbyVFarNOKiejvnaJ
DTHCiAeUpZxTUcxf3hdjqjoWTdHHqO9o8lj+XD9XUksM3G7l7Gkl+kBxD5Xm75WE
F+xlMOekNedE/5XYXohSSYXHUKHMy6j7gmLhWBQgM5Cbeuz6eftu/6JgqI601tqP
v0y8mhLUVCoci2ulZhOm0TEo5uMPzD/Dbvy+2ZN69VxNJLGzrlY2KhiMj5PNwc+2
ykKXuoydakk+Qa0gcVFMX/g2cEIXAejEtflqrtHup3sJUU86CuSHbDX4KryrATEQ
hKCNdSZC8USb/zU2jXbMoI7rSxqkRKIqUOIoUEV/QUJwPMczM/n1Uz6ON6ACwMfc
0rvnNXnENgIvuKzZaX4oGuKqNW2ZqHxIMF4yGBm8pM9vrmthZoQA7xAztEMfww7S
P5iFZhGKSf0auzg0YCaCCbggbvTl6kyEeeoDvb+0PLjACQyn0NAkB6lxDaZGFA0B
7FXgtLJb1fRr/Pa7tWhzOwbEP0HK4BCmwMEVVuhOX+HvtvkAeI/RjRNw4+5PTWgm
76JvY4AvbN3ICwZdrapBdp1tRF6EfadOcKsUquuTwLp96dIM9ddLK2ceBQrXhOTt
hAaH5wzBADKdAFvyRLr8UBEcD98+YiZIDyFSA+S0CNCd0mB2sK9LsQDwqVZ4U3Hp
u3GDgTjUgETJB/nBQ5Mn5ZmbvePZiY3/015qUppH0YHE/xRE+jkjGlWwUvAmHdQt
QfE9rvGI2+mcQA1JHvI/CUJiLuCj098Xt9I09xNo79EPd/F/12l1t+LonJoBpfpz
8zs2LsOtZOT8WnUSovWiCKp46o0fKUZ0ITvluI9uU76JE9J+/zF2l4XOyjQGWajD
lHF/qgcPbuzC1TsUVWUfADml9abDtx2bpFzP+TEkFjx3I28ROphtkIKghJhcEGWV
726GvvTO1pHY0/WPqHWPVPJQa1p/UcNpMhi1OFAXMzkHgYNyfy4BKOWWzR3U2BgH
dokcAQJgDAxJQriUHQJmz6MiWvAMuDqhg6/l6e/hQnzHgaP4tSMpbOolRJduc4fp
TaKCTR3+ogRj+hzVC+bLQSknde7YNrN+lM/X3nFXxHOaC9D2BVa3c4KO4yrAv8z9
Kk6eYmNcGo7A/vAoN+X5J++diIm+BdrS9TL3rdFgZgQCzp5lsNpIDTUT7gM3d2BS
Ld0ATOYcPJ4RnU2UI9nNahf4Bq9FaB+p9WwWNU1zqdXbQchuC/JzTHukB/8FAWxw
SxBKaFVAbsGfJoDEr+MsLmgBt3fec/7+uOo4qGxlQF1RfvGRn1S2WwYNB80sF2Fg
KV+oP942GuhZBo++zvwBiEQwvrmqRfHmwejzQ9TPKL/4+6kQP1fjpN/ZS3LKDDLU
39TIkxSnXCnwvktOBdys0zQkffkdTTDqYqybdQGTn0oCyPZzxdY3QVZEX7igp+P4
StWFuLfdoZhln4BKoN7nj+EN99s3YruJ81beCxfCEPKJjRhiFgMr5NUTo2+JTx+y
l+DTzG660dYa2ft94KTqPYQYSgccFrxY/htpOiYx/0XftVa+nDE4JtN3xYZ+6E3l
uOSxWfYePfyg2OeTgwM0cr7E5CVPVlKpfLuo0wBRvnehQ2Q9f9LFal1fZ+b8PLB/
Iv8GZDcjS3C39v+qUQ/AqI0BnhmShrh2M58Ut8GbUI2ww7VPimhG4CXouRPd7U9/
XsOwJo1eIivjCeGFru/n6SVtvzrkwi0coXQkzpUdwAo3Md6c0ENuK27/yG9FmKYV
QJTViYlcxB5Gu/5NpITrfgg8A9n4KreUzapaV8HF3uyoHGYFT/27Sc6zhmvSIVs5
c3hFnpm7e82TkwR6FqrylNULXbKCh9juZ6nklI5QHPhNUhX/kRCAr7m/sWTe0EO2
IGE7iatm+PGQg4omQ0QPaHAD6Mmb4luaRjgSp0WdjSEF/r3SemTpDJq7lFk4vXR4
DsF3vNApCE2f6k9/CoB41xfnKr7a6ojGZjYdGmijn9Upc3DshegUD9ju3wVJxyr/
y0B8puWPrPMgNJVhx4l6ClaC2s8LFD4YCO4c8PDXqpRmtcgksbNuIff7iJgNf/1G
7qscU8ZE6x7lh3YBFEH68gwtjtOWoKzxUhSil9bc1sUtRFMaGi5Slm3FR5jb/ZcP
PgPPnPiyQwiQLmEfMXOO8VM+j1qYEUIYpSJMRHWDmZYJLzo/jHw/S0BFY/MERle2
nDMNHvciiUZQxwkSsJKKgGjBiOR0m2k0I9vv0Sull/k39EMlPBjWPvm3dh1WQJuI
2VOfQxXCQYCXJftElRHutnfNQ0L9fJxs58bWh5QDY3bp13J8bx3ZpFlwq/O7jmyi
4hgKU8+keHyrC9++bI0Fquy1WHBUhgshqWOLuBkGx+d8A9XjsThb9rEWxCWjAR04
PqXCaiw5XoFN/4tFLVMlB0veNc96qXTBkCzLUoM59LLtHZhzkXDy9ts7kfEIUeCg
AEIJ+xjOovykQo63Q7dZJVEOGr10pP4GFPLTmyrFI8DZdUBL+bKzcTUT48TI5aRo
M0XsyH1ez2QSWknB8WJWhjPtWmaFjeaywGi5054hM9W2m4wOFEkqDrGs4XIJavO3
uDMflugtaYCHAWuRB3nHqvyITjPeYAzw/GiTH4N55FQIBvJZePpOHTVCtq4u6Cw0
TIIlhUHhf/uLCJtTvecLcCCbqBZy4Lkr9BylupiuzFU9hLPzdFcmTVx2/KhfczX+
/OrF2uyIevKmGp5XCPxJBGuIdJ2LznhnOoJfFyNEmlEhO7SaACcAVhOlTg3oa44Q
WYAhgkrK1bm8OuGur1iSPy46PjpndRy2N1Qp+6KHaJoEI7Xg/eKP+BQC7g98HQ2F
EsmrWtSMECLFXwKP5+g08hVSt2qoXtfT8KPuKnq6PIR/vaT3980gKB/upQqLVjIW
EaX/EswqeUYChMY0DzrxOt/5pANKh7uoKe+nXryb3lp+RXmMTjtErnbOmscBAZ16
zpDfDOzNAvM6YfGCgI8VgwEwDR0LYDg7ikcMN0UoSi2Nyz0X9eylIBoMHj8GXxot
9uK0rOKYaDUA5UCNHgwI4Wp+DJxtEuXfK78Z0lxAQ2vOkoLWNqWKFdCZPSVTCtXD
ym1/JnJNSj3As41TAyOsn+ZUpGRfqdLY+CoUim0oUgteW5ywvYUV6nGn2Qw1Qb67
oe95fSBmgjG3Xfe8OdgaiXGgaWUPf0Idi/9PN3upU5l3p33Cgo3Lm7q+WnTiSgNj
hyki+//x7FNIoSuzmbBiqn8nBiFjwhgsKQA3Qcwc9rpdZw5c8LKx9hm79EBCbrm4
CzLL+AIs+9DJEkJqmcf3p+2DIX9ACaI94JGL3fQVXv/d+/ClfoEbt76q3U9l+XM6
qWkPEh5EzL8TDTUxpgqTlVH/kP+xBlnWMfkJtckYBBebSuuaXwTpIDZLsXxNxoTs
E6zp6Cbabc4Kag3AFVCffiMmuneKgIpDAQZgg39jLRr191GOvXQWCHeG6a80uQEd
S1xdl54+YxKaIwSeuko27UCiuvI9yL1R2A9Tqv/5pbzfhVt9FogsAOJfdZHrh/5Q
Re90pGleLFLiAe9E8Oi8/mE+OO8qomqC/Qvg8gpvep8M5Xt1zNwJdyucqF9EgsS4
QNdS6/Gb+OZqFXbtvKNfRvVCtNaJQyr51pdnn64sX6hWnD7ExmFLkFsyG+Lm/2DI
fFX2sOrZUs/pbQtrP/0km4/awKFRMHm3tCzLkd0WMwwZcvCbaKgVyVTKuE8xt0Vu
xfUVUYQL7wHVAQvDZPPdGZk8qlpTleiGcWBn2LaJL20lRsU8bsw+Ez4pZVB+kgMT
E/TNZYa4TtuvsaX3O2o7+LQSIAA6e//wg2aBK5iDScBEc0dRgd9i39gj08K+p6+f
acRg9BTu497ZLD3tZJXcQJYqXgaMlqqPUeBn8Q7QT1xn8p2oyKZOJQNAFfqfL1EU
JyzVQyeqh6aIb55JWSiOGqIEJGnQ4ZtMGUzlcADkDoqWH/9b6TrLYXZ9RVt2DirV
nVx+RXslmNn7G5tJHiJeDsCpQ9ym52ySK0H71z9RiliJGBOzTFK8U3fHOeTan4C0
STxJYErDZfuonKPa5hAGzdEbZv0Uhs0JazJzCIleGunIeuqlap6R/6WRjeDSJzaD
B95TnznKLmq4s4Ty+0t1nkjGgyzoe9p3eEis8lj6yu6sejICVE3Yg3WK2Sb1ysyA
DEIuZ2R8rGBG1Goba+iypBZoyygGuhkTjd4YBEyHsYbrC4RI1DGZ14Ck4RdlMRP6
pcz84c3lvPvRdZFmFOcxYSci2+cM0ivW8md85enlqIdPbbzTDajMPrf/SjC4fMoZ
/Tmab2gVXzdHgzTstqz9YGswoDV/vGhctNiju+2ytzwLR5yPbLjh0lhJ2f7pkgro
/boKQxxXgwxZhBOCRM3/gcYzOEkv5aB5sVDGmLzY8sYTMIDoNQoVZVwfIVxImcP3
d3aoA7iiFvUh0AbsLKi9uMfFj07P/Gwrg91Y/qyQrgY80iHIRpJmChywvPVN+28/
4GPGqxt9fIaixt8h9iC1wkkDdH0+HEtULNPmDMlyUKtIfcep3ALMdPYs/6m05LAG
72HcFgf5OYC5w8n/ODXXXa+Pkrq1EloeQPUTaNY8xabCWPSVHjo3lxENWb5a16ew
UZLBU1QFYjcjkDxPRQpIlVkau/NEpFlWDLAEAjXnKBQzOnjzVrpqtOkXBuI8m+xO
X+O3udKySn5JsaX6XSEu4rxOAu8V9oFbDi6Skvk6RqapRXX4dxbo19wN2VM+r84p
q0hh2XtYNrkgEj70DFPvmYE8TqdgcNHSaSqKsGg9rj8WUWCE3piFLAYUuC+sc0P1
HHSWugnpYYYW3qScTuJJ/ycZ+2UEqGuiX6dbLxH0TcPa0L0MRDBZ6mojYGt/Pf7d
8V/uxeXvFVqbyMMsxM1Y8nnDatCPG6niBvmpzwYdQFABchyxjiyz6c+C78wjqjRa
C7Nfdj+TPBJomq4IGJyClHVJpboNJsiyL6kRx7Czf4sFPYGsvT4N/6ytGlKyy42q
qis/APD2LUKm7RpqemxLoMT3i7cd+A+lQNw+7hpOwyPIO+uy7CNwPRbwrypQ666t
F11qtCyl/GlpnCyzfQpzOHzv8vKpMpm7ENjfCBkqCaDwuR1fwCVwlxwWA3yfhNWv
edF+YyUwXH8cHCO3V0nhiVf3CNT+ojKQwMvUGwMFhUELjbzNcK9bPbCMtCQwMlXi
fzbGzJpX9DxOyveiwb6KiLnXZUVeA/QBtZ0pjYXmVwRUOHhPKVfkghXwuy5/obUw
jRnv5XbmGIgL9LXkqkq67gb8odspf7l9a5Qh58sjS1SgQI4ZPk+BXUDKpDSKiGJ+
hwqjxHDsaX6/vIs/Q/dafuuP3rUTiefJKvaZ3+yRLtk1Cf4kGZ6+M3qrf/61MGJG
gnl3xGj4qH/WJtWuNFi8aNKNYCMQ3eQDwC3qhjn12PzzLO76vhuL9iPMKofJmVZ9
82SB9C2ViOVZHxEnbYvevEMOYNVqt5bbwyIE/gMFw5r1Olgz2A/CXVTtPB2fOapk
V/+qIH9G0ofbWHCf2cOooO1QPoH95AAp4dukOJGBdfy4Z1bMw2zejt4pVHqNHb8Q
ERP+dGfpeKkWo6mivqNdieBb+zY/Cyt64nFloZGQY7YkKX62N3iwP9a0pItc4W6j
UMYNZKSSnrL3lIAydbwKrf0IS/bJiytTREHDcnjMKHPFGTocNNfZLkN7Yp3P0Dez
Ofu22vtV8Xg4XyyLH0HKqrhMSGIU9mFS9ykepOyFfit3IKnLWgaLeeIca1Dy/CiY
nU+U35kUE5JDLRBBIMK+f1dc0eQFpy0JKCGydstccDxiaxIVcOnK+6fVF/x9z2/D
T9XNqwPz8HI1MCsPzctx3Fr20v5iTkbHJl4wChY+xGheQfB5jJBtVyRFo/IkkKFg
AFT2sh1Hfx7/c94lZ1lc/7g+ZXJ3xQJerXsq0MfM3r/hSsLSZhvUdX7g/yfv+/9Z
aToYSuwk5ddGVUDSlgOzl90XnY6bJAGnTntakCit/uGZGFOBiOZHh2VGbDPPiA3d
aRlhX55JAwhHNjiNyB+o/e4gEOm9ArevlAGJF3gVi0IePhYVnoDRjsbMT2RodpJU
FCAnWp7WRjGDk/U66iWm84XHwNjbl++ruwbNV1vY5OvsUbDS30gEd8cAkvzhsO1y
3QQsRIltlqefvtoQfTxSf7GTuYq6mjHIpM5q1H7r3EGrtinOrwzRa+kwdSJ1Irgo
0zpzQuqZaMzLBWnsiHsOU5Dw241Wrh6GzlIJUiKAbZpk8j4cfwKzHVsDWrwY1xgi
ZNV+4q6E41EQI3QGLcHVj8C3O4m1bw6qkgcuwVwzAXTEa8vbKQ3AdGG1VrNdGeRA
i81KYlZPNfuhnj5GGK5FmdDYWjRmVsWVRiDrGkdohaMrlFO4iXtE62FStniwqy4Z
E2xjHbQxpqyF6StAQT2eayYNuJb8vUQabOaKUaCh7knNc0U/g6OZczREuXEKmTLd
v4nt43meYDu+cpVMoq7Ny7+Wukay5vIwBZWKCnKZT9bxi8ai7lb+QqMATwMvagEI
+ljOcldEOTabduXq4Fyphv+Nn01+mvjYrMSTS3QMkaCkZekAjmg/szV7a3kWqG4n
F/6kd5KdEq3wra534az2YI7HHJVnsWmzezHCiFWLGGQbmBa1OMw9uU+/gtyKWnaD
v44DurujfJQhaR6JpCb5YsRIvXeRvKpoIdTKdLrEGBnuBUvUNoVuCLfSccuJdb3x
3ZLl9EgBhxKRQGcwnCWgIpXr1/BsrNWOser5ExjkXIH6kraDyqkpKEQSYhDy8TQY
vBEsVXqQQL6ABMq8b9muzpfFqUt+Qlje8Rdmj6wgBRDLABeJUPh+af/7enKbzBaJ
fYTTSC1gZUbidhSnLFfnoLzuBThY7F8lPYuptVv9kZm81yOD1Gq8pIqaIELtXSX9
aayX8//bTnR4bd6kHsJ2OLTW88z7vlM6CnhsUP/c5DaokIe8vkpS4N+0y/DTwagF
BMS3RQ453dViHkAL+kC4eEDupp7REM1IFs15R/fstGiVo8jTETVYIYyzHeKAKD6v
X3//WdUnbBz1SE4Jau0j+2oJpJ7vK+lHsiQBiI8bDA1MsphbqAbJ23zBD0u9kXXN
pqeyn4S9Ivd2hgSP3VMl0j5FXJkjzwwD2+NzgL+BQRlpd1Uh/HGOZHZ8408Ab6IQ
C76hOqlNqOoa51OmyYe+1f015Otg4zAUr2chc+I3/ssXTV0pE7WZJxeljWKmwuK7
3WspvXMOha1heNSBrrkDuF0TShft62YyykP+PhzYsJ30O69dz/DMuRPBNdFOK22X
4XfFqSV9lHOGy4nJhu+RXg3FU/vKW8BuCrKEKQcfDpJjJvmZ5+c9z1rbJZI534kB
wJ703IhXfj8QF46DzVxVIP1M+qY53maDqPZ/kcmTCJWORsBVvroSuPDXfX2OKswh
TycHhmS+a9DmF3PSAsBXNdme0p1w8sGOU9nxkOZaIrepAK14XpAk2zTxgcxpd21b
d1xUDBYkCKvfloG29D329fiIZkjx9eaTCTbV0W0+idtT6o6DRvMEejfyTaW4euDO
6yOckXnZExqnldfC+7dmPbEsV34ixUa+txwnUOzME9KurefXrn3GUFR3U7xzKdH2
U8vkJY/ZT2XPbrl+y7sr6/cIxPrMie7bd4U3YhCnW2QW0g65+fupUAbOEOzmJhgL
qUMfOXFwWMrx8O04IKSPV0MEzrygv2Otz7vOkW7iG9bhyphiHIss7FMtxEW9ECxR
y6drt9iiI2607FwauLpElv3r1scoQ1m4Tee504feYKv1gr7MZK4trTN/biQehqXf
nk3ZrFHJJmGMf+1qfRtA4QO5cpgB06xHVtr/6Cf5bLJIueyuypyGX4j0UGIysDft
2niGftU7zH8rYY75qSNWhldfqzGqezGXy8/0w9pv8GPkfx4R4LeGGDMbIFucwiv8
nwDAXZSHfD+pLPXYQC52khJtpQ5LbTcoxewxkaa7MVwIoWgq8mhLuSlmEmJPgm6G
S9iWVoheQhEpCKH3g0oBaxuQaXk/yjL3avsHYEXAO+jJt7t+kyL95q5YD5gmR7xV
WnAMOrVsdDGdzhc0NeihlIEigutntA63+U6sxGNWwn8=
`protect END_PROTECTED
