`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaltUHWIBwxBz9xpY3TQnoO1a8AzL/El0FlLSesK8BiXztoqGMTsf84qd85wO4d6
vVRoQahxltGBkm3CnWGRFKgE7kqvLjCrqDOpRY08SUyvgNYZBvJ7CLaPFa5RXWeB
DhlsC5DIyfOi6HaggMOKeSOps9OU0ywVxHj2QIEVMicfRJa6a2OsiJmJyla8ekPM
lDNNzZdN85vevMcVHDpo4iI6yhwPtVilqQSaPeLulF9reIWAF0hUPj8spIADuPO2
WD3ta3asR9fUYVvMn21ODAowcWIOr3SbfCEde2BtvAVUmtx++g+WPr4p61BFuqNL
PBvt/QrtHZAQVQtm3qzK/EHhzxsxXIZjvadK+JerKmKeFvlYgpieAI2aO75OaOpB
L8TnRRgGR3UC7N6ZyIZYcscaqWVbGzL9VM+97wUihdFzISPeJNyEh1j9wNoW1FN5
a/VGBBa+qbK4R5Amo2hBGzl4BJJjGodtysUMn4Mv8xuM56KHot+a/NL40ceGdR75
ghNGOu8bg7IG8T1N9pO+0ndalkR0a+jMK1vWotQsMkFmU08+UiWdZ3B19m1YGf/r
9IM/eO3Cu1nsH4G1bgRUbmtsZ++XFJwYeGdOgTSqQmeAX+NFMi7mutyRss1bfNyw
er3KHYR+3V/tmL8RHSe0S4+Vh3l83lnvr2p42pYSJggF+Y8ncMqWdQokuSflVl+v
K1TEqF8Nj+Ao5XzGaiBXgEZAfwnz6gPwd+Ic+vRRhzlYwu+fRGysr7bN2xVZCxCf
POJShBjgk9M/shRMZ1FtuHx0Tg5uWl6mC/f1uTa4HKzmo3t3tE7n86XahnfQ0qH/
elpLUCdc49gO4xMkl41W/uQ0JqYVQ7w3acwJaLCrZ1IzwFJwMpgLLp1fLP6EWjtx
9+ouYYDlAzyslwyEFcz6MRUhH9OTQYpVPBkFYeNt9lUdqeanJUDjqg8ZX0JTI3vV
iat82sIHrBeYlbZxHf+9Zl6A0OT2FkTGkdd04Y2I43KuauNowe0y2JU4g4jpr5So
17P0/gQ+Tt1d9zOMb5l2Te6CQ0Ae6Rr7diK4kjdl6PzCSQEjmVwGZcWwh1wInn+I
O/YfuOEDmPKZtmxXvtDmCbx88Ysn4dQA57xR8BICiJoZpunDEiJ0Ny8e2XT69mU6
auQrbUODRmowaiR41K8RQS3EfUbUB6fp7gW896xjW18U7jF4vzzorpHLHpSopEO2
px5l9PfhxpYRATYy2TnvCiw8sZ9sLeqxYhfCL/9GrqdwNuoTmIWdegvaizduc551
Xp3ILpPVaKRCsncIeonhkQcwjgZbXYphDWQyFceOmLZkbO88D2gJySW6grzNwnV5
E0xHHfLq9MIvE1yy1vRXwyZ66IllsAmX8XmqwUcOG8+P1L0z3xwrXET72sD8In+n
Cuj33LbmPddnhpuhqciBsM7VRNd4HlMrrQUWJ3pEoCmLd/K5mmG6NPTZEzMzQsWn
`protect END_PROTECTED
