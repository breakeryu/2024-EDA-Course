`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkmPMzhQpS4tVRAdig8Q5XhZlGcOoyLVIW6O1+h9RAiZHLzhB7+hRjnIoE7gwoNa
pLJgmtAcbiUIgyC/K7p5dxS1y+r2XWWxNsQEDRjFThRF0dqguR3/SRlTyiUyycbt
ec00McmUXZx7SLbgK1b3pkgnjNbvm5RukBrqMCZDFXyMC5Prx3aKOa9b0jWSBkLZ
xp0bzNzfINqgr7x5YCb80IZpxNg4V1yTB1ktGzJhdE/5HJqpWp66oT22s728CWz1
4Qf/DYlNAMTqsvsllMvgRgobvrZM0OBsotCdpMCevCk/GK0jEvf1nuU36iYRd4P1
f+gOOrSb/cRyw/HWFBPJoz65t7tElOO1ljJ3xzDQeg0nIXflamTZptzXkmFROcrM
GQ+bkCH4qqBKz2rIVNg2ad1igvh7aX555Ka1dNSFc5w0H8j7BX6BxYIcHLgWOYvo
yFrFv+wrLaPF2zjmYyQ1+XSuQcqVRialltMyv4ayR1TheivY10v45hFWaLEpsqv8
8+ZzEeYsVJdA+NDdoFSj6yGbpnnjhMFvIqx2P1IZgy7zsM/crEOMmVoaWMqGk/ZH
5VGFh5xyvzzvGmT+ZPJro54tpxOkZVx4hLV8/mnqCWIp1/ibnBG6zj85LjykWMT0
kqjeiED0UODYmVv7oeCnUVsweBsjcfOYjgn5dg70K8ua9S1lfWb5PSwdu/E31r1V
m5Ij1O0hjgboBQ9r3MFdTc22CJULRv4GWh4J0k89NXDz5BbB+nQn5bPdlmvOjGL1
rlwlVSsP4ALIVQM9MQ3o+0AZLw3HSKaP4YoIZsXoz0XUTBNGJ+sqazaHI16cQQ1U
myu96LxaPQISJSGpnQNg3W1Hr6YtYc/SDdqTveZysbemjRx6AIP/nVIlWK3fdh6x
t2h5XNdpb3UAHqeTzqeE25OO/yCOnVjFIi6mdSREqoH89l8xY/Bst9UU9pbXp5xa
/yVcflOGmZhmwH5+rMtp9n4fx8qKqqL/Nvku1o9/rPnNVp8dDNz+VZTezCnSLWd5
hELYMTpmCwSzEID9sbfw1HqGGFfsg+LzNBtBjRz+wrdalDiZ8iagHqdYk2H+3cE5
B5ELLI1OAnOt0W7afDLEsPb3ieCxAbAvASvvJ37lJn1ZjP1TlixYSzsKF/vc6jAs
tO4eE7uoIul9nzY/a5O84Uj92Q9kbxx2rBWdIRtheyhuv57RY+pmdsPlKuc27ZRs
/Wt0Ih05Qb2QFIjRc9z9r0bvVVJv425kedrpnGJcbRXKkvqoFi82Z1WyAAc1j2hY
Ev2HbPSJ5ZpR+4xRCrQLC5fwT4WIZImg9TialIbl3ThbcjGgw6ehpb8Szn/c3uah
f1DMHfdD5lUO6pNgY4PzKcs2SZnC/sUDo4CVmwskrr3WlQW1aUaRknKyvBJXZBMv
tEtMBFdnjX7XU5eaDYDlX9COG1+3Gm+7CqcDtImBygn+e6zz8sb/ra7rlCmIoDWK
CkMd2Z24gBd7Fic2qo5zo6v7sHuEZL9Bc4j05RBkuCgCxLs0UslXNJcz/WZ6NQpy
jtvU4xOELwSCsSPuLHzVDGtmd1i0RzdRuWZ8jQ3uDj5SC1E5uuHXj0aVyrbnU444
Xdm3DUa5WbthObVsjXh/7WSLZFaJ9otjq56w1kMUOhF0nBmP7kU2Taepl6GGR+85
pm/pTHdyhk1e5TH8mlLnOLxpW5kehgxdSvupXz1xu77d3ebHSYb4CxN6ApjuKT6a
hMjwsrPVrsIjevzFvnShPyAxtiGMdnUCJc01zSUTrgJiLJow+UAi6woUM420t5Ap
AF6BfMeGR+H8/CjA4kfOpuW+yS11Mvll6EZrSxuWUBbBDoWMgRSdUhb4JD98BtBf
LYXDFxUFkmM7lv/faDq9Jfs2rfghIJDXcMKXYTfQlbp+GNk6DOv+lsn0+XSMueRe
UhVCb0yV+T3lOY4VV73mlkkXtHNhjS3pjlQFdCKfcVJas4RpuIUbtF+kJVrnOeaZ
eg3aB7Orti7s9TUvKSl820s76hYUOlYT+YRZ3O3yf1H7JtgwfjvqaL6YC1VmVZUG
9mJs0qM6o3Vpc1EWMK+oE0Wzjpa4HNdFgLxqB1RYz8LHmAq5ts8f4L78E1gylVXl
6wOLVu4/z43R5GsP102iEu3sLbYZN3WVeTUQmv0/pb4M0Yi1kaXqMZsqrr4lud6W
5lz1CuiykGRST92AwRsEALSrLoSg8/HRFJS7a/teRePba/VtN/xQSBU9HRooiPhF
OK/bS2lDDZaoxC3QH/HWMO303+oV5s2W4ip7rU9SK8wLzUH0rNgdMlq+qcxxnsHA
gesVmSxOWYscY+Qxm7175MaGrV5P09efCFCNNEJPAIjDdJM/6Uu2e0IuclsYdF8f
tXds8J0VYCjBE0b6mriQzAx5Tm9Ypn5WZNsrdzYI1E25O+PXYhZUuzka2GnV0UYJ
BVOz6eEtA6TfjrWp8ymewgB3ieTuGcUGtGMrTox2u0PCT7zNvFgvciGfTezJwXqm
q/i6OjDvhEoQWUd0VoW+Y99refQhZHmyh+pTXIU7hhjQCvTDiSuvWe/oyeC499me
tMwhJ+v0bysLin8moSsGO254MvrbC/d/IHIQYsAUlawTd0qIr6hclYWVyHw7pliJ
orYL09tpR2w3YfhzCGdRD0fFfgRsHrsk2NTD8zeP5JJWq1L/Qi/fHOVbUII70s9+
BnKicjgVkA0gU55pxhPrf5kBAMrDlR63P1Kwfnkx4TeM+NyaKUUitmC4MUKa+GpN
d6HKNytTxCfkBZd9OEuxlE8M3Fco8vZizrKxFceEojlusZ1JCpRdZAhjF+4f6GnN
TAXY2a1As7gRUYYAQlfdz2smutxvAsJyuGYLBsk9OedGMKY5G1VuzLMEx3J6a6ar
atz8bAexkDRhRJZHgITxctKIaHoKGfoW89O2/gG6oVKkYt9KYcE5z0isa9+YQTQf
x91A9tSx1fKBww1nC4FwqHOzTkayN/UdAg2jongplW1SoOE5uvnTetzI9ozLpmE7
GRdEbj/7I4fkBIc5jpfIGPienzX0cTDGtIbTDi41293f9r5uyt8tNBm5Vybv+Ho0
gNKy5GTjmY5+bPdk0NiIotQEE+zuKp2kQ7XGE56KH755UmlB9BAPoe4q7tzLQRkR
OxA8jjc6cfHU1kY4tIeXpDlA3ZK13qlNG5eNzDI92cqKGNpwfw3KbYx1Shk2yhsW
fQQ0xxiCQQJ59DGiftyp3+H31C84dKf1M+Fs9I0tX45WkWEqebZq2o8SJb+9CPTv
ABKOb5YhjJsuXTAKUe0+ELJpP8OCaH8nMpYvePdruaIZy+pAvJcNOUloAO8sKxs+
71YChGR3hkbNT291RLZm8bbGeM+vlpEYKKLVriyfo71GtnMQ3Xt8NXWf+mZPBGjm
Y/kabyAOecms3SK1dMGjiq8GteWBAgtPkCFyPd5vKa8pn3PiJsyN7FZnfCVV1V1w
WvPSH097st65h+8qceThq0G1PYcQoJtEuitnPc+i/HZgC2+mpwmV80ACBNdP1z5Y
kCN3VuT2Kb2dxsdx9dsVo5tpQC8Evkcmr+gOWL4sND+Acmmm4jg8JQ6mQKbpfqwc
zxAb58AYKK1Df4+oDeQ1rwBvUFGJREuPvlDBL7X6slZ5axSR+9b9TNRDKCjbNknw
3rycPmK6MGHHxy1iLr8q+xxZzL79xQDVVrTuoOXOQE38OdgglnqP4n1famQn+N9C
ALFk8IBXNYCJDIfa77lg3beetHC1jWazbmH4pNcNrm9nFKHdbWx/AS7R0HdWLZDd
rDOQ0Q4f40g+Ju7Esitu0qczk5k53K/SiGG2KJ5/TZRqPODOOhPWSUbkyFp1keCw
HN4s7W9a06g7BZAd37Am5O3iUIFy+iaB8i6jM/XA5DT/EgfeS8etLBcOI90G35KK
GZ3RjxXPN140RI/NnUPJHUnp21sPiPgtmXXN8ES0KLxVKB8NltPiVgN3lV3fl/xT
JdWv5pYSJAxD0skUaIzp+DlNMVbc7ppJv7gBkOKLBihkbmPS6TBQGvMwopK/ST7d
rO1vz2P+Gst/NuBwzQ/os8r0qMFq//WGmc08ey4A8nwHU6sx7GfBYvnBM/vCnw34
ZTGd/XVWADGY0s0moEsLklSzIobGo9/58mEPW3Q5pQ8QTgmyTvnJFbdiLSbhu5Dn
Rq6Nkb3cdQ8bo6Zus2PCMR3Jy9DPLzpaIWoYQcc1fUiPgs56anZdu+pLI0/j3Sce
MbJ1Uou7XtqfbE+8OGe/f+mZ10HcxPr18UoS59pP59hXigYHOM7n44sRbXJMYPvp
OQXpy21AakRiZS1vMM1E5pnZFTuvS8m8/3zkv3HMp9oL9UPLyObUKF2W1xgeQPks
oQtdHNORfaKQJC78q5wAR84tph4bbQf7jQi0sH/aavrNCKgpjfaBGnwEGoNYVJiC
7d8FMOzM6zSIZp1uuA6HWNw/xBC5WW1gNnU4DngWUpB0i03ECRTg5xQjWMnLH5GK
NDaYBXB0sBQt2a7g8IhPT1ARt+MPHKnj1bRK2iF14kyLcv2MB7nyu3Ev6f2vUlpL
Fo2TKF4bl5lJZdwbvwlA7aJnjfxjU9DX3GBzTjRWsWMf0V8CrXDFdZ53KcKqOIdw
A1PHwX0woZY53PA+ulBtpr7JpAUUmnKOZFF1oMoHvkmOK5VuNb7fzJmkmjr8AbxL
dFnNG3NokgXXB80M2IJgOay79FPlhEap6t5Ts8zc5vCV3QfIQKvCzJKWLpilQ9xB
hKRuGxuLYWinqLgB7p0AcnBsWJyNiBUmUXkBnTxx+bx6M7DPH4cvaHcmx0HAGTCM
nCyYgGWtRsy4GRIFfa641YEUZ25o11SEmDtMfdXEe6P3ZGG0fSLcOEQiAJxvnLbi
Xnn+/lXc03GsLAWNxFlh4Fb/rSthf5ER3JBSyFfda2CRblZXN5Gf3qaKwCGc8wcF
KdJIgqBlWNBGib4SY8YXzmjGgcQu649djnhsALZq3n+6eMgPkteJIO7hIIw4SCFz
Bhq0OojU/kYda0eUD1xxEb6Ugf8l9q2SYvNNJ+CSxriVGf3G3K6jYqIoYkjQhsoS
yDfTNMy089/hoC/QcEgpqji7WlN0q9u5b8S0ftJ+nhN8jtybbXqQJKJ3C6qNZSpu
iMIs8ZkuIlFGZBCPMhfLODvxs3hzVz6UZkeXGFEYMklRB59rDisOkzJ5hyPkqpQX
5bSM/JyexWWaVdQk1C2AKC+H/EzPAfhengQpOCsCsE17b51af1Ww6K5NE8pKf6cM
HPw2bikj3umH71caIOLaQRtC4taN3oW+w3T+ucHnqIrJin88ei1QB7WsTd9ay38c
t6fzMuhTFCZav1V9QwAHEvXCg4G5daSoLh9n+z+K775eGgQ+2n2gTf3Lg7us42NI
6b62uUpA5d3Abfg0kVjyIrF5277HfAk6LL80V057fkkiGuxISqDD/zlgZXVIpH3e
9HZFFmr/TCk19xm+psPyHCwCIJok2lthZbcd1GO1jIQwRtY0Ihd9QAEaw3BxCW34
Ib1GClmAdLaMEHlqzqY7jrT02lAYuALrrWAFuF1vmQ7TuRucQeuX6K/aw8hDkpA6
OAP7OOP6j+/5nMhXlO/FLv8nflKKXSuwgQ3saBu0CNytFXS+U+9G1YV1+RS1vVNo
4/Zrt82K+kbwVmjzTMa+WyvLaWvGM2IfY6SDJKZfUV9UEesni9whD2hNedvAGfzZ
eiZ93xVwUzQhXsYd5eV1NYdxVvZC6k2o8LOZgNQ70obCAOihvo1Vlg+ocq/DUwgo
D1Diy0hQYZ7WLLa75lUTZTkEjiXJWK58A3dwjQL/wlagpQB7OGfx9TN/yCVk3a7n
r38ITzBmJonsDy9F9iyuuVvDGtvujPPZsu90WsIfG2JcOjy6eXy48c+ogyOtVBD4
/hxIGPS7NPa7aRfJnAPxRcWkVsYaEgzLxO54i1ZqSaJ3NuxF6/sORypr415ARHEp
Uh7VBnlvlvyhHoZELccrNN9QV1nrxVaoehKyyN/APWVWH9HN/qCJTOModwFqhauV
cT9w/evFoDKiL6MRmWEsR3d4NDvqSJhoKX8+OqCkKAUs4c20+si1TU8LbBDNFEMB
M4QkyLSI+NeR+UK2vzoBRsQJNBlHsOPj/dMJZcwp6M4etV7ioP6UhSDGdYGVnCcH
AGP+rI3IgbYpJe59zYUvKLBvnL65OHlmIUJlnJEKA221CsZPTfWk6wxkTHYLc8/r
h4xN3cTJpLDWCpgTVPQdVgYIxIWYPYhiSqYe5VJu+5Mnr0TNvQsFNv1R1dRwQrhZ
tH+KceZnYKJ+wiOIbjNk5qRD/PVRKTuSXFH1Z505d9O4IGC9IhYq3FgwpbGL+Sv1
LMIdO1KDhD1FirpOLOADQ7N7pVIQ+Hpsci/agRgLaZ4AuJ1T2v6SUcl1v9gybmhi
4NWWAtcGyY3Vm+igVs29ei0CN8nnrozmGVnOyCQhAGPfr1iAqsMVvnu2e7U5AHA6
L3kefpYZ34HCrZawC8Xtgi4Wj1BpOmbeYzAdp9KDw/RbLvxz4NUwg7Eb3EbOAZUK
qE00WRi4Lm48eSdy+5X9QXG1keD8K7N3WMdpMsIt9awsJGd8yJIU4ZTTjy4S7y6f
Q7tnCR6oDnRN36xpFtbJSF/i20el0EZPQXbmBDK5YLNX1My8DRGdExcMS6B87ykK
MMQ5PvoFAmx2k3KKMBfFxubGHASwYgK4G9KKq9RD/ahgLdw6BmDAJtWHFzSrwOaT
3WiLtQ7uY4IuA20ruKgkl6vM20ibTlpESrCY9SHRJ2z89Rb9lzpN6zn+rLXHDCyA
10FuW5y/wEZd/z1q2g4A/cPfQ6qR+LG7HIvsvd3HXWfKVdOXkyxLYPwsW1gMz+ie
wAkyw9hRuKfw5YNipYwaegdqhRocV0CWSTKaHsNfHfo5LtdsteXlJkjG4N9mZjAh
b8AfBZp7aW7iyraiEOcXDC7fwi2VwysRHff346x/GHy951b5dmE61mI3f6gUZghM
Qmng+WYtOgZThVl567EF+rpttZJxknI/2NUyEYefrI5F0mFC7E/Z5eXdF6O/SHX+
Myc+1++Npgtsg9K4yOOpnnupOlUQ2fpEdfc7Duk25opy7Nryeii+XRL99Zuu9N9h
4vm+dIVnREzEh7ldofuyARyIX2Rfmy+Ut1Ps1eCqcLA4EjpcpjKyH6ok85Ew6dk7
3fbTzUvTwxitO/yzP0Lr3ukEFbuqq+4dAsD1timtVBA1rD7l5dKRaz0jmQgYw5dw
XVyDQoblnjBPgruzxVUVeOmPAHsYf8TrLpUc17iz/FSo1jVAwwLj8WmzyXSBeKBN
/eVkpoueFVNVuinVuThCIpq/dRtYSMdMAVBDHX7kapuhwMQXoplrf98UziPmrRYP
LBP0qUOUdfnUxmLiflUjRTJuWCQaaUgVcZVU/ZnBQeOfRTc4mnjjECrAnJK61dgm
3wAWPhh2xDCoTHfEhvak/Z6UthEetZ+dqnTiOuKEvv+qdJhozqEt1gcPIU3orDvU
gpqNTCst3dTG/YKV7n7T3PDeg4ZmDeD2UTgSKY29BDndBcQ77IYeBWz5IDnie9zK
tJ0KTbPpqOQ378F4GKNz/1lHHGgr5MtWp9DM/LFc1rZo9pqxvqp9f7p2h3fafeIC
/xbPf0yYX8Bfy2wFHbrgt93VQwRKfAIrjOk82U3e0gyteiA5DVaQU5MLMFB2U/GZ
rO8sUavCH/i60julAWPhJTK73L7ieRH3TXjO0vedSzxflciamWfFYxYpVxRsu9DX
JIjA8c9nNeCLZYVGeC1VKdQN6Hj2h9VRH0VDcbOQgySUO6ofUWhRD/Xac7y333Qq
zjTouzUxRckiKn7XQ7YGp9FPAbBgBWc7mtz1foU2fkAkxsoXEZnd5WvaQ+Ra6txv
T0wt4MwCB1ndgYZ/gREJYjTo83Z8kaGYJcTuRRNiwHkVrpoU6FL880AOWk6OG7e6
5XSSrF+Bsv/TKVmT6WSiDtS8OIooA+OIJsu6RUDuw96skdHpcPG7lwR6ASZbDYCr
MmLJJoRiDNRVK1BPRXtRixaRmQfCHzNGikBkBRL1ZOaehjq0iG4z1sZBIGsNbv9S
thqgH8dyIdQ9lX3wVTq4jV0gTb+IPuZhMhpEfbr19kmQW/G40w1Xwusy6hNJVwTo
G2th4hXqwqGBqZXiPt6Ilf/C+r2LEsVlAQAmLRlGE4Z5VRLc4hXRp23UONssHZPF
x2NgecSg/8me4HeWzdg78iubNcGaGUTYmkbbXJKe7cxkLmfB8zLnpfSVFt6PipKT
QfQ6dmsYyjVsL29fksZkAG+MeEQ5zs++CjUNcnFxw9JfIbLr+9HW4hvhG+inCdLh
9fTpw7Cq0gohjfIqgzNU0v4+7MMzKykhKVCrzcc2SCW2j89DDq/c7jTTD63OgbcH
Hx4olbCA8xjzdQfb8VvFAPSbdYvTynZgUPOVfmL9HzQXIQy59fdfmL+xBJtT3I3p
4k2uCGhp8EMH+ayPMYwOL4UQAYaRe+icXWlF/tzG7rtU8pRXpBSF3VRf5p0RxTAD
DgnSUughtS/Zb6Fcn11LBfHNdjq/moil+LH7V2AAFVIZC2uUD4OguXrdLH4PjUjg
vJctUOqJe1Ki0E/ClVHyrjsVKCIFrTlrYU/8e9ia1dfPkLxXM1XNY7wC2GaURCmv
IHvtqr3IyRwviMFKyCkglQvO4dqGc2MxkHAk6Du87HeDakfLs0W9XOC6oFVq1OHR
hPn1Sjx3jWUpR0Vx31rFyb5F42VSaZxeYAoUxcTcneT0kI1jfkWzx0Ff2VeHE7Ya
6lXsxvychxjKtaQa9oQfJYheUx3YQ4sd5FLMJyRK5c6NvAr388R6dN/6EnRIK/Bd
Xxwv0Kz7MOQfAOnfgWUMbGqRV505NIO6ATFQL6IYxNoDn4E4dDdDN0f8EDKCtQFo
7klo3nRY50sy3pRgBclMW3Ils/i3iTzW1vvSH3KYqPPy5FnzFo4j7uIsTbZVOeUr
zb3t8/910IKxd6TJTHoz9Sbp6qHgCDSBrWr4OKzN4eqpYBSfHqvV7kE1uNu44ePH
D+bUrZBrnXA6p9+7M7KRHCU9lEiH59nAncsrNpfpFdmOlBczWk5esQq2Xtycu+ss
+1yas0tP5pIREJTPlBsT9MYHw7EHbdvmllnL/Tc47K39QU1q+PPDJK0ZUCdVcoIV
XsDnnpMHbWLl6zNj+4CVj3NEtnd3Lc209b1TB6ZnH48UD/9Gf32CieAyt9Nl2+d/
T5FfbsHl5dKUfN6O0VufKLMaUwJBc7oYne2ANAvCT0bOm4zQZaIdxeC1zsh/N6az
UwNCDgqIRzAgRUbK+bW9Lw0oPvsDNqXVsPjHQ/tALP/uzLhj4nOzzoUZMPssqSNV
3u5P4jRRiDLxMe5M2Oy9ZIkJHVBtXyb4wGtYIvqrzaIbOJizAdC6nd5kL4bjy1Py
zSrT+bvEK9vbY61sJlQPw7U8tQD8jLgJ1UnkX1V4FMzM07y7Fnm1mr5iMuGAtByl
yCQATFTesM7HNFj4WXPHswPEgs0oGRe+z2tZhri1w7mmZoss7Su5vyKQlirZf3r7
MoIS22OqgEDIgGZvEAphWqLbiWA9vTOT/E3OF4YRPr6G12pPIonyJzJ6kiNDznAo
THJONe7US/nxCqqCmh8+bjy+4Bv0pAe3nZyWBtTUShzfGdNWWz4G46NCvxefRDqv
r1NkNR8QR4xxRU9mIoyZU2WMggs6jdStx+MiHkdgMBLXBR0O9m4YSr4HSCuv5p2S
u8xVuphA/00cp8uejgxYIxS4NY8jXTsKC6huDEPo+fmY29FFGCwVsu9lsfQx+oEW
v+hX+C6DqiFrr9AVGDPu1CitFMYIuwgFttjXFsOf8LCjzmw7IScDW14eZ3fDFsnm
VWMaSG0i9gqb77Rib1xWjaV8VuT8ePuJUhBfGn2YWwlzIR7eYu1iUO4dGeRQstpH
3RQ7wGTssQ62f4KTbVp8tne6X4aGjxvGGWv7wCafsvkqc41HCKpdJB6tdAVGyyUH
7Ht/p1l+0ZHaEgG/G7/xTPiT+b5JRUFUCR25eNgX+h4tLmg9i7D9iuJT44CRZ+KE
h4jLQdLsD1ZvvKV3PD93fmjCFXH6CXZw01fyB7h9d/XL0Hei18JCKiOJad9MB/FN
W1eaSsSYsdVNn2EwD6EAADm6pbhJg0eZFCILcQ+dc0hB6reL/XyfgWD4EobhW26H
jeeWDbFkWchVMRT62eLgwtDIQdVcqwXgxT3aDoKVbO5z5e9j10T30jBIfCCly4p0
ZE5SVYrrnz3tYXCwsJYtc2wUJon1idFdN2yvtSPO1RC8hUYFcP9BjOZzdHJ6CkjQ
zYoGVVIBq1BjO418SDm9qQAhhbIQym7aEtV3u0X+DH0eEkI8s0lODXFOggMGxzNU
fajZzHmqeR3ZFX9GQe53KIK0+skg7om8yE7RSU9cK7mKyaxVc4T1wqyvHENHBx6x
jPA1HSZPw2r4L+O4igVwzV0Q+X1QV6GOmiGFqLOEBvM/0iOwnTG1s9wCAf5AVX1x
milNwphXyD4ZsvgbV/JjycW9PCt0wj/ER/SxEqyxT33PXUEb5wJBkwduWBNblYZF
XTc13qW1GSpZROYgTaDiJ2xY49/zt2mJLGkG//7vWAmS9qoGGG3GqMfobuYzGNW+
1k5PkUFNhMsX5sbaLQ7rG8291Fp4Q3Q6lvl/bpPHPlwodagGs0jOXm7DtHo55dFq
NurQU5jjENkiTHRrl+v9782O66LK1MtCQka37ZMTBot6JfD5eQR+xUuxhOYSKbbX
BvtHzCZ/IICsQh7iBjcA1wlweHYnNLh7itqgialV92gaIMLFOOjCL75MLWr4TeFp
V8lFEl98AeSPTa5AogxS10qTpvgWdLlkS0lAEnpGGzBpmU+J1PL1M7b1km3cS+Fl
VPjrcMJhmIpEo+MI3YN5mQAmPPurQkhoqt8m0YDEW/tBTSJr8tDmGhF2DAxacseZ
xzkLqYw4oeLCwWUotyAGmg8fjxvGO5Iupiu16YZ4peVLJSrIXL0R5QGBFPsG72CQ
FmEuYxc4om34AHacJTyRZJcLfqEmh4LXIy+/TOpnUBZSCwQx3DdtDNzLmwyRCfUS
w6IRDM+KVd5BFsx7+T9lxAMgMPrpSfh/Vf6pkRBHrAf2EeJHNUwOHjZYHw1J3riV
FZR2Z9nAFXZ1TNja0P4/1IxKWbsYkNPingXS6Bc0emkm0WQRVhR3UQpqbES6Jms4
h+HCa5x29sW9tszrr2bU1NKXUkiwcKXN5M+RARCy/RTCZueCi5hWqLCBq8zKlnOP
UQvkDDDkumfSVcP7/lFqIkz7e1vMiS8E1gfJ44HwLc9MRAj/glYpP73YUzNc0j1O
U0jmbImqxLXoIXKSNzeEIak4yYaDP4XrhIt2kEW5NUf7bOOlqtZG75yc3Z1P/ftW
FGUmfkprLlnHRB0vdr07U3o4GOY/yR3lW3YHl2wylUoN980Y6vIz5P1f4bw5fQJ7
pfEGlVEkTsZBrwpgdtz2ce0foV4S/TK+DK2FchJvmMjVdmm61q0YU/6yPRRoTygR
JkzIYYvkAoEsKQY7MDmVxifz6n4C9djqGDzXKZsHDqxPhVnWVcv67LgEpK3nVX+M
o8ZNeAOcB5t54cgRG+uB24rsArKYGZiaTy911WCv5Xa8yWqKWSiNsqv3CU3XW4D3
UJughqNHVg/4vlnesR0/LlkT6edP8PL4iYJssEMFtNg7nTfAYkbtUW7J1Is557m9
hIDms8x4xGoYDv91rM8oTUWnIAOCwQ3Cy2g2MP7IU7ufsWXXioJzZF/tuKfDxvPL
ZRYMJyU8twtQskd+J9NHPppGlGYoOR4TFHw/aVr7vbu6eFhN96MzxMQpb4IcA145
inVYdw/qMJYLkFWbVnNp+fE0c12FCVwrelVaiaOI10m85NdExK6lFxoOJRJfvs7L
VVRCzfsKkabo0Ozuc0x5Wn9/L4pI4bf8pWDpDAXAjfUvjamMuWbL1jF+EguiCMSK
XYQF1HxyuNE9X8kYkYM5+K2J4S25WUsay6EabR3hVirSP/P9XGamXFPK07dxi8dg
7BziYF+FDe+3yQUc9Yy/sj7Y1l4H2C0mxe6vZ3L4pqq3jxpRvu9Vx5FwImEu65L0
EIAY5gSaKmdqagYwfd8aG0JU5NpHiQwH2MF1CvvmhPsEfRiWISwvv/+yt4qYkKx0
xduaklDfPd6kzphmrp58Q5A42Y6ORg8EjOKA75uDPMVx7ywooMfhfTdeuEdtFjOh
QpC0LhKt3ts4Ujk56FaIr62n9tmgJdQoA+9npnnH3u9iq8pqiVovBmwpDLt9yuhR
IdRTcqWRqZnHz/lH/wpf3Q1x4OyglZ4ndn35pdG5z8MdDCjI7kA0edgtSwRPZ9B6
jj2I4atfCmLGuW9+Ipl1qydNUNEU9XYSnT74R6WAv4MoC7zRHHjUb2Vob5LbTfHX
ERncZksVI/yWA/5tykjFv07PlWHzfrbTlegfceNGre+hnq/CwMHLv32XPMDVBQE+
XEpRdqgM3GzkCdJmNTL2RUYoGe7dDJRH6IAainUBznimPhaEWbtGAUcP6CcKMGPt
QrTT6la0z/9NxhelDVfryoOdWoPqyL8Qkiy4/eT3DHV11RqVcc3mFIkdeKlzI8n4
LUlOze0TNgBr+TDL6RvrGbrSrzqzKNIVDB0jIqV8lufpTyMIuNUzBCOH3RQEFjme
7Wt5j+C/XW7mXvW1+sQ49XvWp5Ry8K5Ul6tX+21EYPYGLV7TcO7HbWQc7xM++9CU
neQT3akb+KGSPsBcq3IzOMga66wYJNYyGX71SpftQfdCy/zcwWRrM0CN8ts/Y3ve
DBrembkQjq8PP0vNOcZgpPDwAdLZOOioh06GMaruQl9HDrMfXpTex1tv3Nt0bikh
M7++KeEalJbq5rcnue8MvqyotmSahwdETgHlfhRtjmi/H/KXCZuJ3iUDZqJy6key
c0IKFS3O57XXiTiIq9BdoDtwvSY/EtZHvh/cZ9zBMfM9tXjuiIQKlIqiK8J0rnbO
rn9UOLEABf+3781fqC8PaYeE5Xqsr4WJLWKrYMs5WAM/L0Pt92RwNN7sF+KfPHkt
u7lT0aRKp8kxAf4xEd7Groec7zkE1A2mOm+Qs3ml67+CROUnlQvlXbxSDL3d3Jtn
08M+d5a6KuGdP2NJRG6uorxoTR09grG6m36FcA75l0u/eumlJp+1NeHzipAAu07W
rnIE3cyHvBvJKuG1NRcvc5SfbxoUa/Q/dF/CCKvyqPK/31E8h95f+aa6AnAplEgh
aqizB5aQ+NH76ZewK93aCYQ2+tYuBKJNi+lrs7Sou719ad7r8ofr//x3InCPX/BO
oEpi01lMOZ9ls5k684ijbuZNzS+WIvLyHRje9NWxib5O0Rcd+erItUMCsg5M96qw
KGDhSHR+2mqIoG4LTxIWjpLYd/xv7+tw4y5uL3pYN7LR1Nha/BQtYPxmhrmn75Uz
TqB+AdSEgcwpr2Ryozpi0fO8KsBmyu8G1xRm7bNw2T730OgrhG9+/cguefP3lA2v
Q3SqyI1fW/asM46JKpn4O3xm43S0MtpXHQISJR443sPMLj3HZC8NTUpnqJ8Ifxsi
GUZs8fhS4cJ9wbHDgJUa0xGjLMZeNdFhp52lvBlYSnzGRsQyaJ+5ZGomZlKu2I6I
MEDbGXyYPPjTY2sEQCvWH0PkTnnwZJB6H2bmy2A6grmOkghnT0lCDhB7ufDkG2TU
QadaMMMyxe4sUp9z9SyrKsAY5RMifxlhRiAKuScquR4e4D2Z/odV6LZbgpkwZipl
lg/4qgjvYCBS0WNgVuWoOErNRPMUryY/TC6tkk1QsCXnIp6IBsBaVMp7dyAbwYhC
9wA5bwaTDmvtzYWuvJD45iyLb2KW76kzzlvGiP20ASc0FPzuAE5zEdYXriCuqdgs
4xC+eGW1BhRZsOK3NTSHmpUfntVsIvtsrVWQz+Kr9CzPer0xg6zR7tzHejaKnJBn
RGukUhE3qc4FUD6bJ+QN6pyVvGGKx2Pug1rFoQJRoCREpECElV1wCjaFQJxJD2o8
JwEpJsMqEGClNbOOLhrJLK/5bO5AzwPNqmH92tq95zRArlJoRXm6AOtda11+xrAM
w15G/1LhSadoNurQ93wdvVM8Ljdy41AxJQDYK4fqsWz6mcKmff/Ogt1vbHc2kIpt
0dbFnj/8g3urhXpzFj4lQFqzxwI0GXJSMsqTBDymrUvRDtx4YonrLsQujzsg1ZV9
qAdGgptX65RVOaqst5q4CcnsPWQEJ/iVb3axbmF9FKsLOhpGN13hZrRiDaZ8++ch
OomUN5B4u/BLIx+FbJdctak6m7aIl/5tEyIXxx8H3GTvS923HAe/79l1TQk6Hq7Y
C46U42MIgUAv7PuESR/BGu9uWohEddHV+GgqakprXF5mYSPdcaxeZdLtBLWIa2lw
REixKVlZRND7vTqMN8x9P7N2GGYS22zCpcjoENbXsdWUzRRqZmGz5mWLsKCgt9YT
NqYr28DY8ZV554konXLwI9wmwwh5ffdU+BssL7eOOug2Mg6/uJngUSIMXlHDEtUf
O8Yp2VkYbDaIWhfJPl2NPi5J2TIFZST9aOGEm71y/GA8V9+LUgDK6up93+3tcFpf
thETnhaTDJwHp3kr1qgd0Y9Yax6GtIslfj8o/UgYpgBIbi6sr4OsOK1IZ+UGlnu/
+M+9/NHnTTGeGiFSWhKe3DiktcsHhoTGIgG2TeFL9V5M7P24SUA86yEvq30yVwtc
sUwyjRtKMEOTW7tBN/xJumFLElzBowdZYFR1Q+nEXRBDpLqpc6GBPi20cCCZqrBR
MCRdkYBShByMEsWxZG7C7DOudjvEMYLhcdr9QlqjQ71Zv08GrLZvPwbxddziYpCG
Cvx0GCkw7FueJgeDn0+4tEkLEO+GQ9+vUG03Pth+RsSfyx/9U9bHvBsX1TNe3dcH
FiPPK3KB/ACDL5iQI5sIhxp1FIIZwLoSv3+7HMQ/fyEE2X7eNwjmKfCl56ZiJjtw
/Tf+13L4qBt+7hzNNTLZmBAi6fqXnVrzNFYEnS71mm3nTXTFzZQAdPRpAMjWd91h
Z027iHY4sDABLIX2BdlFE6/cT5a5RRZj0XyOymGbn8NNQL+2KZzoLn6xH7B6jvR3
IWF3tNs9JmfZYxFda2Jdcj/xLxegADRpwY0LBAZw5ZD3QBdR8BzeaRpCZLz+gNob
QqAd78HO3FGGUDJSv7nJioeltWFiRHmfFDa1nstI0SrqtZiDLeh4H/t3dL3z5dIr
ZX9gYA6TdIygMpHq5j4KatCfffejSDypiyPIwXckA1e9ohze4FOpbcf2Ziw+U4dx
Z3vjLfOFCyUdbB62Eum610Avwi8njJodas+AdIwp+rWVIPrmFjgf0XHbD6Wfn3uv
Ku4m4BtOjLPCLbdRuYBn+5A9VCL7OXVKaUZDVWArbBvOZKLGq69RnQ9+qHM3OSKa
mC5CLv2VpwBt3y8FBxxAQlAanMZOJxJ5ejNMTPcEEJPwCjWB8ux3T5ah0/ggyfTl
D4UmpbZHvXfxS1hOec4nwwbpHxLTD19z/hWVzf4ecC+bPyz7tbZN01/HfuCQr4JQ
ozNosXPij+PNCEmDlQdj2uDQgd+0ezBasU7uAyGXzEsNLPVam83Eft2vuE9nuPaI
8Czc/lKE7KIHz9ItAT3q4Wtxuh90xGPKX3Lfbyg55z4pnro3mIDLk7hBnxc4fJUy
KGgTKGLCK476BgI2mmAI78gjbA8iwE13WnnbNOM32awqzwenK17ofMtYvfnQwTSw
5tridKgbHqFEQFeBSvHnfW+gu5Iehg5Rw6NAEd+OgT1hzC6TKIqoFUOfH3LjbWD7
5lka5BdaAnMYwix7xfuyqbuaeGKj30i6fEM7hjmM/Q/Bewbfr5qPjtpB0//WBiys
k77CtUMARzSI9X/3K6QVXwuuN3++VjOnJZNMALciFBiJ4ydWkEcLI//dULdVmS07
uXljYjc/9HklwQUV/21nLk57V0Z+LSeLK/xcgh188BMYWINuGBKMug07kb7Oqp2o
6C0KcLf9MVKyqNkAIu1Adu6iMGgc0w2XLh2sxXk0XKftkp09X/+uDikuy3OY5pCd
cH9EmKv66TgTdLQcVfyt4XuDSlFNHaGGZA1HoRjAdBEvCdwzYo5XtHv4VKQrYmiN
NfDpO6xnTd1ZQ3qu6E3+C4zw1ZIfiNMwvqjfOL5wyAggQzrRPbNL3HnUZbnoSMOY
OyRExxRC9fFcR78blA17XDumM2cHUWL6fBS1+x9mmMYOMEbPvXi7L0uS+/BdTxv3
+47DOzNcqVKd4FaVQCUE+UjZWy7y3ZWX5ZrHtUuM6KBjAUR1zSG1bcGM71I6EbdG
/TNBIttmZxPRDnUdcdKlkxpfFg1qcEA8qfCnli55K1viOcJO9/bQlzdIeUidUbhA
AS5CUPkTWLlM7p0YNlOftnXYPp469xl76vd2XBRMzp/jNXvo900unrHXdXOKQ2Tm
X3PtUmAFw5FDNIupzF/HZMNndnrvu9Txoy9aDChVlNVw+sZ5KXx8hvcXcB/WWhgg
F3chvUuNENNbMlpOEeKy/cozRAcucs1pXm/xM51TZrY6Fa/fKNCR1rPgV6EaE9v2
fLBsZD41rYgfnK+bjoJs6vYQqotv0/KQOdNluiFt8NnLISXz6KIyY9NQQPH4HJXC
ShecCqh1+8J7rYY+K01E6uKIqnDEYbOVLEoFiHVbZoGOK/X+QPMHn9aWUOHBy+pK
4qxhBJFGeIJttDoAMB0pFiM6/3G0Z4Ah1zcaBdHqg8T4flzxR/DGOUqb7qKPrzx0
gAYp1gufZRfT57iNfuvSz1cjNkvWsbWqNFzo3WQCr2ZqJeuBhkLrxp91fwe6onp4
ovuAcn/CZ2RywsawNkz44kONwAQaTDKkZKKFGDUNHRHpUjLARYa0fsNFCvwwxB81
bO2yBXZLs/D6HOjiRb5YsL9UGqPvn70/q89NG6IlEcH7ttYgfQIr8le6CqZOvJYX
FtAIrecOTHHpIobJ1fFRvFq6v/QTxzuzDt7sNohRbwxMb0hC9Dwpd39hNB7Q+cfu
Oes0bgiJg1pFZRAFAAmtyS9WElqjGS5zeeigon2whZDDzSpBFnSuJ8JAnp2fjfmj
3FmKpo9txCRMX0Rfyh7d5dZ86zhFaz7RnhxgaAlJevjDr8Xsq6IQZa5rq2TbQ7re
e6U3typxN9UVs0CQe22i2OExPtZm09IFsD4GGgNwYP4hP8dEU/z+aZlHXVUuUSwO
AzUg7+UC5NUogA7WTdYpXttms/oz0knMMAwr78FweWW26tcCQFRVceSjOh022CcE
NquOOPzCCAAu6OP83v2BYsf7HQcQjVOFsBo/Ukl2xb2hvLU+wFYc5xXN2HQ6Ayxz
KT3O7dnHk/WfaCJyv0sGxXFUycZo2FW8/6E3mfkggeKgJHZ/LCsY6/TPSJsLti6p
KT3mufDEfp0CwrryIm3b5RYUBn0ZNNNPM2j8iXMyFOM1fES9m9DgeYiNlTJoMJ38
Pqfub3uGeigLcyLeHyWPAahZ5safhlOv6iZFg1XzjVBau+lFYaofDHB2OQZMVIWt
/iILMK6M2TKG2xKZ9ADePMKKtGtoPNeMmOZf1N16xytwwlehUD63X+j67z0d6OKg
0sVT+Jn/PrvmVflsLsvA1ODx6yiecG+ku5iGr4NMREW9ABUvOMCKZAMcSp9OcBYz
uCYd2MDtYvSuceRnwlIoa6nWnYDoBDJoHEkLSnLrWuS50pOWCGjqSI0aVU/KShGw
2bJuNuFnk65TONHgs8ZfMzaI5cNQLPnGcVxxKHegA9Ip55g00DTAEbN3TJCMCDXw
JQj6TdCLp6F0mmIk6dFZRddLYLMKi0EDwt7EoDmgtWZPdC+/Y6odnfiNQG6p8aHQ
LUmhew5wAGRxd298WIPLfDQlBq0DtB+Pj3QptYbDOuZ3hIA873qBVA17vny0eI0A
X79OMPYn7wORgf+OeHUq6yC2zadPxLtFRe3O6jgJ/VgJ3mZMxKCk5+kEPz6h9Rtb
K74+2NoBcNzXUZJfLjNGCwNPspc9b7l90s2G5m6OBGLejz99xyVkt3FRt4XvXXff
nlnfZ8ViTjNzG3Wr/1Q5A4Hw5jGM9gy5I/Sq05CJRtlN6dj2jj4EnmRtIUvHZMSC
0FA3FgMdVaJsUJmomT4614u6uH/zDYKHqZkToG8anFo4ntZTfj+1pdsbptaTc6iZ
rYL4xCQWnPP68wDhRwWxZra5Q99/LF3EAgA/6uMMvthCAiiVI7IhFECpr7sqviVA
PTpGTCkTIDbtPP9EIQL6w0ZacjrsX5uXwz9Qpa1bcZW22OvVKenbzqJ1rCKkGc4S
hohgO1adIGrDzbBoldgBMBN552QrtxdCxhcJkFb5mXSHaxMNa6qisc4YHwpVj9a+
k+EtQcebgJ45VZSUA9LNmnJrpXpdGOdaQIqOLiQ/a/uWulPY1/7b3hUnmbdxh0jc
Xefek2rgJogpFJx4AdY15xucf6jnECW6v99GTz6LiWXTMiX6H6j4i8cHQHXA2y52
m2OwQ+5swt7t5mFeZFezeXHTMZMX5r9lDdSZ3/oFSuLdzhjUuVSqhCRR3UwJ9ktv
FQvummn8CANmvXCZH8MsIGmsAxgjIpeAiRRjEO0JmYMS1oldkE6vg+ZHONisL7nQ
BzZJubFAgKUbDbwEkTaxRtPz/oWU2moL6aEdt/YI0vAv9aEUQ7/pFgj7IyMrTRu9
iBvjCTIWGt68nXwao7e7G+aNgrmy7j2Zjr7PW+GyE2kONauRNQ4wbxv/XmOrxv9i
p1vLmST61tYMiPz9Fo5VfWK4bjONxpwOcc4kAlhE+/fZRYWIeJvERVPFNLI15jOt
2+2YGfz0R1MXfNez55UpDaHVGh64GM5foZnA9z+JU3tWBQPgsQnZpOKvRU+iisEe
bNFoW7oobwrKU0qbcwav0VmS1AuwbUYtaVo7SCFUYhjZyLXo6JT6KBrIqqiUbfAq
nqPnR2Q4JjW9P8yMQ0BVEFx8tnJA8FMByHz3wLyn8uP9w9XJBT+7s80P7d26gxo0
vo28pjT/PtR6Kbj87HI6VEbO9cznFI8HDPVRUYXqUSmEcSsZg87D5qkSNuwD58Ge
HtnXZw/Xcqp5exgff8DhuKTomx3o/fpJLGaJ7Yi4oXP9ZE3tWIGP1u3Gdp2kESH6
EBMUKQCOH9bazVo9zVIe4GEeHVY93Aog81GmBTDzuTNe5VmL/ongVRqpVZvK4Wqf
JJBV7H6oc3dEvhOta0uTCSD+3Rf08S/AE7o8rYvvylb62ui1l4Je3FXQppb+bjAF
Z4y/uJpuVQmjwD5B9be9AwLN7YsPvTNQ45b1BexsCF1lx0dZ14sedVe2S2nqD9CS
c5NCkjgoROPLtByPw7ohXBo3VY5zc+LY5UGMN9//xQKBggGBV0EFPK6voTd6Eu9c
9w4Q5LiD7MKyBDR5znIpkVs8IqdvrarIHiR+ivP79nWIpnbCz3iVY55jHnt1qr2X
jDWMy1Sxqe0MNWSw23lSavYM3ds3W07bs555aUQeqDEv3G18pl3DbjOlKcdF2fVJ
jePKaiMtizc+J4S9+6Eyy33WxHHZm9yxj9HhTcohPHPkSCbaEzk0ujZ4Q11fuw0Z
bwqY/NuS+BivKQwW0IaY/1UkpVQrtVCVZGHPQdSC40glxSijD7vb7o7fX35yS/1A
rJPk9eJv5OrRkNh27NfbVLrznyLgazIsKo9UwJytQ47HsqTDsCNV9dgfSUqCXBNU
zxE2cerkEVmDYfdPWVPaOvSAl/FU9hPT3aI0+WSeERp78BGWOCeChmtawFi4UfzB
f4lCoYG0YqwTyDocAp51Uez1ZGuWlSgThMXCfA0Msn8AZvw5NOFYUKU+yALnGRQ9
5WOUxPmeGdhIIutmIf7sGQkDBlEhpQbijan3CR6jbNLjPOnScv97zoffTk4SbqaT
1wDxG7y4mkL12TySU2t/erTPOsNLM/qzoTprsZcBCcdRd4DK4Vny9UicDn5TZ1dG
3NtUsbwQVegScYsvVZYmiiCgl/aehdYAkZqiw0hSotiSygs1dt7sTl03NRIuBZER
+Qcf/U+mnm8dzjA0Lw4e47h4jhbKpWoEJvNaTjm7HZA5wQQptUJbzFe+3DS5+Jjl
VSafx0kpCjHucxh7JxqDxXpYzANxa6yV2GYjDw7xUqRNdcpFkH799lwXGRdUHSZV
hJgbSQaHn+aPfcc/EFc8X96Ht3+K5yRGIhOHRfsrEYdp+nRgj9rBAdzkCsrUtmRH
lc4iCYBzJ9Op/hkPFbfOJnuzyZtnV/vt3yWrcH4eTwDLv52zSOmmXtV05HLWCYLd
bF2Si+zUYEt6Sy50BqFLIfg4DJBOKdTOTmeiibop6ZIizYDRQwKgDFh0ho5u4CIu
mH0X4km18yZSr2InEWxslIjJhQNzGYn5Iov89jpq2iKy3cWfqJbY+ta1Gyw41nh1
nBNQNIpKedJkmcWUwhxmn0nEt5hQMFlUOq6ndBdM+u0RR0ptkvgc/cE9tiOUmXFt
CQAPJXPqkRqV/3LhgljhsoTijuhr+ewqe6xQHfiMFAvUmcdi02AKlKa0gYIVVJEs
E2JX2wykFRBe/E4QUndR+P+waPSY3kqRgP0XmHtpJax33gJ80X7Mx3ojobaAXHAi
CTbVMrvvWo2XkYI1DtRBa9qz7VPh6qFmTUObHCq4Zf1m13wm2Rl0bbdQu+wRvCBN
/eNnYd8WXpRCKTdbC2lLkBzzjIMUG+w0fwezHrmK76aKwnovfn3eD7VBjMN+ybcR
5HQGeXVfVJpy8+T5z+dB8DTlZ4IWbbGEzrQJO7t+BtKTb8kSd0Cr+eeF9LVHEdLJ
Qs4J7OyS3HR+qe0M8PX4Gb83daeZqWZMB4RXWMzHuJUFpt3Z29r2snR2eIA2Q2V4
qRf91MrXLHZ7b+agKKolWEHjkTZ8rZA2XsLQwHSlAqA8j8gwftvOjUaGomNYBSkB
CaT+sjUJyv7tzOFZbQscG4wNqbzEUG5lw97cGVLXTGEB7D04YYjVXBUCRQmpz8gT
TDPcVxeKXn/Ikf/L7h2UaWy7UU9haF3ro1J1juE95QyB5HnJ89s3no0fuEEXHP0v
Fgbtpy/vvQSWV9kdvAZbM3hDbH6KErY7JNlUxXtpHWIJg6jy0f+K7CL8KTNUFi7r
nAuSeJT7ibVC9+XJHq3Bq/ITC70UpH0NmHlQMvTAu82MpsgCwxLfl7iJSpR93Qcv
pnc5NoDjIdEWpkw5WjV5TOqruz+8lH7Az4SC4qC3MnMGttEdOBrGuO+DRWaO+9nu
t1bc4yS+9h0sU1cF8l5uNdocEWpWOHJ1vtwUNdPrPK1hHys7eqRfraty8PaQimZ8
EmBFa43Pfj9fqsngff3JHYSOpMpX184FMhEtUvoULaclGtlCpvC4Rd8jSYOWxRZE
imtq/RZofF6P5ekDT/OefSK4u3VMqCtLwL938HWyQwAylY1EI5LBY8Bv++fz3aDa
Oh8/l8ndDfwrMiKZ3Koxr/mxpCpQNrYtfe07UaiSUagfF0+2E7jZ7jXaowRxBSYM
R1VpWKasrkrSrAiZMmEIdd2/Sk3FtcmJ0aqW3eO2hImzLU7OMGYnZ1O2kpnYtROY
xOm5Yyo0AaaXtpaV+iSNRe2njrrsgpQN7PVVvOr0O80HZNl9bZaUzryTl/Qb1ef0
nwimPsmucdad8f6/znxVB5e82M6rkzJxaJ8MB7klMC5KxgV10IrgQ0D4OYAJRUxN
E8Hd48cldNe9QLvd4ASOXlE7nBdRA0/T2S6Jd9y+HH8OeUN0yijXnn3HSz4ZBhXq
LuV5ip4qGzXn6wzi3ltnCMCFA0u4dc7I2XXCJnurQ37CsRT3hq9QQjx4tgLL0kLK
4r01nx2Vk/5Hq9Ttto0jO0RIaZ3nCrWDxJ3TtRJq+VzvAX5hql7hJx1UrA1CrBsA
x+XrB6GwmYCS+fIVTMsw9RqcowJ706qwdyb5zXlyrwWGaIArMaI9YZ4xbZMopeJY
Eb7ZWUqBx5WmB6C0ZYR2hDWCXl9h1SO+1tfU0FuECqYIePRjZPaNt7jnzIiAQNyP
4pvBNBKzmnzvYqCEi7vA0zKhsd0o4xn1i/gahJE8h2ZBdFkyZ0I/HhrIG+wRbHlf
0dU3WA5MphdhUYoMJnMprhgr/sXM8/2GuzsMVGZw0Fds0Vg0/DVIal7reqcHm7bs
khnkVThytgh3nBwaHxsntPFaDh2Nn2gqySF13ec1ECqax5CibKwaX5K6dPSqB57J
s3ydATKuZnmTCcGQAE0o3VvrJW+8k4H8UarWPNRbM9YIWWDpObRRarWbAbwieGlt
/MV45+hMiROjpi06UpIZ5bTpy4OzVBtNP7c1u6XSm3j/VOgIV/Sy3gnjm6P8q3Ss
0GvFHim5dZEVyZ1hFpomGiraK0y6lUY1CG8YzyVQQiT0mPO2ouFelQsBVOvkhb1Z
Ael1laLnkvg4vQNy+EJcm7w/PwoNOH88sWc6ZkpHd6qfOAr0K5tqXZT5CfP8JY8T
2Ch4RGtsZbjXMEnHKq5OU4WR+31QnUEpEQ/ma+mwogs9bbK3xNBYD1TwjAdG1J0O
aAUCenyb7jK3vcO0ZkosylB2cJOb+CpsIjy3efZXPxC9Kt1L0pSe9iIjEkDrmEoi
wwFd7KHnz5FPUHqxs97Ve1/v6o8cbVJ7UmWvQsZwzE/YBpx5i5986L1Ibb3iWiAv
NRB2nTKX6PuDBsKVxjMj6C5B/Hw+YN0EfHo4+9D+svBy1IJfYU/BPpDiyP64i5Bn
2wCTgJ0654g9s/1xMBVgTO7Yq8hx2TDKAfqujBddLowmxcx56BmU5Rgy/GCNcNpy
/XHxbAZuZpbHly/eDruhpxUMZkQKGHBLntEyTdLZnUiFTsWVQWRQdfTECuk7aCA5
EGkFV517ZGPYgn0OTrHwzYqyDgND3lA0wUmmsB5BCKeld2zR8Gwj9JQi9BckJdZO
OCdSzyQwyNMiA53A+MUVkSvekjXvNWCIpJuVFIv0wYyHGtaiAeSqQNN7sTFImKkL
fSuAlhSW/y5ehBkYOdDBIw7lcjGQGxAvqg25bb/uiLZuebiTfRnSwQf6l5RKF00p
jVNCu/r7GbHqLlwl1Z5rorQIwF3Gq5r8lrhhonkGEAKH8T11bjKOJGa+x3HHZBXw
YcKRePjo0PnzThqjE7k80gst4kVC8SsDnoj0Vx+nyjHoD0X6cCivhuN69fWWInap
LPYpqotL6oYYqu7kLUmLm5BHZYNrwyoCc7/AeT8hA+U2FMTZ82sahARMgoDkCRh5
xpJxZc8Zf800uRrShATU5khMz8GIsSwC/plr+G8mkIQ69jTppj05/4Bkfh3lJq3t
BeBPmY8KYrrmfWtAl0WTZTAkxL1bWqRRuzASh4axjb6z5+ROc/NmmWcjyQJcrkXt
QZamsVEM1+lvlQoESf8bMydjJXDERZJ2aiLzrvapGlHpT3FRt3N6ubVmDDNfUUzc
H0BDLn/W/iB5XQe4fJOu7boRXQ5atnKv8nNCehcoDN7NehCtLM0z+F2yygsg+hK+
3IEsIY3yCtGQOknFBHdBD27RlrtCHvT77OwEVHmGgF0cLbPbzsd9Eb9tcFdRfIrl
wRfEfjQG2nyEJBSrWbzTtTU7X2F/+wuOGZl/DmaCTP4z8sRMOBooFWos9bjGSnr/
BG6uG8QgAy9cqKMZuRi1nz0t3xaVHnS68BLazgRSM9rRpdh7bLKPDY5fRNI6b9WV
r91cPeYl33FpxeM75N9cjVIe813AeKDZ/TBkLB0iSbiogE1MXs29/ccJZHF3MzB1
aqCt9Wqf22fUyN3tCC+xp2iEPlJjQ7+swiIDYumlj11IhimUKT6HpvipKpCBZh/5
6h52uDp3cQkekwc2GkSM+g2hjiJvaWUxkbVr3gAe7QnPEKFhpN+tozV2bIBTXA/J
7HRdZlVNqWTZhcYtyC5+4ksdLTKId0MUJmrueQHiWGoAg9Egj0RK4OsaYyrqQKqu
3GrOlNMHWH2uKbeRbX5VNcSG9Sa9ew6j3QdKikD4c+5mjpOVdTpc37k2tmx1ku+9
ix60FiqzZxeJ2jZVq22NRNd1tWgvtqp4RNf0B/M1q/MfJ/VDAijYixD5/23uLp+v
DXRGtBpZuQateiZ82Kly/qNa9x26MpzY7dgspSgmhmQ+PL+K40Jy12m1nhV8pXPm
dHt5XmyZVqYTfZ2VHHxmS8pAoGaj55O5iVPD/k7wEMl0rdZlB+Ncpgtu/trwXiUm
DqtoigFP9ETA4If3uxSCPHz6d0XioX4y5b4mnjnpDep1mwB4UBZ6+p5XA3vmEYe1
2yMB5vc16xDlYp3lQ2IOvuVFEG2Nan+OJy5LKHY5ymnkfZg29nu/8xdHS7/pBqMz
LHrcXXHJBUoyCsxSBDdmj8Oh3YPRHpzHNaQahan2T3IipzIQ7hn8ow+2Em15gmhB
EyHUrU78+KWjg9mOLq+J5o32K5TjKOSEXDRx3YrMCtWSUoM8XVjCdKwgMBTqGJTd
nvR2UoIdJy260Z5G0bGstJ0toyAKv/ql1kn5ixND1zgNp5VW1oB0E8ou44uxJrfw
I6IWtl8M9OWLL7jR5oqvC8SDdAXnky/WZdIlMeiAi98zjVh3YT14Dku+FHC0vF+y
gy/mToIaRBLEKJeqdRKRRUiDsuycGeCpczM6kLyztsfmQIp5clKQQ/+zbvu7SZkm
DT/Pim41LY89XbF113/2kTgmwWNDHHA8sKpM6jpBa9bHyt/dPdgjJwBdqP6NMX+T
oi/aQvup6pTJQebUJ/Zb4xYBGw017Yk43NXFDnCEOTf6p/LOGUL7grLY5eLSS7HZ
g07QQTNjqbunB58Oha9urXlRVszyq9OqM6O1Nm7TDptNTWskTL20VtVK6RtCezJF
QcFlqGNiW4F0yej5N9sketx03xm8gh43liI7uiW5MEqjnBxma9bWrtGwGglDlSw2
Qddr1hKgqsyF3k+Y7eHvnUci7Q+tGqJaC1N4oOB9uXHL4gJa7kfEx++EJpMTQAnJ
sI8fAshJ00+2Z+mVNXmdZIT3ehEugvUaMc6RMUdDI6W2nRWnQocLMYLnwtJZrX7U
Lws6OYOLDSbgpgvG/VfsL81L/hW9alntm2tnaw2rT9GHQmAq3KMtvNRn3QGt3UYU
OJ6I5CCrbb1uxV+zt7OBN2CvaOL9KA1kFso7LvnDSqQ5u1wKdY+cFdBlTiTb8qky
m8dsUzLt64GxwAdzgVkDW4gl7DpczmbOMT1V6XB8vB8+Dr6UolpQLeG2hgX4K9G3
7A91kAXGaw3b5ESOAr2iCqjEBDBZasSddHGv8P8+Is/Tn7EO4tMbLviVLRbkxReT
RZsAIqpmwEFSFqIDUKLZ4tq9AoRvLTERGDHH9y9wL3Sgs4FVITG5zgCxWHiFM9CL
trvna5mWHAf6QLqki/vwL2aW5rj7YfcOV4eZq7kmi7K9GsuPvowWDX4BHIJ8ZiTe
7gwcEJdXXynlcOu7Q5zHyLQHegICsFwnBprS9C1uROW87K8HDeQjGwEYo8YtU1fn
qRnex4tAdzRJyDzH5x7RlkjXlJ8AKPV5DTn7bGWXOG42OuI715g/i32Eg9F+m3EF
CADabDeWzDrF1l/pcDZPqq+dMWKBDcWs1v+H7YL7V8GUgqSaE6wTCOlC5xMN9Apf
HvvaXe3GUt1vXN63IhhR+Uz8pv8F1AwM119K66yn0vfVABgUCjKiAYyqQSLWKqRT
FtItDcCxcw9pHlpi4XvgvpzGjdLIhoTKTXpy/6io6qBxGLJFBLJn9s0NTocB+TUe
VStJZ521EGsNI3BbYpRF5OUH88vozqy0DgsXgkvHxJWTemc2QiK5Sy6vGX+M8X0r
iTsrtuMyBXoXdQypT2/Fb5rbioHoEOhJ7l3+liJ8aAP1KgTJUvE7yL7aA3xZhIy1
sdIsQ0s+8A5ZNLAQDbviJC4i6mY7C8d7d1iDO4wbVK1wYppPVVA+ZImnujzW3xhh
1uDwtPx5TP0ZzEpqwq4RuAOcRdJt0NAmWp8LhkK9lkd41CpfuLTfn3knCFvG2rSA
8CzwuoerMPNTliFpI6lvMAcUD5qc/7ZUBIEHdeVChkWqRWm45vdjRb0SN1dG5S+0
uyXt/4ZhQD2WuPpp2nzBbza9if3J4xSDVva7chR710dAopj7d/VIeFPcWCv59vXI
HH7fi97c6i8+1GZmTEHy2AmwgAONR1VGDShXRGmi8fcd81UpSNQwglrWV663U2LY
BhwyOwOhzFOhFK7EI4V2QpkfcZ7vzqOZb4raMwXsmPlrjE90A3VNYCjSTGJ/2PWP
SyfkwgPzYEcR8LJ+ETlN5ZG5wYaLqFrQp3hQ6vWpEV/Kbpwo9oxnqJr1mb/QPHQV
o82PXXDZczqJyj1sfOllHw1uqsPsCPazgHBi2XGQCUy3ytxKHaeftom7JLOse5vh
P9agLzFv4X0kKzL/7P8xWyet55twh7qqp+Mj5QZlbL215GFGiJkcnpJiBXF8Lk7C
GrSnajE9Ubd2JcUkHw+ObogxrjcDskef5MadsrLMMRditSuEBQtwGbPpFAkwM1vI
2zRsc1tRXtFTrgIs3V+q4wIC3xKj5MMN4qSxuepPAUrZLncf6p2l+++rfdW1EZzX
5focJQsDMK9gX7eqHEeozscBHuOT3QBMZalAHXszalUKKV0h80LPi9sDktjgAqwa
zA/EcgAvjk1Nf8nwLCbJy31moItNnijtO83D+aQr7K/MAYlldxXO32KFaH7cHPu/
7Ju9w+mqzOTBOjkQJEvxvRsmg6LQ81+6LFJcAAGtIhcEJp3wgRV/+CobLVbypOm3
iDMz4AQCivJtuOeKiqFkEsT5xKdwwvxU+NvfbDv7RBjBqnLq24nTey7100Z+v4zp
M1f8MmFigGv3cmGT9j2kG4Ea9ALQcdfyDwAndXzvUxcMlD2m8Oy7Yk8qoME5sfu4
w3Th/+rWaQjiN5iD0UU5e3lS686kMtgK8lCBnIT+b72QUbr00Us6zY9aFXl2BJMi
1/bxGsqvnOdjvDFPS+RspjBDXXi4uv0xaJTlfVW5K8ExU0IbjhdZ0W5lYxnr1Ee8
nhqlNrm5eYh5XOsuqDtP9GMU5VeuiTlL8e8daPDO9nxFc/ZwHW7RQ6vYSTHEeAPY
73Pt6IVQANqp8X3ESyZvTA9R717JHPKZXFJWgY4bqYeFlLyhbjBRwYr8H4iE+qGn
3iQ2hfrBU6gEd8sGcExpq1X6Wrcdi/rs22wYzsBv+3YdGLtE87Z403owyW0K6MaP
R8tqHrj9VMkb+OXwbyGmDRVxGzQdinWshx11M4s1n2ZBLsA6XbM5ojO80hxrqj3F
1DlpW40khgsKDQ85fYAUsRBCzWQz1zgxpoiMbXUOKCNR8o/wKxrpKSBLXwxGAm4X
bkeFNgvKvUPZhv8msptrwOKbz0ZQA/IgTEpd1gfmQAlBibol1o6PJDFdsEyvooS1
eIgMKLHUi1vATTTqv1jXXoPZJk9Aycdl+JYQTsub/usRwH1gq3byp4A4G9DcAN2C
riY/oAh9RxKss9bPaAOYOT1VdQRI4vmYrVhcmWQeUxdQn2aPyljHS1+iV1UtMnnI
MyDydITK9y6zKBOkzjm2UYA81cfZGDSDvLYV+dC4nR4UvBsqRbkAHbO478ghlcr/
9ftjrZlgowvHbrnxpNAlga2R6g9BNN2J/V5mEp7XjhmSXw5CCh8lKBDOiDM7vehm
UutcaI8U2zHcOV+Uq+KmhhK4sY0vbbmGf6UK5lzpZ+HilsqntnVJEKJRCbBpHTQ0
AdkWt0IR7x1P5rClb0DQz1P7aGb6+lblQw/207BIxrg6KUFhCs8eoC7FT0d9frbr
N4xOtTzJ2NWXtn+ftCzttk+ZVAn9CGy4srqjBXsW7eZ8S9MA1g2UqyLin2cZ5H8E
sPt2nlmKUgNTvIn3uo6YJKCPKhbohfA5NdLqOMy+zZxflbzA9wpy2+lURELCkuMU
lcsV/nT4HcK0iC+KForzR4cNAr3BiNzTqHN8RpSxgSoQYwOuaHIbExf/HgZrfXBQ
onclzX9xSD+8IQHuFeZNL/B1gsqRbyal0sJ92ZAOaoc2B7ZoSjdiAnoqC6tXGQJI
+I4xk9IYxdjVU0PwJRBSGZ4PS/0qCx6yeINxXjpcoQzMDIXhgXJJByf2RecilSao
KEOB3aTdPoqnLdwcJr8+/M/eI9RqXRmnJs9ti8FO361JlPoi/jFGbhFF7w4w/tqQ
xJvlJWtHbiZvdqGZtrdMCKup6zR429o6wNSJBI7KdtUeHZYmQ7WM5UqLTcts4XYJ
Sfn+tDnzeaUz8g+lv9BsU3okGoQTp1KgnJ1eHGpIsH80k1g6XAnfMPIvLnCk9zEa
uLggZigA3FXnQdRYO4AK/dpjIaHtEuxaVc/bpHNlpEv7m4I7tJKBMJgRRCIml/zK
IhqICjsL8ILEX0/04+nQD+MoZS3WYBo03gbdoHRfeKl84dZ5t9MKdQlX6jwRgT3N
hoB+u8kF86336P/l4w0OsrUF9CqsZer0sKAK+Sk64Mj+1eqw3ggO7cI19N95PgfC
Pi7GS2RN1LOaTN6e5TKnH7NT9Zf9fTkEaCKqJmi8O4V+2jByTzvjtrZ+NOnyLmaO
NfzEqPf2sOH5BTw4NNVnB61ym86mTQgWjd3sTwRPtATB3i/nTK43n4l3UslvBR2+
/ypjeNjXDXcPlpFD+iHX/SxG1BSZMpxw426qhln0/DfOM47Bv5IEbKU2OIGZ0R5M
cWCcHgUgJiFBzN3t8SLQaFTww7nXqLlPDx33VMPCYXjdsK1DtSfKA/m3TO+oylLS
PdKKa3MToVC9j5uXukl183P2S0lmpsAT3idwrEWnKZqomuQpcif6a3R3tA2QhAlk
KSaGzBh8tc8BJnN4NhWHTsWLe7osD0Z7QTSk2Ht3A2PNiQRPgib5cGbaef4EDv4L
5SKIpstrV0xVwtJalTPaM/84vmT0QI2BEmlq70+rQMwnN+MCmUf2ZztO4UWqYhZ2
AUK7Bu3ICXdh15NQV0YiCg+OhNgjKtiGxSBXM4UtDEVfWRcXXFgqCXz8RyX9cLpw
Xgb6SLO/EfpDCr6Q+3IKdHhI9+7GQpPupONk7CYyMFSt6hEUlhYiNxtT/NH7Zd2Y
3B40FJw5c3Vv8kc5cRKWmYmUHXDidxg+2Y8se5fb2JA1RtUhA35LiCpngkWId2wP
M4Bt1Y2WrBDsVR95n1eQ5eFL6wHAG/2l5fL/dOie+MLNpUU1XfL6KCbH/LRTAcwh
piI3Lfwxf3fgCmj14Gj9KLQX0afWyi8x4JoJVxhvLwB0e72aTvJThMYER3TAxUop
2lifCAOsPSRCjB9ZM7oCX1Ely/7xxXqmcudbZhD50ddkh+zNsCBpCN07xSNrVHNZ
WiwGGiU/ONiMj2p2rhFEjFcsJybxg0vob3jIw+bPuXmYbQJlCfMa7sQ67PTXdBmx
mMrkI3k8SZHqDOxNCXxihw4zGv/yMtfEKc83q+f5GrUiqQH4ZKDj5y+EZYGlClOt
4+vhMo4qE4ypGdPNgZCmBdbwn+qy7TAqxQOslbplaJrEa9pBOt7HwyhOcQVld9ag
w+tq/SE7FhwZ8xUN7X1lJZrF7XSdqLAZ1LVfeoEImKSshVzHGxcnV+Ao8jA2CdV2
gtER7nBN7Ypw6fvMk7UK8dGwR4oAi1+kOGT0UP2qtV1JnobmN0YfJX61P9amIaFv
KP1xYS74AACGBCz1A+SfINiDq1G2MiGY0KxEndOGlvxGyfYEiuK8QEPseFpyWbiP
WBqhhcF3siLAYfJ9H7IjGoxl+R9ABMop5ui3Di9dXmHauhrlMXQk6/CriPBXJyLK
d7A7Ml4BnmYidl8a5VIUGmRjPAVZYWxsMbgv1kFrv3QqiCv1eIJF71L/nKZdKDj/
PbRWitnphD/ZUZ6UdT9hqJZfAiUUj7e4q5b+PWK8DS/hrHB5+eFB6Ba9C8OBQyr4
LefIFflgCcl/lkaJd73ClYFTUoHLInnNhdmI8AUN5F5+JKMVHKYkV5B31QSbw4R+
OBiFfP0zNbNi+Ndr+panB0sx8ulJjZCDyYkqfapyPpBWEAJdsiNFO7ADtMWcUIHA
rcspnwUFb0gkV0y4k+fhU/PpOBGTjSDOkz2rEv4T0XenAn+F+iu5OjeBjsUeIdZh
g4MTc8ra59BVXgDVerCYUA8beJnmtH5XVWiuduBJjzTLqpDzUYWVDisFz5JTwL3m
DTSpw+fgoGNuwt6Yq4Gq0ALt0FHSZa1XW6cwyF7vr3aNW1F+y/DYHfXWj4Au0seK
rGxSEpZZxAu9wv0KLbz1WWmcTKNEwzD9911KG7F8JE/dcJ7vUtbyA90KM2UxmA3q
4LQTtJu/TtuQMe+nn0/ZxzmIxf203Dk108oYwNF416KHN3Y+Yn0FtvUZw9ZFjDqE
wTFcdOKtk0vn+vKKfiU2JBWjrG99NLFBTUM7cKFzHEs9mZeX9RDE8gCztc8zZR7m
8gBOysP0qvJt91Lf4OPzYuCmR/xmG84lPOqUlDblbK0kWbciJohPJ8YGcrtFPKyc
CP27k0RLH4pz4GQCcniW0isJvd15gAPHYkwiOpjoow951I4VpKA/+T5MI4LMiCgV
NpYkCtkykEnvjf/Xpd4LVtuS3QVCEcsop8U9dxobw/jbOb//9w3GUZN9aKtg2mvu
d5TzvsWaghHwMH6PdlOMapTOfvQrUWDmqFAdS0dOFZPM8nY+XlrGZbealrfx+rn7
g+KSG5gHApfg1wJIuvnErbN+jKX4DtTNsGDXjZadTeyPgFt+XlRrX9p+MpLU2Fv3
WW2cfI5Pduy9j7PQbaS0NTVtbKB5mR6FiWgNsxuYg4n5G/7Gcw/5AREHjVhOWV5H
ww/A5EUDiYyn2+baXPlKkI3jx0kZEmJJDAYH8HGVVZI5+4tHl/fziCBDKcKNNcty
3Hif1Vh+/DjOC9MYxaaxXNqkMAOHCVw+EIY8rPW9FLbdXNj5mzVN7y4kjN5jri+7
jSK8jar0r5+2JA5wErRlz3SW3CFYcMgR8BHiPVIUeqImYtJfykPuZ9v87ewC9NB+
u2gBpT6f+GTqbL5kP8ZFJGAlAO6U/Nn2Kxst6nrJl2bfdADQlPzL/DVIF04lmYAS
vzR/pB6eyIS+S4hinaZ7/VIh3OyiuMfO27Dg8p2csv+Sg1qwCLyTdimgmxYgYfug
vD4xMDkX3UlyH4YZEU+mW4ScQ7JvHEzFedZVE+D3jSsbK3vNDlgorGBskidNoo7s
GOtYp2THMsrQzyQAEQrSCR4RF2IwHfNkovlyQ34CSFFHE+/JhRepTau8q/4w0ih8
Kcf4XnWC1tkPboGMqwORfrVCUROUlbTiCFRK8BPmS85v1LQnHpbtleNTOjO9QEVT
aGkdIPI8PjK3a5Na8rGUsHK5C0xhsZPqojGUjIAuWbC5/zBAd8rQwM0hR/5y9VPh
B2DkKMy2F2/VMlABqZntNx1GSBLIUknuvUoAzqxZWmXC0s91BOcqApmaYGCFZCL7
OgEK8Z/xYGuFLyJ+co7xrhdWzTwhmXcl1JRRRAiUusO1bZ1WqGKIFAazaF5dKcX1
c5GEjExwxbT2D/iNfcg6kVIk6jcbvNSVm1F+SO9NEc57IyhdRHM582caKzgULAoT
ABJkc0A/QKOCqU3blQLAfxkMl0gKulhD70f0G9lK85vD1rJQ1X5ZnNelmy0S9e64
zTUGZXI44fdOUM7NrAXs7hmsyIBZHp5ZgBuwFLpScTCOarUHqM4aBz9DXAeTm/1D
tBOXDe2aF2qpJGDrPoilEX3hOi6jJO0YjOGnOWg2jf6ZYmTvLwNht/R5A4ggB4p6
rh1w/kqpP7kYmwSPamP/D1HnGyngf8vEmlXiX56Mdrmkq83ZWIFA3yfbIaE0CNxj
14ZoUCZ3b1oXl49kWMbvd9l+olp9gua3zqSH9odC3Dm6/gx80UKUwWB002jLfUZf
PP2YFhcA+HOCRuDuiFOTR1Z8tcrA7KjaUObZgsYJZnRQpg7EIMDJC2HOnCYdVSR1
Y944fBM4YdHXQVFCsxFbc591miNZ30rD8tMXHo9LuwZUzQXe8uiordbvXMU+eZ2M
XT8PoypcYixPky4l7A6aLy3gKHIR4IRiyZmdq/sKVEsxwftgvlnN/WQHDzOEiRFL
thfrBr0OhgWn8UEKFZIe2zwBho1rrJnsJfQJUeNUDhk8ghV9349KX/fShEJ2S/vl
MJ47c0LlQaKx9yEKPJHXgKjpYH7TWsXGN2TDY1qiU+UBZrUrww1UOsR/RF0AowsT
TK06zYLiGAdjgm7vWUgKDEeAeVqQRcjRzcuKtNptrQ414hGR1YB832j8T28SOURw
7apseDXx6a/mBU7dMSvroLPanJyTsXAJM1/VGwR2dmNJdalgB8zM0OaxaTJoXDk7
YH26+zTFr50ROAOXTtqOXIxrg/qXg6pQwv+nl2WvJs4+N6R0x8UqtXrX7rhp9O94
eDngOdMEeOaMDj9y2EMpB+70V2vevMq0zhZTjq5uWxp5GAdDDYibWq1oSaPsIaqv
0/qCwFTlmrCDwuNkgS3WQn/pKktwDGMAIwm72L1dOwjF0Gj8w0JqdPDatonVOK0W
Ryp/fT3UtgyTRohDSgckwvmAhQsV1zvt8r2c9y+O1xGwAODlvDx/TEucejSkSpaT
umJ0yLVT0t0phrU3AxifnZ3j0nCOZJA/FzXhaJ1NBWzm70KlFhPooEInDJ+tlZq2
RQ39E0GJfqsVgLrmk5Algd8/KdyblzMs/ZEkvSG3EK1HI77Cfid+tM1aFrYBKuDr
r2JZdPHsJ7KpNNAuPDdZkuqEBWwS7bJx8tCj1tbouRllbMYDp1aeUfQyAQ37G7Tw
pGNC/alnigbOmFWZI/WnTShIzoV/YygsPNp6NkjiksCxkx05CKaYYm4LVUBhM14F
vIKA7HZsVfkRqPUfi59G/t12rljXW3VpRNPuzhcQfiuaxuYBLuk0eWUY/e9VxkpY
Fas7JTS0DDfR0GzNLNalRcrFi8lCBJeE/By44v1tKDnffOpEmudB23rwDz7nYyd/
xbH+PCLW+IIl8LQWNHTLeHcsU8Xlsbyf5da5gvP0ql6Znd4HWvib0QdPcVKU7MvG
KZ6Bed0E4tt3LE2vPKYMMJ6sA7aE2b7PDVMm055IoZbjc0HjEwN5N9x8fXDmxiNu
ui5bIquIswI3KK1FsFI4hUGIA3INy62nZgAnEYLVc5OYAlMQy+hUc17L9cZYSLLI
HDaJjXW8NyIVIvoHUxFPf7QwzCbxak4EZ2yN62C4HEsUKnPYxIDVPO007yVtjSyX
BvKRLGCP8gean08ovPTmBd5HScVOmmXTevUP6PZpB2cDLARmgKRZKv+XmUptNF+8
p0Sn8FnmTmnaFZYNc3QicE+vw438L1N/IbvfHa/7/5iGGrvJrZ5n9Ml0Tz9ScDIr
cn59taQIlfnBCx+pcgpq+M6VpP2KegEsyS0RciQAgPKeR2Lf/34zLAlImM5Yy1W1
Le0YOwx2uLyZYv0TbAOTmcfqLP0TQWG6/P2SsKeeBa1RSMJ0/1Bs+NEfVeYHhWPA
omxv9+9Sne0+4am3oJP3VB6o+YtEgf/sTWR/hZdiCJn/4UOyUvstPAKGLjcgPr2S
EYq6BlcHAP0b6P3l8GP6ft9UnuB+5WBwcdyIauERwWkWbiwUlMSVp5GtVini3BHL
DhQneuRuXkFSXp8W9wed0NWwDOfTY3leYvNczjvmOpVDnf/lDxkUagZT9/eGcZZi
0c2L38NoVlbkMRhBL0ru8VpLlwgIVWh1vz0jqW1xsqUoxHjqnCLhLyHWsllGv1bY
BL1LZP+b7cLUJK9aP/bkitGLjC4HKdZFLkk5qaA1MUGS2iuSuTqje9RmahDY6AAf
jY3fMo4KDxs960yGx9v0DqJUT7XMn0AtmsDaGOpSCFoOva4GI7zKTw4W0dd98vQ2
8jaaWZaj81a700+FSiO1WUTSDMDpLrqOLgQVCEEYfKIl5KR/4jdOy0nPcm//D+77
eGrTYzoS2bjTu0ijCSbEzj/Q4E0wf4twap87t00y0zxQsA23Tgzj+/eIttk6gsGi
hPpRoPjYs6eKiBWvokovbBgMMXpeg6kX7/ch86PWESRHSw3gFHDPkyJoDMWWHgpq
8ArUYnD51Gj9iAEkWuq3721Tzn9mDROWpmxne4T2PNfEKtNDexggixPVZe1usaky
tzTsbifiU65jU8OaOAubo2eVqo5Xg63AdxtavRkxm8l0npnbmVm+Vb0snDZgsptg
/WgPlRB+G+h0kklcOQVjBqg6qSsXGN1waRkfPO22x0fYkKl2OCxGPjDj1Pij7TNW
9etYmZDM0AM/ZD5VZYeGhmZ+El8wIWkIbwVch+TZO5SxUmcf9BkVz9/yr2B1iAFN
Xfw+8QbWJxQ97zQeyRG6jgewFmvwir8FAenoK8IyAAgQk9Buz8ee9E6KZK/FJubD
AazKut59XmH/JYYojzJh+AY/wg7DUDcZndmK+uRiUjKfwzwyOyyvht9Z/aYinLiz
MlZLr1+DgP+Ka78UpNQZgNdH1ln2dxiU0oudoa6E6/gNiKu9z99dNWbGRT7NHobX
uw1YrdBm4tMwz4aYqUJVgW4lNjpb51S4LATzAoxfcRqkksD0yr19u+eW4kRbWFKQ
1XGZXrY9+HW7Su3QPFq30b+aBchGilAtcZod3Zh8heFYZzV2chb1JV943rUssaoe
qi7q3yqREIBVD+cJ2uRbIn8v43OIiZqJLq4VjkcM8GWpH/eSK3GjTRATVIpKKrEK
en1rPdH6CQB1kJpY/a9wijVHBFiyb7Kw0NOgNgZ5ZZhn23NB03pkh4VgF64I45fR
dNb3ZHRL7j5Vbj15Eio3dpUKl0ge4aeK8Usw868OgZAFPXBP8hyf+0S9bTL2sOLy
0ZBqGC3Qu6LFRjW+rvh5fk0NBtc7vHYwMD9uneQ+HpfXOseX+OA5qobQTEKzwMk7
5pcBbsZzxR4Vr0oJ2mLpUzAkOlMte1x/EonoVMJ0aA8pLoqaugCDDnNk6FivHrRx
jX2f/TIT2N/YKFl7h9N1f2yHqapAbf4jh9btLzPC/3vwataK10h5AvG3OdIVN/7q
CvlZfNM5v08/5qQnTe+t63pkM25oiXWPornAfFMtp71rFQrdSVTSfWLzZmND0eax
b8f1N2XKgHE+T3EJHh9fRzcrT7SyxOtbRsuotRq5iDR0RtlYro5XnptsqZYxLYeh
060Yw7aj6uBTSqh8OG2UiXx+ALyq/vUixRqWwkKEjQSF/BQOSxSh84Qnk/UDTOQR
Zfd5GUlh6a1vbI6Yu1u4blMTYTjNVtlEpbGfqZwMwOKmLBFliGzmPUwPBo9kPA+M
uCc8G6muPci9BtLqQwhR2tftktJ0oK/pgQ9A8LRy4GUxiCtG5IH3xytskyneKTLE
/5sD0/raM38jLwT1ip4xHMjoUGedR8huNuQYJw1YjnKJPb2eASsTJONPDh6MYbCm
Y9aiRDeTFaglAQp7jWMC5EsaH22RIfX0Tf4NktmYTBLBN3M6gEcaqhy9rh3EjHV3
AyudFr172daLzT9Siaj2ZFqpTAc5bZjJfZesF3ajTgxPcYc2dG8U29Svyam0fpim
9imyy7odI9ASUvRxGPlRBJLPOdz7+oKZueajCFfXm1oRaJUpDdUlCpsOzuYa4Qoz
Fn7xOpO4mOFYLJzHUwxkalw+zsup1DKG55J+V+VypFMnfpFLD9yrRVzIfvUPm3i6
THyFrvA01zApFtDzmNtnieJgbsXvtqUAgf0xPifrdkNdCXF+NQtFAkggQeWUyd7r
x3S6jilIgygE0J4oTs1qdHORYpY/2fcx+7YlxWFwCokGwSN3UBOJNnLjQTKkEbXf
Dl6oQiOkx/E64L9VpmAmOlcOctNtToRtVEcDCV4AaanBdBvXULRMeAAr89rFVvwz
71jLJi97n94tGL80yieu7oBnafIIi1lztEYLASOZCdJfqXszzekAdbCiz3atUEoI
KNJM5SVfa+rYhltRjmamWFzhNYG3XAdZ3hcY4NSqPF3tLKLTANt2+AySd0bkLSgj
LeAFAKs8+YVExImC3ducc/n0/EW8w9i41PuXDICoSctMv6HyonqfMq/Y3lKivRbT
bJ2C4s4CQsF/S2Fdpuji0xa3SkHaMT5M6HwrqHbqbTcDj4+PkmRbSlh5X9tUbtJb
7N3wKlPm6MqHIfMM96kNK21kHW9jRXMZv8VpcWgc00bPSE6PRuy4uoW9so+4uhyN
EkouEE76REu0oPFATHFdZZb8zmzmVzMSH7MzGUazzHPSQqTSO1ODDncR3njv+KDk
WrYFe7Rb8wUQSnbmNuvaGSQ0c67PgDH3h3aJjFKHep6xBL3epB4JdPc6O/j6g2gu
g8PegMsF4IObNOntaSTwbvbF60KCnw4C8bOf4pD5IoPwgIFhV6X9u16jg9Vpu1ZG
oZICHlGfcZz9n/OvvzDJTcrIWvcQtxJ3IpjqXQ4qqKh4elO5a3k5vU5tcxFrAbp8
XYM0XgchwvrkTEdcALiQPfJ96uq5zRXoIYUILGYIjJiKZdB2urlhevGSaxynW0Qn
GPZHMXV23fn0k83xsmeivEpKWVbKhlruHxICkSz+J/tSpmZRooXKW996choqXIsq
oljg1+H4N0oe5KYZZVlvh8Xu3CRfRX1/MvSX4IEHlGhyGZSxDuDSSZgPx3doS5Qh
RAZz11a+qiI58c0juTb16d8I54PM8z21FzfVnakH/yA+44ffLMlNBKwNW4b+ALZp
LRpq/et9guSeS6sAt01fiVEm+PVBuccm15OWSMeapeQoclSNgO1w/oYb19ro1Jqx
JJ6zzNh3NXvZcFFmJNPXJ8Whpd+ZK4VecmB0XHtv5RvluIdn5CNxqGypJNdPZu4Q
rbHhrKUL7RyPwKM7X0HNjxeEexnEstNEYhFq29hgSvNOIWVyWQ+uVR+TSvJqUuJK
S3/e44k1w3wQ3hJUQmfRDYv6bfyuGeCOkZz2Sv/0i+0Lod/qRvFqSr4eGxWo7XWy
F+hvR1AT7hj1sKBBunHj8rJX7EOqM70W5UyCGF0QLvFMaT+sfbVnTNOgNy6OFABF
bs+bUK7DgEE3/cK+kR8HQBFtmIGGgikIBm2yS+NJc1fVpLd1TZ6vnwKs3q30Pnld
BK5xTPyW4n8yJw1jwcuQ5QJ5tGki++4gAUdmB5qBNihw5/0LLk78ZjUlv51hgSEq
P70x1HIW1ggJVSZ/nOrzyPiGqWkVeCwNaD+iX/YO2jR0UEotl1O3xzlYQAWnYG//
veqVFm6VsK+9FXrIw6rNHr2RYoPuWC9kYsWdrjpRYacq3oFJM1u9n6sm+fu5uQq6
00jq9krDHJvJtAHQfGC2NA29zZThIZwk96kBW0o4+xEmbbxpz8OCjVwDyWE80AZl
Hc6gvE03sm5/CJQYChLjygbSm/ndRJ06XHijsnMsJGYQCFE3RFATzCyS5i596614
RgZUd3nWgdVhuAShb39mxwgcgTuJBwp1XFzx6FhK1oNZRP/1c3Zhe6zHwgU9aFLm
E5tsfnABga+XUHJgODHnDi2icp0dAtMPlxeZKUWFKrb/zjSTPRG3raDPV5MQCWrW
iSgvVkjM5FriQHs+FrD1EpyKhPl5xCmfgT4t+eVzuB+KzNS8d1UF1KXx63IwD5DO
ZqL6TungNNcVTr7asECajoY2qQihdXIPWwR6qkPniw/zCLC4VHGLFcFCU6gA74Pp
qVqJCoSgiN9hxgqOJsnSe2nhAIvS+9oPXuAHd053Z5VBR+dX/r6Yh1vUz3V2jp3k
g3CxamT4FCFz9DjrHRvz7tY0a3QcqP1sdRruVc+WRQTdu8iEGlxFsx8VqBUNk8iQ
+MVMbQiRBPjgx9jvb9+kbFaodyBA06gtSTnAHIl9+5Zq4Z5pwCY1pUZXpY2GYZyy
UHLrrMEpK43CqnoZ9KR6uzgYoZAPcnZNI3uQEC3fZ0//sf8+Untq9tKrZupS8t4P
rYazo9cbqKAXAUXKTuHEyg/kn1WDNdPaydMu1nBylGraYjjql3KhLhVsPRro5kRN
IGtlV9QqN6dfmRJvUBfiTss+KfQj45BWxDyEI6ZN6WUevH6YFS6zToL74IOjca4z
TnzJsEZA07kl58ODntHllGVJc4yCvqtCJzp6cyx8taMkSJhL/p4PPU45kvwwWNAb
MvZzXuQN3fzVwmFeGyCEx79PdFP7GqcCbulgwIHdaWZv22wzT8ZYpIP5XUEdVz/a
bVClRxIvuGxRLUVXFDEzrcDXef/JVsQ1tWIONO7TelKFquwPswxmbwgeZejJRNOU
T42S1rd5yxzp0naod5mmzDjvNnTPFunTZaFsSnUnoNC8gBY1FdDfC5yqug5LR+I0
6EtF7GY107J/fo5A558/MPxn5KZ2cFwIAGzYeo3R78bJTg3pBc8/7peDKY/nzF6k
orLZtuZFWaBMMQ0Joz4DHgr47rZh5/R+faBmaqLYWH+dzu8KZoy4PJmZKQdQGx2U
w78w31sh7pSJXHuQtaiiVyxO3mkKCxAmL68sEmkN06s2owPyV+YWR3fiY6EIbHgc
bF0PSg6hVgxEC20/jKgQIiz3bYs4Bmzo0VMT9jMnuiioHa1i3VVF5Fi/fh1SdBCx
iR6VHRUpm8fJaiKwqZ+UkCGfnaFz3gdDJimM3PvPs3HXHFgVInLJW9xW6lqGqb6d
SoQIpuwPccuckjJEdzn0uCDBmT++wWB91vy5LDAReHaruLmNF33knYbTWy1KpAZL
tDutBq8/sbM2+DR3ki6Xb1+8Q0rNJ9P1wioJWtzvdov7ZV3Jlt7Z4C+POpdjJIvO
mLkHQy/++IyseUPOP7WAlO9vYsATgT4h80C7BAp5wF6n8+uwTRARjU3hETWtq3TD
Tj3HDm0eMClT0rqENREna2L+AClXtb6bPBmH9Z80aUizWra/hbQSzRtf4NuYYKDq
KcU4qbx2vviuWJW6guuZ3LBGBNxMXzbs9TcwbIOLh+eWcVnxQLlG2fahb07p5que
5LOcHuBIjGzlDWRqnsaTsuNLkDe4bKKhB7RswIlnPem41RFwLGXW887suMclM8fl
GnVN877TI3uanTRpqNWrULXQtkvxsQK2ethme6tEz2iUkX7RWeOVliLlD5Tfjjwv
+WgHyLTegHeq6is9F6XAPysrnoKN4XUcmPnp+n6l7eaMLuDunLvUJwEsTPz9JdML
zaIwpKISug+b+tx5XFDdU2p4hHDktkgGw2w5e3mclWBI+DTPs9g6T+woDFQ7XzpD
xmIaq6mc7PfgZgq18GgL+3h2x+Mku4tdGPOgpxY4XXyaZ1UTnKZORP4kiXju/CDq
X1mUVwaGSd8BZIs82ZaVRvu+NzB668IG8mXyKD7hGCEQByce3sfn+ok0LKpYpDTY
Tqo9uXMqUoeDVXThZoV9moJj5nD6iGWMDQKUT2NCZ3j21paNS4tzIrsPriU/eR+n
m2FKOIOHUsVbnzaVReEKdhDtsJ5Si6vwte6iG8udH85JUgKGMGp3dnxIIdLCK28b
X5Xd+N5WQYg5ymcsscQJQbmePi/E0pAFLxyaMCoOCjobf4uPfG6lDiRq4d8Z/XQO
Hcg73DXzmY53jc/52mos+StYTtUCYOeD8ZwHQdhTezOB7lqh0ULADGNF/PZR4Ukv
wQL8SjQejGamKEPDue2GRCJnakrHyALOxsqcgUtUNrlcu91n5pdWKoAUe+x0bVMD
iiMmnT0BHWBEkIAp1auXsFCkG+K0tH7fw0c+xidjfNpPsaVpb3MpNAF0oC4roE4w
EUZREpIka0oGNy+UfgtBphxQWgCy1uTx96UTDMcS0NcvnUPtS7R0DvIoRxInUkk/
IDBx94NvSv5lcTUm4rnrBZafbl00IDdS+vAmWJ4Rnly5B9e1xUnhrrXiQfoDN7SE
y4YDxSby/KWca63PBLtYBcngAWkVnmpugKZQQhf+c7SsYzPLZFPfR5QGxZ9BKdBR
fnBV+eALDJn3pnUsatQp96iB/w6Brz2O3AktleimZHsgJpx6yWqg3XNSgmXmODc+
F1iZmUv3xe/RnpYwpFyzjPsP97BE6CO9woN1H3qwA46FKnFuIt1F/effm/My3k15
IkbgIKGxybJ9QmgLW2ow3AT502K3p+YOGtskLgMFrE2o0dKiOqQs9lOu5nikncKa
E2bMnEkZCGU2riCBucif5rGsbpisQbCOgvGZGxj5xAYuXUTaxfJ1ACxLwcXcXZGX
627JW//vrm6fck/yXJRwengWmdQFBRaW0mBDrFX3j9dQUi/TGIV7kGqpN/FLa64b
lUrsmWl7FL6x4R+nWbJ+8k90fLSH+l6L20j/KGNGc2UA4YQlPoylUIVbkhlcHzkA
m2SfmsZTaPJ6WKHRgQAuUEaCx1e6xX8gb2K83u+faoMZVnLkhsSvPa7IB19tQV0k
/GW9a+IAhZM5odES3J1g61MvhgbmUulFYtioQLwvJweQsSbGFdduCBWtq2DkSCXE
K0ZTLB4nUkpHlFJZ5Q5sa2Mg9kSmy+H0CLEg5ApIUcmT2ASEz9gW5tl87XNgxWKB
HC4VkcLXEic8BNKAj6tVr4uh/sBmEhlO+lklaCVPGeVcDal2FCqLqKdAa50OvLTc
VQc75mxFfr4YkwKQMVTSOJyBAaC+geY+T3XSnjX0anRT/OKMvBlMLwpdgoe5VbPK
hQfl8L6RSUCjmhuqjQQ9aVzCeT/uURdtfu/kA+6PaQeJ9yKtCAXUF3T/9Fiks28Z
XJsuN62dsnKqCWAz033teepJbTVjhqJXco4cb9/GEDFmdHN8hr4gXTMMyqduqMph
60cHUUQFX6+flNJRjxjNXeofgDcHsS++EAOyMvwtbIJKjqLmaMVGh4Gtg+fvyt2g
reRrVOzXlrld1zIQuVDmU6XizI06YjceKllrU0zYDrZKbkN4DydqCYgr6vpFPDVz
Xpu3cHkQmSoatxEqoPHHXh/9j5nwpsqKx+yFey7U36y67Ol+DW3q6oMusPlzc+mN
o1gdqmy8WTDSUYCZezOgz2IlmQw8DKyUPXn/Qw0ixiJ1i7JQDejs0ldcaZ0aTISW
YbDwpotsYF85vMBxcuh7gmkA9Mx3ojlzSc5Uxyf6HhvnN2Ik0zgM/Hq9jDTy6Waq
K8s/0ot0/Vyu770ECrxMTSzt2vUL2mvYTrMwm1Z6+tWD0QmDBxAS1BSO/u3URgm1
Lp2swLBvf7yy7I7dz8Z9dFcAyhiUMX43AwtUIpwpTs3K29VTCTObm6kBWuSsxbdh
twlmn5HRhFpTDf6Sj8NSZF/qbsjhqDr/XnT/m1g2R1BcJfAFgI5SLWSruL5w+lZ+
LUh6FpavySzqqSu6OJa9qEWn+DgAv2rdXwJVkVpRshO/CvbDd8dlvVvRV81OO7A1
mY6+DEdYbe/AhnPznedDCBiKz7ckElGbgNbh+yzLNp+i4wZFu4Tzg4oA8lJ4IIjK
W4bKPxA2+V7DJMVtW06W+HzZxQNe7Qhn165+QbMlqnnreth9HUkrPrilikpvCOAd
N/JFrb+ocI+xigGslNaqnwbiWs2pllYxT104fZiKJEGIkrTOKjvRPATAOwWExpr8
BC9G5X2LLrsdPAoLS8e1YH2lu/A0AFCUAqkk8dWI7KmscxNt1i4c4132+xepEIYH
HbyL4mPp1CXibVAYeNAMQ61RkRGi8gGJ9lpJT4Mbr5U/o33lQwW5WJjhO6PlX0pl
047UpDCVZBuHrZbxxS9Lrf34Zq5nAjeukNzBiEN/kyRo3nEX7i34/FW2U8gua9Vo
CZd4ApwZd0E6fThPFmQmcVhgJGqHzw+clMXi0sgN/WsqI9xPt2Nd/fTXZPF1k3dk
XR3O+uI3IZRc/BL3vT8XfPEVfI6DGCj26baVt/IDSNsC6qFdSddH55/exUjho30D
pLpyPwhYKg20hoJZoMK/4rc0fJxtTRGvlTKABdBeX9pgcZOumpXVOe4x0iB0gPQ3
Z4IOhGFBkFqxQsc8kwzT65681uL4Tv9WWl61/zSZYYi8ANViqzvk0VXPgoiYzINO
E9sw5ZS40fAaI9HC2lpfENh+tTJA68veqK/GiW8IZPCh4TAwh7MJ4UUsqlWWQVtE
yL2tNs7eVwMDCffh2qKjpmXJRn5AWC13JMczUSA2gmL7vwPL1wFGVXuIKyCMXFw7
GkXuROikeiP0Vqf5WIGjRf5Fr8VLj3kbz8RFuN+YfPuKrjTLdOScrEk1zq+KV3TU
5NeE2HLFMY3vUzRqi3CSmdooo8Bo1nP7UaS6RudbFrMkE1YnjzjWZDsTPUhpOZD0
w/uWrI28ALJsE0cdiXSXafF14A976TR8qS/VCZruvOCaBx2kmKjCCBBLqv2JhMhE
g5+ixUMUtHysDIFUJ56vqGETAOySE0DH/1rupdQsCH7UpTx68w1hbdW7r0NHSJaV
IF7uZ7g6HMjQF49s6KsUCjqE7xBbb4B6WNFYg04+uT+p22dy2Pssi++5Re1TITGa
zJ15y5+o5+T4nPI87QpXIV+TG06nfKu+LkN1FZcjB/hXfoyHt5TBTnzPO9vtq89m
JYljBDufc0qQ69eOPSF1ymcwuEzC2nfNWMr2kUjHzV6+/IKeAD16cNS4c2SGTOHJ
8CaKLGvxFAvoVihW4VV0ej/KQkVGg88ldW2h3rasxQJMNvo4EAfkirc+5UHm0bac
ocuOanzwvxgJu4bKu+GpByhSIwVPd5vVqbCBnAnY73K0PMRjP/uet9t+1CeKSPcp
MOu4cGFWSYkKDg2qDbp9P0+vFxQ2PqM10nbp8Gdwb8XXXiMlsnjm5fZKZMBXWQXD
XvQds0h6NCo7YDQFEQRx6sTVcXWxL7JI3XALKDD6vlkvWHx7hZHiu3gsUL1RL2wH
o9dP8epiTBxGdvfbqlyf+UushXV3u0UMlVZssd4ShGU5MYYqQfDYZpnK7WkzzYLp
NwXLmwRSFjd37NyiPCZ7eSsOhaw9pnVcHqZVTYLLUgAAB5D7DM1C1jSIn8av916j
s+9ZDRNksjDDHOyJAkxLgfcVEtTUBC7KrCE118SVoajU0yR0T+kZpvfwM2U5mOQN
FkLEd533s4msugtWceFOUdIZlCCYSZpvOqwxKNy1KwxXReDzAo0/i1Wi6ppLrsfx
wQldd1lA5L+YD2M9CqnUHzu1YnOmbtayMyalCuyYZoEEy9991KLmZq7qL2ReRIH9
tFqmUoziNmmlxsLPk9y2GzX2bt01b/Vqw+uKCaoXfTwpqyI9qphdpg6oXcNYBjn8
74/5SSP1MMNcSz43e9qTWd6uWQspCW2xEvO/egsdfiO6IBXbxcR7oX37ZbhG93Px
DYWD0xy6EjmpD13nUcR29ZIgUlwWd/Ty/xzfTfIB87SzvM+HyCMFzeNdhEgwZApk
QVEwXpBK6+zkIXv9CCqs+PO5Hb0ZbHrc63w+sV++LgI62VqqLBmZ9FU+u5PDJrh5
DX7kcKIki05ax/C/jDHW5oHTRZi2Ce14Dl+q7TrN6jm5tZECQV3TBvBZC2vQrUC7
HCbnaijowxkmuDXj7N+8msutXt9yPz1Ajy+lXkU/T3g2EDQCEWNTj2CjWx7+DEVj
x7IgZBMYgiaxMG8Qob3dp7NPo8SpFWyGi0MvsnK2cv83fNpSyWVscs7mT8fK2CYV
yadFVD7RLwT5QDEPyxcVNPlDRC2vT8r3Yq4tgw+emWhs8MlYyJwCkRW8jzyjbJzP
diWmQYWdGfufWJ8LtrEJG6Y94CNVEbMML54byjDZzD8oDGyeMRs9A2SS6VILW330
viqzFBBaqX4ecHB2VPSCFXCrCDlrduCCU/lHQveM4EeJBYPMRKQN+ZrJRB7OErrg
tKfAzgcUXqWgh4rxZEfNmcR09FJnuqVISY0WHWBZemb6cYx+63sLcfbG//q/00Ji
hFjVgYc86G6UQTBKDLLFWF8Srk2tyubWBTXDkmSTJQsFw90h+MTV6mqyVfgCixA6
A75syxoyvWd98SQYH91Xjrrg4E9q1MBBF5DtYLk4SF2cZ/pN204PC0fjdOxejSAC
cNR/C2vVwj7vv/aUIxfkVbDt4hdmMNvHqTt4k6QxU4xwA5ArD1/WhBHNdLnNHnVd
RBF86Pmu3CWwEdBS4XYUgfE+3j8Ti8/WYPQ03lsQd93ne1aY5BEm2uAlCwnKENmj
ckWOssflrYmHH+Eez7n6lJ3M9zwqPULtI6H/Dan/lkxnqAb+rigUA7XB8tYTb5S+
YH8Q6PKW2nFjd48XzchZYoH5Rl6HFW4KvlKHCieC7g3Jw4ZoisM95rTawl1E5J/4
3c62wkzbacymE4B2tJBd9PKCcb8Sv6qvQ3X08YOUp2ZTe2CoK1QSAtXcUnePj7ir
H2fxYX3Lx1Uh/qlVBkDt2co11wqcxpGEoCUOsEvJe5vQewE3felCG1ExKOeZsD4d
TbVOE1b/vJ/b5tleyQbT6oxPLBjFcgrHF5eWdSHn1xTXtBXNk223x9+yC5gPdurv
uINqXghGikKc6xATXZbsu4rGzFgUgEfvkiqNzjoewetnE9uj+hWtpM27Pm4qQVse
vkH1fnuTa9JUK6MBC6wrKO7a34AnDKI3Tm4vQEUvR6G7Izya7EU7aKVmLppJ/U3j
FaUwXq/RKORcsK0ck1jwnf2plmSXIzy7lJkBdgwJ92oBuRpIyCvEyfwNukGhzcoG
VdIAk4M8OnyqbxfNj5cPKsUtYYtmabEnwv4fa4tSvsAUQZ2TXlU7E1hWCGn4R06r
fKrFq2LnuM757Y/HIK7lvHXqAeHrkKU1S4Axo34qy26YW0TalrXRyc7erndd+J2q
C0CkYHyonBllMF5ruFMDcqgCkvPVyMdwNjs1OccgGKSSt+LsiNPKYQ2CasW33VCk
JpoudyzbogZFgtmudr0BZQCSOHazBXnADPrgFn6fYLNNtuLIBcIqXEiG+BXpszAQ
qPrAMnVTj4yVhB4C29X3sSyNW9b4dh7diTylP1ZVx5YwZsXmrYtLUBWU6gDNnaZ9
bomYoaIn/7sZwNUGtt3sjtx3U/tFlVa9SgiYZLM2QYNxHzZYhC+kS0sA2J8Bs0/+
HeIQeWf2UIDOJ8D21v18NgAyts5TWt+o/7Bh/ywln2xNT0ahUigSiS45zrOFYZ3/
W1z7jjMgJNOU4Zk0BWTkNobAWwIoEH++6oLFmMd5rbP5z72st97OhqYGV5WNWsFS
ezStCMqVo0b1LlwUMVLl+b4+LQb475yXJEzfJGkjnSDI18l92bi4PadZdZ9QZaHd
Sicos5RXMndsAE2P8j2SsFbL02orZSprKyVF/53W6D1L/mcYFjGxq71r1CcKphai
/1d9a1N/YfXxYJsn7Ypm6sIJs6Y4AZvKpbkbbyPF+BJ8/veDCGz0Cl+wnkduJvn4
nD1Y0B4KoMccvKlbCP+vO6wt8Jgz/b+m9vp/KItlvI/BZ2XLBayl3muFHoy83EtG
kfEyIIV7uwlF7DfqrK7fQXBlSa+EqZ/GYKNah1Ms1vBSvMdzmJr1Y51sf6LgQG8C
/4JNBOHUcztSK+Owj8lNJvzweeCTfsz0Zp5UbMLlmG4zDmCM/rpNs+T5r6TYcmNF
BZr5yXZauLt6mwF4uGTM5vMw/1b5GSFKAAoIqLGkdSsVq7IBczgoknn/VNgkC2s/
Av4Pi59SogwXjOLW5QQf1TNJfnnIMO+R9UbYEZU3mJKxXE9Ix+ML3Ypmol8cnF4h
6P4CBud3dQkKTCsExVOHJk4Ftzb3u4rbAPF+Vv02O3+nrLEbSiQPL0wj5WzflDrO
KNTWUu4yJnKQgpKjxK11jOQa46atrB+UUsdfIp4Fzf5k0xCNWodnwGJxBZJkRmcf
dAxzJ4PiyLhVuBhuc5qOXE8ftLFqJZSL4DEBUCljTWiPKucwo4rXAKqpXkhiOP5h
CqMtpbq09DAcHlgWj2mTZW2kFvR/eANaBpfU+1MeY/iznD6PYBHeBh62ryntE7Jh
3D5rJZXafStDIBLXvNL+nWBrlHYwf5I9dx+JHE/K5u45IsF8672CT9EU6YxitwHz
dy6V2XyRf04zEdFjhKPTVHTa5sP8eV+9PKzXC40JBkodtA3EMLMA7q9lLRLVvLrJ
saA/JrUYYpIQSFubg6HmacpfwdelK7JAxnsosfibVM9DQguvE0DDv4ANopMaWuOQ
3n09U3s/FP7i4wydrQ2EiM49KjR3LBZM/toLz90ctyXaMeTKGETK5mdxOp6/Qeo1
CXSOcPNH3DVJFyw4pNYHlAQ7scfvQGFxK7Pknkf+MvtX27MF5PX8I9DQctTmYKF0
8BoGR3LbbJFgC9LRVB0E3RU9jbm3bxYGOu6EH/X+QRiZMcGyxQWVej4N+JAQc8sK
S7f1Jd2jMkwdEz77L6Kc7qbzR9M/+Tzzoh5vPT4Y3uuYxlmibLtr8yoU5fWcBQ/N
Kfvb4GcM3lYw1sHDgIGwE2+4NITrmPqCcZJM/SBvIgE4Q+2sODTjk+7IGIyIz1ER
8IIe0ts72B7+lneibsL7evjAcyoWMkUtSPkA+6/zZrZKyCA+b53isNAqElcgnFst
uUMzgzuHdkU6EoKvI5izygslqcU/KfZhT/mz0+B6jcUMVaVN5BC7G/F72y6/7Y42
9vRqjppyUOLoea2ogbc/cCUK1/FPri8qxE7VUT+M9r2mPH6iChlIRfkD3wic4lG0
f28SQTgwNzET9aJKSOnHT6B4Q20ct2teeeYlpn0j44VHPcxIB6MSxE6G5Cw0iiG0
f/qN69+bUc3zgRT41ovEU3RpYsjgcHuk64Vh8XVkywvEjQfusmDR0mzGOZRZk/I+
KG79eOqyQGDZVwexCVY13Qe9M3exmDaodDhMGws1CrADbx1EGvpG+7WJ3pTsJdtY
zpFopVlQBPvpd4DFxQDzB6skCwP+Qz9L5j6qZKmPa5wM1BiSmu69//Y/M1YR8+r1
hZ6qXDWX4qII9b86GRvK7b0nKMG8vAuC8s7/APC2Si7zqvvsfACNnPFEZxoWtfPA
9A7krRwcJjDzS7scYumQvf3PoYWo3OBzpXklU+iLRZjK7pYeWIrvfYU/4Oano3SB
dOSnm2x0HNOcFIvs/wTCuIXSEanN6LLvI7Ta827v84wYToN6buUBRMly8CdWAj6+
xUT2hfvIx+wWnHdrBQ4oqyYNQs1N/b3pjSvVL5HqaA5gkH7MsehOcZAHF+8HuiQ2
5rTLxr9R16x9q/97sWWMbDfOWMLMRGaB3LC5uUG+W3VhsfA3asnNWcfVM9jzPl8W
YL+Ccu4x/PtC8tjlLlR1nepQPHfmIjtSz6VZL5CdSpQZJdPICzKAjWHrnVs3JOc9
Bm6zwbkhaEZUQIxpb+v1gSaykv4tQ3INy8JLii2aJ+1PCAjYTPUYJUkHFwx1tlrn
Fv2Q1T9XxjGyjAGi+EgnpVeSdEnVZJYj9QABhG1Xe5rKebRW8b4KUwHWluBXxb3e
vNhxPcjwMcDrEAgpnqzfTIEr/IxRCV+zZct2zDYtLafTswCE0HTGpJHIvPSQPnv9
nGERT58Heur8H0QdSJdlZQn2LuGGKIHkVSvYbmnXe+7iFw5bofu1l1aGIUfvAH/Q
AJzivW2hSJGfFUUhCRH5i9m9wHiAS4IMFURzR8vDHh2qC0gAc6Rl5R6Jc/yJWpu3
+B6j34+zvR1TMOpHpFXr2IYSaYRHgkhBZgcE4BvcztHSehaQ8B5rSofNISOZRuWt
fx/1hmddvZrdcIObIuf4Y07zLLe6fvum51kc6LYC/94L2w085O9KqRK6G7oSSC0v
mKwn8ykm32urW29eWD3pzVMxZrBRIEmS1Y3Red+KhsnEqA8oX5HATUfNeFw1vejB
6lVy/v1dbF6ZaAj1xn/Rv/rVfF3YFUXzdjchj0vNuYydnVJTDBtW36rBb7tqn2dq
gDzXsY5rZQS2dVQ66lh1sozkPbPagGJEmZ8w1tpNVSNSbTcU+buq3joFz2CDVVsX
NwYo8Gwldg86uTCcuWsVvXoM/8a2zhInEes+pyxMU1nGiYeEMN467tHUQqalcqW3
qvKpSgbaySfALOUcQ7t1PEL3Vj3LW1IFSw/b7puD9AOO/XqkCE+YTiHXZ3Lyy/Y9
O/EvHvvZI92HsaOJxxO0ZaI+vLSsPeYAXpKrmlLobILUg1SpJkeCA/YpWUK90zJI
V4wqRJsheG0yoG2GZ4yxoxYzN3T/FD9i/nCNqf3y4CY2NEdIBpsghHc8amwQm4wW
kREPYCOd22TA723LdI9yjRKdRUp0TbZy4ZKL+KZLTEnRPu5pWPcgr6fp/skVdIjL
KDgbM5wJAFClMAxOAhUH6PQnYVPAtTXTqqRtBrvN7OtSC/+dQS60OoPjGO0UPyKy
EKf/6YqkMObnNNjdTR2Lq7Kec+0syS/ojR4qdY/WAJWiZlMebaG2X0QhWiJuelgr
4kBSB+rGgA2oudUPTeklmv0APLV7jKHOSmDYevJnoPm/TqR+h+1YX++M/ruAncLC
smuRWMQioGiViOjAppRyD0qEbz/tT0h6xQ1G4xcn7PVAP/g0hi4Bnc7GgrqZ0sgr
emlElYVLYcjhd7BJwA0O9folb/sKXdCk6yvUceJl6yUCZmPg7/A++lE9DSnxO5rw
SLazflGRD9DYIY+8ZKTJH7eUgpc0a+/Y3XLRrBcZ9lF439jlmgsxq7rgQR/eazUk
wOropRUhUz0NdDhEVnXcBgnXWG+00dBamCGyU094ksPrDmPgY3XBwf62yJxpnPVY
bNG1Db1BVreD5FVsFsttO1IVn6B76YB0q465JjjstO5vE4KVAYZV6b8GUUTrZ7xL
xtsJ7E0jxXicp3r7F1+87TmLxz/ov72Yj+AmWKmS8fMa7MP+2wEk1f7xTZatJ0nh
bMDpEHlH3Wla37NhNp2b+sS+0WLNgzk+Qy3akLH8z+yP0GLncm0TfOEufZAr+Sb0
1HV63BE+S9sRnD95UqeMS75u/TB2sp0mLlxxSEuZufOBNCKAPhHisBmT3SebNg9w
iga9xZ2GIZNLln0WbgMqD0WLYroYtjLrj8FLarWmshPVp5LficJtmMH9hFhOSLwF
OkDeeN96+qOkqfGqcMCPlX6x1Vr6P2VSvPWzay4lra4AHlz9rMCsngZ1lfRflLZf
ycwwqoeL2qHozIah2fXp1T7RpFM7e54E8iuOVK7Dxy873Oe0zKNuBeeEwmFXURdE
EcGwEDf9cV/6i+Swef7feUSX+7WL7aTz94NVwRuTpIwhlv/gY7YnZT/5+crkDb98
bPdM7TfknDeR2ZzBtDc4NJO/UujilurcAXz83SXo7dmGkzgLJR7a4AkF4t6lZjVE
RE0JB9LAFbQqdyYll0PcM62s9gQM2ILNJSzTwoX6lNFlAMGtxyYr4geWJr3++mul
Z4vq570snSXU0Ew+GJY7gQbMj3s8AC6zRECedFgAfAjTUR2rX6ZkoQcnfER75UuS
kishz2143iTEgj1Rteg4LBV1rUAV+yd/MFzHV9ILNV1OaEw9rSfhTM8upncu9dpc
YWFYL3F4RBv/+wNFqwHjbvYCY91sKPh0YVCGrdTIUApFiebV1/LVX52XfUGx1Dbu
GqisS25I1PBCCvad0rUye/IFhZY/vYWpiDfFKAGGl49i5pt43FGRjwy0hS5vwmZC
QVLzS2FnImZo/yHFcvr/suBcsb21yOKteb470uTTk5GNq/FM6VXNE51Ppeb8sKRU
Kcl/JqGbA1PUPCG9Ql+2nxI7EIPXf9xqTsKvqz8waOC1v++K+pAS0WhXpMLoFPY0
pJizpNOULZWKrnCAIgD63y4U6w0bBD168f+5NqbhtiyRUCjejpGcddcgc8SMZrW0
ArhhEVZfhCUqBE2ZlJA/ygLshuYroF+IVOrmS1XsC/SvDzufKJi0SAJtAjIwVYkT
PVYrBGOxlLXXWLN72HS/UdH0U9iITLz4GdPINLj5KPTvQehmIj4O0pAwC80PQIhO
osJVXakGZpmge8FIBQhTP2kjT76gvpS0r9QIRwNbeZFb1XhTWVT+lG4EBQpFkcIO
5TV8lltwUfCCiA+03XUOtm4qboTE/grw9mlg6nKjvLFAUbgRQr5lXfL9KHzDyyBY
46K5Drj53SD4NvpVZ0YTNpkyzoPi1NkGZhlU+5ph2Zlq8+qEKmf1KNg/ET0PaXUZ
Nm1GRsePhMPAT/uE2pD2LEEPgcwuzypgm9t8AsMT9jOrQkjF5RPpvF9pHNhQejQ4
J6COaiyb/37ythDtKszR7FGCBNjZ6GRTXSKKoxFECu1cF6AiR2bMGBS4JwMiFWnD
7yScYWt2gws2aBfQ5XVugq4Pqdj5DiJXRTyaumphMnTG4KhUDZ74ViCuf8A12GWX
QKEfn8pIm6Pn24OqyvX0YDzsrwngAHZjwNqbXT9uSP5sSvmYc4Lxpp9C9F5RTsLc
VWkcBVKy09BytkHNMg2p2FHs6EA8evqrNicMzFM+gMXh9cVCGsDx3a7pknFx2fCn
asWB1UZ3HQQeVsUUGtpmZTv7dXN026XyvwzMi1dito3NkndcotZyv6DOzSOMjNTd
pq6aIXDSJ83yqAYkVGzq+vPtTrNDAbJPbgHGyfA3TOZ8am+9NPsOie4Q69ujTxD9
EM1iKWaj6OYWuiuRAsUgCkNtKQOxuGe0c5ZIW/9sykqf7YHRMZWv0xiN9UE26d9A
cdxpn8KIynjQfVJfNmpy5Mj/j+8Mw+UIETC8bNA+nmQeGI09Rew089743CgCC++z
iFfjI4VtdQ4tBBtVdCVeLUNxuRFGv0dIL/AjJXpSNsnatrQ2xtSvAp77vTRuARCV
JgIJNgZMcEo7kCjoMpj1rVs8ae/Rbn1hwU6e5KqEUngI1W5NGqptZWL2ePi6ocXd
/1+DLNQ+E8vqUJI5ghziMvemL9q9BNtFXHz18vulAOzXWArXqVruLNoPs2+RaAgv
quLa61l++4O5V5GEKSs14K/procP6zg8/0rWb9ucjRvA56/GDbGG1Sm93opH3qGF
0xj19IHNy+dtrCMocWOCIwdWTkh0d8bKsooKSDtQGAA/uUGjPHvkgxJ/UtsDmjFo
ZeZ6D2aqk9X3bctXQ0e5d7pUNdDtW+/dPyFT3xtuOYi+iDyVDWndCVpuqthKYUiW
fOePo/2aQq/f62AWwusrywXqkM7WnNn3VXyO0HU50my+s7+EEFbj/G00hSIKBtXh
29Fa81bVP/biiRhn/DONssWp2EgqL2Ea1L4DZeYlJv45BBVfE7SDNcC8JYeIMxSq
f02TWf3WXSStvojQgRXJk9FZovGQ8LDe3e6POSfAnBLgYfHbIg26mlrPI2hZFgTK
OXzCg/3jxWvomy97f60p4mSDyQ8YAF6vQGRWyb/SbZReE9MOFd1/2bDz3mf+F+0Q
RF9BFR0gETcryA4Sv+i2ldlUr6sWFh08QKJZCNicDotJPbqKpVaiDwS+5v9eB9o9
JhBmb5kT9L2QxhXW0I5PM7XC8YpTIkPa1oRIZ89cQOoIyAS6okif3M6aQfkz1Bkq
jtc9QMs2nBcZjzEznfSymuJrJz1jEODI7fQFY/vT7IHIGMP4I+ZfCBsEn5it5AAU
94lI50bxOH87Dei3tlKvZoR2gA4PMXzoFGpSVvOt/EkJ07DDrNoti/YXFx73tkgK
LmcOmphxXCAvnFcdfGkNBVlEJdut9ejG6oO520nGsYiYphw/iX3IGIwaG6/TPMaW
L6lJak7FYcaa2g/+SELm/RV6VblEosGx0Y3VD0qmGcqTW73x5PzLD6xC8mRAa0Ib
Qzw7tvBA5+22mSHHtw0nM1YEzb8NfzMYjihYqsvDtrV8Y5PgpmNZCHSayXaDLvX9
rvWRxYqXX8bKvBv/j1g2ezJt7ei3nRymYFUEM+k8co+7TF6+HQyGH/n4cUKFu8/M
N7bDOCPuisLNLy+eKOEZp4FT+OS4Pp35de6KIViO79bCtvdgdGKw+mZDUNAB9wEz
DXP84EAQTnKpckUP6u0yDveYSEPT6hbVYtWFZ44CHJhd1JSodEknhTf12iv1ADEh
CoLcvGYTUn64Q1sWGlciM0x3w7PTBJ+yAuvc+QtGRJ+uANFvCzfk80x6lb7/mUBF
RTFypjU8kALQduVvbEoj2Oh/s2GmQWzHtITEMmT0gPxfVjCbhDkscJk6RDg2D3P/
6/Xo7H2UHgtN3GI/AIB7NnHU/j4Ib9ZxGqi3xBVZcROERdNlBfWAfwMs8J/gm2bP
S0EsEx2p3jEoh2iN2dnWkH7BnrCh3Ow8APJakZ0XqbEYWCf49I+u+zWV1JO3HYTi
YPAS+wLOIR0UmNyq6BrrzQAmfjh4t0K0Ss2s9HByGBgTKzpLtSVCrRtzQs3IAlik
y1gzuSr1p5bkfsNf6leDjJ3lmOGrsepTVNE+RkRZoIYMctdnCfAh6YAnSLyPH/o2
XCUFZ8q1Y8ZmjCJlYbn3kGayFvzBcb8SlpqFY5k+ROLT1KZqvpZi/O8CT4FU2mH1
Q8/LWFIQ8VaqN0xwffbWf/5BFxH/2qrdy4n1NN/LHCPCzUNacQHaakhIEzJGY2fL
fCGzLGqMLShJwlA7PeJs1nYk5+IOWFuoWJ5UqPR2vm1cvJU8ZNv5+/ZjyW64Z2fd
LOfrcGIoeE6Cbk4GwYFUrnv/2dKIr1ZnXFU4tLR33ox6b4SEZKwbo2vZ4AG32x1k
CjT0Y9XhlyCWi8W9400ge+LAIrUzf+jXZjePHyE+PztKcAYgbvTOXu8/Fp4nBJLp
GRq44XCz58wo17IpOqp++yh4a7bUAjWNZrimFAyewcU2+W9IPLu6qygOE0SIbVg7
brJqAAPrisv5PC/WWyNwX9rqqrqDJ7AphZi03qTN2jmC2JYhx1aKvhrBP9ibhcJT
eyPAcp0IVu6z5LU4vgD19rdZngILki1BuqdHapXK6QrfUcO9VC7FWUfVcxmz6w1r
nYGuDSJxDKz6E9j+wWRprnYuU8UZCs54HhTaUttHvJbydoawG2LY5+tBp6TbejUw
7L9McqkJl/zejYOwFoCgNdg+R8rKdWHl3LLUe/eFG0ScExf82TL/1E5SUzelo7/o
4fZdktEI5KQkM1ZJ4Fe7Xb/NcgVifltAu7ezEr4/LSTmvf6cmfsznZRiUe0VyFcU
ZhE39sH/5Vk6Di8lvVCVAnGuB6zRr7spAImcj8kUPuZVLre902Pl2ioP2ymbgiW8
eQmKoreK3dQQexDb27E4dDYEAabZMkKSDC9i7/WoqT0YjhY50pfmNnSL8qdS7J6e
Qkg3eDfjfYaOCq3pDx4MXEYgZnCzENdcYVMnUcOkcr2XeOFkNWBElDdOhZY+Z5Sn
umVGZJg1LpOtJxbC1BVn6nYWsTtH8YN4kdF91aNcV7qwKSy54ZoQz/Q+R5bc2Fnl
qWfwbiFHVrmhYyt1Lxv5kJLRCt2Wfb6ivveUkch9x0tGDRIiHidehXtFnS9GcxP9
rP2a3sZkg19ZqBJcI4JLpqpVFv3ofHrY7xkMjlDt8e06qGjylZ3nxJ3GswpdYuj5
N3keDKtnkp341z3HncPWwue8UgwVF0AmNMOs1a3+KE+R1I6dgogmadWO7XklIcK4
m/Qjk8d7d96EzGTNMO/Ujq53PheACCueruRMiAfue2FZNRksjkMeODqePRKuoErM
5IV4ABOU9LDYj4wvRUJQeKfHxup9fFhXJWaqrGmLY12Gz5sNQsM+DavMGx5adWyg
IVte57Wg98/bXTuHpMu9R9KMCJSdFUylOW8b0UtnomV2NNNxgpUkHnuxTXRMFbyl
c+jvlCW3/8Mux7N1IrKb/R858dID9PymjIvi8W5ZVrLPCosArkATNRtFfoctRu4A
XppuECV7iHIZTRYa8W60qsKvMa/O8P8zYMSRUXlfRX7rkmPxjo20PIcFLV2Gi9OE
AVJCc+njl0qCAWh2Zu3KTQuvys59q+gsFOn8plDTHwQTf7qLrjummuQdoha6+9fH
MJAcqNdocSJvFg0N+iSJbXPzYy9mvbjZMeXjnQKcjRO/eoVE554nAtrqj1khbz8B
Hm8S4uRLh5n2+Qvg3fRM+diwcAS3WREo5SEPHdVacr0gtYRtNC4cKaPdqZEoD1kT
VWInAEUQ08H/uH7AHYKvzl4XeskBgrIev/C4A4qS5hH2E2O54G+BT2uZ/3ivxrUQ
s66j6HQKfLVCO5hwJK5UkJX/SXJy1zF7jCPsJb0Muz8BsV2oyUxVbN352Hzatf/U
xaJ0SXQSa8u7EVjrMlsPaWDoxh5Ri4uqjPr5X0GVXIbhrEHITgHc+orZMawC5iq2
nSvNen5HbwRRAin+W3oFx02L1XcCBzBf2d7a9dD7ZlM46ZynCtN+B/z9fhU8/vKg
r3aDUGfYPQJFBPbqAdXDRiSzrl953xcqYwYAT0Z2YROmKp9J+cEJRsVTDQlwkG1J
Adhp0Q80fQ7LYEsxkoz2rHNLCMd0k5Yqmmy1WOhRXhpjytu7UNd0dkLsp5xXT7/c
UsAfqc1GDO4KPH8JPV2hGs3ngROYs7pJ3+SHK9g5Ek35AncFcvTYEHrnDs0oMaFn
e2A518k9cJzLVRE50mYcj0NM1w7S5Iofjy2LmYGepaWKXez1kxyIxjxp7L8K9MgD
07lJqQ2qPGdBFM4GdLape3LO0FUdG2Tj3EQLEs9lTf1jGlSf6E4Dl1ITgccnOemj
tjD+Iao/ZY4TZmeUgEoEDUhBv35OipiUuo77ANnixDVHcLKQw3bxAdGtyMyDErg7
pAk7/m5zk8WVpcq1Ii0fNB9/EoSd38z6f4doJ6i5WIngoGscL1edVgEBpw/UkGOr
irWrFszIUQMtjp9kKWUHqAkAPME/H8JxnyEfNfT3Hqx6//exjbC9/mafbhEoFNH0
aVmUvsEFQMnsiAqfZ0u+4OaS6r3lTWB1BqSMA6Gx+mehTFKsqBv9tTO7OqWYKChs
mYZoG/q9QtM2ldxOhKWMdqmYVBXTUlw8KZ3xCgBxkEyZsaNvbLRDwfJHk0JrYSQJ
syCaSDbUZcr/L85j6vbjm0ruZmNiXzov9LrFB8Z0+wjJF8FqBESNZeun46wU5gYh
DGFtkdo9gGdP4o+j1P8Jm9RIxmW7oril9pMVtiKSy6gIIIUdp+22TpN1CsdWN5Rn
YuYiS0okj0S97o70VMgb0SQRFkwV+0n76dd8WiayXcl6W0B3hBDvZsQDz48TZpHv
3sQQMW1xjXUOk5Gt5eLKZDhHBsfmUUK1e8w8iEPDzcs+iXv60tfWtLDCoH220R6s
wtM8mQpurysoDJUOsLBhbjdAb7GnF5bKpDDx6RuGR6tab84YFCxc16PCvqNj09WL
0+b22ZhJFV7Oln4XRpuOHhOJnh2njz5y3jOk0pq/iv0lJqqsaKjMW8rTr5HrKCxX
4TbnJnNAxAfbzecvcZaqI05BcUE4WLdi1RMaHviA6Acb4YVPLiGI48wKQrbus/8j
Vn0owJjuevCJsnWpJhea7VYKfsVrDWtpFCRLWO6oU+vdoIJF1vCmEdPyaSBvpi3R
/fhvyJUPsIsa06O48DLXJt5LQ0gGpjJmZ8ee0nhkBqdLJYgIht4SWpNI9y+PC86F
Pbiq/gBm+coISVN5VNLFDbdjnntsITWXevXh+AW2/69v7eIY0rll9K7eF2oQLeGG
HSmIA1MiEE+xx5ji2o3lvpzyJN9cx4pWz4ISdvbHtVYNm/fBOhsg0epUWR01IjK/
gENaQpe2iElT902Clb7Jdk8TZ+wz/tP36TCWFJ4ANvT/ZdjkD6Nh3xgJgsA4MbMf
QIzSFTCu64EhzzXDToAZMKZtGqoIovMR4OVB5mAEywhNx1snjA5+uQq6G9NmQYUX
QbULcLPgnlLvcRY4vhr9PxG5NXtv3FK7brLwHXc2+fWfQxC7Ge7WqrzYTioAtxNc
j2YN/6Lmvy1EcYFyHWapYRLdqYUeaN65IxGx208zRdmx1iORMKXh7PV6Ke+Kbo/n
VKYxcDMad/YemA7qAfGQ3keLMHGzy+KjIZnrpuOskfF66FLjm4LFuzH0N47ciTra
3NLDKwqCejTiu28DYYSTobtxA6CSVFtM3UELsdrziHgfGCc3gBS4GcKwEv5x7oQD
m6YU/hIgDkaB9/0HE9Cxqb72PY/KLQXMbb0xpvKqRVWcn0NIB7kgq6vXmoUjggIS
YA7SxUvz3Uaf003vEcdXjnOmOuecsvCzW5sA3KgG2TxxfKuRA36GK4CNkm1LSndq
16Bojilh9UKQCInaqNBh2nOFSFrZirP309DdsidDqLDyBrZ0wklNIgCHTLab3R75
O3oFESler8LymsphKGfKh1KpjpIVIVp3WPyDT6B0eOQlbRPp8p1tE+nCM00Srh5i
2EQjo7AvmLvgeCw11DiMJgSnwwKh7pdGxAGB93XZBqO8ghUIozgcubEG2k8RYLdV
iDey+gEjVjtTLHKRPZtQHg+UFHex/FY5yIETHVxm7W36N6K/dg7k+kkHX1+FgEZo
rqzamA9kzyEUJCOxS1mISIkHWOf8iz/l3EYSxtGGBFEvew8vrQHiafShB8+2VwhD
pS8fHhuE/EAKLiadKfUp4S3NfseyqQEth05ulBzn+MMz6hFoD279QE/GItlWAN1T
UtvXcS4qSzD9fLsRl3H/JKIDTTUSaVcO8tlMMNtj3VbzjFrqPtcrFeufRUV+3EuP
eUtbh7CLfs59djpQbs+xA845fKgvUc3ihvuG8h2xZyd6Ls4AnkKV+3/HUCAayCHU
pPivb7Dv1tFFqQ145aFHtpeO+bmgOD/fhdDGeMxDzwqPqcqO3aj1ZRRMW7L4ynmw
DE9WBa1izMcllTK9rNVlFQ7bTm0P9TXg0ptyKstHtOoem8t850GfYwLQeodZdjH9
nF1QhWxWNMxp91k0HueoKONX0TiGlx4B2mN6pLoFy4aokjghwqkOV0Ietvb6XOmh
DL8sCr1CYVyRI7IAaobMNSEVcdfh//RcZXYoSOduBRhevAMJU/CBpXkQKf9zVnYr
Mhk9f78lBAG1kYiydvxUXdAH/y2Ke+XGuQKAVvVV5iM5DG6Mt4cHXdqtsLjJtaKy
SUUup2Kbi86W/+cCaCKMZ+Ytk7mX2BgTUyjjEaO+v1a6QK+PLj6iOwGEG0th2b+D
fbIc+q+1Ac4P+hcKkKAQJc2hC5BRkgwbc+h60h27kjkBGMW9qlU0UpG8P4V5PeMe
5biGl/AG7wbKOxF469Dihnt95j1qMB/LKo7ZliP7XVIp7+SoIOatRsVpKoZoR/8+
N/wFLm5D41IFlwi1jKk5TCr15fOwkCliMWNwdERiG8WVE2lhpOZLqqgK/xvPGQrZ
xEp/4kZKLNitDaIokCND0Pzrs1j7JADFJOU4wXqaOqf5BK+mGdNCbU56gLcqZvGd
/IgCxM7hJasBkjQbJE/7ERlz85hy5FUvoYh0f2oy5ir/+nBR5ID9vYRho0lzloJ3
WLZe8fgHb4k14NhTMKtZB9HcIYNtaJgObZjAj3bad0A1TEYqIgpD1uqQCDswZlpa
s5WBmpJPzG9+n3bEx/+WOWontUMin/WEOhJsmVJ0P9Nsh/kegrgFQWn3jSrpj0xi
grRbkwzdIWSspvRq0rmZ7jtU6udvcgxmHzvgxtma9XBl7vIpH8YQH3iYiXNs6FAJ
ksknM3AtYb7LM83eNWq3L48CE3fpzr1z7XqBWjs2Xpi84Z1xP1b6MSoCdg6yWdGH
vSr44vUxBz5ZscU3kyR5Jeb9rfAcRTOBufqpmZMgX0mJWqjOaDo8K6EE8/IkyIc0
mM7LnMNiiYkwuKa2a1zSu5NZzovDE9qjGRcIM06MrCTXx3gPESH6xkombkgjekFk
RfYQkTtM2PdT7k2qet4tuBz7nbc5bklqAgoSJY5QEaFcEPYMjy85J+gYFboIaKp5
+lq+62FKxswczK5+5vi52CkR98CCP99HuxvCXvnsw1OEcAo3XBGlXBsb8646YnaC
irIoAJUA6P3KVEHc+40vcOTs9p4zAduDWKDrJqnTscpXAnZs7khHmsBRlRnSzVp5
APuC9Ve2vIJy+sAUuvyuKkfkWGP3USBO9i2SZ85y22O8DxwxLfVM8K57zyrqd3On
lPn8PnXBduQdVSXCbKjN9EhWq13GCwFyBc86hoP8vz0mTmkjdNLOUwlhutfg59gD
DwDD8kDj2EOeeqfJjswr6DNs9iqE1JP8Y9Y9+S0vZ5pdipaqD7WRe6fVIqGWxPuB
ds5shiFO5wYa47my33m5im34hJGNIPfsXA8pnMGSAwqptvRMV3D9On7m3+qNel0z
4ECQULLmB8fQjC8X2Y/mPesdjhiDabDKiDzNCSUUjyTonxJ8QORA0qTiWmZzSg8S
UsYs7TAGDaMEm8AjR+eORFcO/hqPRsMiBeyndvq6NDKIiStqIRGhOdaMusqazeZ+
Zz7vphu/LjKfH7vKjOLTCItbwnRr6A1gC+pg+GOIwKG/z0Ahz7wVjU74U45BvxB0
YGBSSTSm9s7o/oQisccImg8P7h3iTDaVcAnQUDqUmHBughztQcAh+1R89cMgxwCd
StJKX5Vg4/xSJP2Vax/ClLIeWfYC5u+9LfqsYlygInNBb52PUoqPiEf4o+rnFrGK
UcTSENvvmmC8nxvI7cmSJL0U2Mw8qnp2OJ7ThXm3EgzrVi83mmfguW1umqjhzYHl
GcHZGfuQJHP0YbouHgOBJzN52x/cPr1YUVrUjxZwRsDVaXhyQMQQVVEaXxrHuAYa
tdpoue0TKRYOJvkuILm4wiiVw2qVHtQF9KPsSKQocQRMPKIIvTcQoy1bmVbqYAnJ
2Cfl5mO9A3f5H0z6e+sDW4nbcxylAwO8hyhJUIvBhzfXZWmiv7bBJRV0+5aQCYP5
zRILIaxRuAoHjVlfod+2EB0Va1xWEz+M2WNYm6Ha4bFS36mReAKQLGwOrNlqQ+NS
P/oGeHXcn6gLzx8rtIjHzfkIzB+bUJQ07QUNSaYbP/OUkvm5KSCkIQBcyAiMIbap
aTbltap8QCmOZGU4xD52aHZfacIRJtsLX1kST9ku4OvsYOrAQLOjtnY3RJQRKK/F
VKc4ZpJtdU3zIS8cQdhLs8QPpPnctSaw0lcnRatqWLfXeawDBpPBk0b6x+OGLPt7
mT0I0ot/pp1HC9qkTxYQwwWYWgItD6O1t9gCQAy32/P/BcvfOFqPGpN4lgUmOhDO
itVy0NfCWBo5IUOO5u6kQuPqr3d6OdHY6ADDA1nx8JtVXV0dkgJUpEY6wI6rDRQ0
8WOlon3QwEctO5rmrsULGcUtpeksJFp1el7T2md63onFTnMkw6vkV93gXsqP9R6R
FD8wDuK2EjOUpE/sSXZaGkJOVsg8DDpnFMo3G2K0+sC747vC6E9UyOwXQu97iIrk
X6kkVHVZSrXTIspH8KPZ5h2cKXTw7c+DxOGYOnRouCHd6HoKbvFPOY4hfxFbwx2f
EFTnAFh3rUObNs6hyDBWQYrknH6hv3PB0e00oucYR503QnAAWfm0APIrCkVnlVhW
C1JeB4R+n8FLUJZvslXbKcLEc1OuiZr3JA8k9z1plJaVrzA9EEaswfNCYoVyrolw
KaEXKrZ6JGrJ4CLogsMGfpOfLBwvZJLnaj7PK9NQpnnPoBDWgslfg2HKREpy+4rO
jX9ksAPucxDb/gwuSogpkEb8U6ksr1ABfX2Pxilac62JefVXLKXxtmXC2aRRtCzK
OLAgRHMiG0jjuU7cx0nkiYP5NkugT7NM8U/MmLbQWo60SbxlqPfJE1auG4a3Y3VQ
lMOeH2ks5yZeBVvxDZpOt9ZMpiCYS95ezGCPS+93VnTRnROabjCeaBoaWrQh7dK7
kEIT+gNahdWnnxYl+bp6dQmI20J8Yoeb+sHQaS5PUDr2Qn+gCty6DRiX0u1iEnV6
PZMys5LU8Q/Ff4UxayCri8lMh5rqVJIUCx55zekvDnG63BRRwmooeunailwQITOP
XlZglVXdPsV2nQzpoYGNizVDI7Akb63NdezOy/IaYCfg6KdR700E+cwn8dqhpTDI
osU/JLssfEqigLQhX9UqI/aAzDO/bePo51Zk2trrDcc0lJDxh5YQKNkpyvL50VT4
99pSR11bC7QNAxXG2lfoLIhrJJiA6SubgWpBOPT2V/pifxNdPMGhqDJdbT4z1YQm
OC8R2nB51Ma5R7Q24WvhWmpkjcr9gyCqBrL3kwErCIl1w0o4V9sWkUW4ua/P1O2I
LYq3rDiV4LFMI4SHt769aQegn0AaRYNg5OyE5EVSWaju8rHI4F7ZPpp94XbetfCg
sceZm4+ommtl05GBhjKrshAyVxa0lFcXrlZVuIEZmnGqno8im6efyxnyU2dqcWe6
ASwmzvFiRkr9YreV1I+FdZ7Z4mYi5R5+8rZ/14G07zHAxfCDpfhmqlj5Dr6geeAo
9RDWjGO0OTjwXKLIrdSJ6zUMsz2S5btLH/FX65rgO5qW8E/T+M3Wzqom0vMJzuKF
pZGoHAthkP+DVsfMA0XH1E44nnVPJ0UVgEk32W8f3nSaNeN9QkP480sWTm44KDQn
hUmY/cg87B35xzkypnulgQr7EY5wbpBfu6F5z+enRl/ygcN3ZTahdiEZlJro64F6
hp+Rb3FG3u+lOEJjCujrZp3L6sIAZRQ6FpPfDDDlKlh5h8e4sE+ZbdENRKE4mJP7
qjfL/Z8wjvMoN/g5tQJhbt1uwLqhMK9HXOLQg2ryUn57Ui2Cje2s6Z0v9eoIYCj8
u6vJpKyiv6Co0wLb6TUABpzHWkcQyhNclEAWV42cFzX25+gsxLY58hMCMSBplNrm
J2p1C8QOaAXEGxVEUx2gAv5IogqFtCwdjSk3u9wd++9tlEWMA2o5LERHwTe4G+aU
yJW+z2sVEcGu970TVzezwDasgvipiJht9KfZIvuRpvj7UxQYNPdCntrMgmPiEBrP
kAzQSUSrWacu7l8uCjmiyA4cBTJr2MSQudsZG1fZBI4McoTaOCRt+TqpCqSDvOn3
e+LQadHdYsl7BKB+yjusUOENC6+WmZyB9uPNZQx6QrM7ZWRS7gAxVCpOiMoCZvvz
ou+uslCHo94guukbb9oUeqyMOZ0cuyBFPUWK7HsvC2CWvO3HFAKSNLhwD7PKoKKT
HGV+S5WZWRnajla8/HPkK5gbXD4Czqwz2lntXr3HG4kdv5judxsbrc9IPR3XKhUG
HmYr1H6qPGajPy3bRm6Iq38KAr+i8m3j6WxHfxjztuyMuwCWdhD2EQK40dTKCS8A
oKLTRe2bKfjSFHAmjEqhz1sLmQwffnoSpZ0OxXVgMP2Z2TgfKf9mNATW7DmD4iQj
xppVGVoiGC8I4ZoSetEVT287ZG2dqCyv5uzBZtw/IBXPgwXZ0iWSEdApC175qGs1
RaeyEjmVcSu187kERj05iLVAwraa+JGcFBryuy8d1H96PJ/e7p7n+MuAm+uIEmmj
1JFfwE+lzdaVvwoQ8Cx+QV/hRQ5ewlcmm9ysIcXIWiF7+MFa6v399eU5vNsPnSUP
HYAodyjSWWFajuE7i5pKW35PYYbKu+FgbwhUttH85QpmFR0pt3eP26p9L/N9+s62
xa79nAwNGx6ssqDW3QtWXdVpgMskTZK/azVuWipQ5aLqDdixOOt37jFh6GqJqpJY
7UAI2mO9Pg/v2ICMeUx+en+M3s3EIwQ+fmTEFVEYnvzGQqBf4x5tIytSJPT+sTkl
0MB2GRPJTR3uwJb2mRQmKdSwnMEGkv2WYrli9yR4Zlnjzx/b2uuNsCD3d9NjdPIC
bsQUe4sU3nGWCGn2kVL2yzHKMvE8/Fr4zQUhsk3REch4kdNDktP7MIOWdJyDhYug
4tr2r/1UXopBVHaUvvid5vkPfyr4DTY9JQ+MNggXWg1l34FMQVopDa9LBe0MRjIQ
JIBj59e8PvuPcRZ0yc6UzAGhZX/051109KT2ud+JkF/KJXQS3RuQVJWRUAm7c+MP
5Rr76EyTbVM3b4kaWpuINbKSEzRnv7eXEtuoJB9ZbdENLR/7NW6/lnGUlOwK9B+M
Jq+d2UufGtLVvUqvihVrxuQbgIlnTYqRniiemICBZ/6rXGqi5QUn9DZFduAyNfIK
oQMbUjL2fv7VFR75eCtbp70E+e7ltVd3Cv0yxfGnAnMmNvgM1E70yqVCJ6S/m+vM
bcAdzMk9193jvMdBo1vkfxQrxfEvouCeUV2bpgcABCVDZHRiNhnFbkoPK3vnQ7QU
eAjZ4fSzfHoQGdwkry3u5mZi4nv+hr+JrKTyEaMfM1xP7IvFuBOf9bH1C9Ebtr9v
G3x8OvY4dBBdxZCIzWvP4KLqEd7J2YMdPurXYFTqH4vrTbaXGwvVRmFZo6gLPX5A
WiIpBIXccgfGyPaSbGORhVxxBFP+9CQDVbPeJQg+s+XoosRUaYGwY7OCJ0BH5RcC
ENSn8qs/MT0AgRQQuta/ac7m2DSnrfsxpZbzDYZ8/Ht3jZLSTMi+4lO7BVUGNciZ
E8gIHgDGIKGFYg7uddW9MIMki4bPU8NmUeINzDkjINAQ0o90gfvSq2FLVGVh4qC4
+LNXe+vREBiIFamn/IZyE91gDCqfyuwNrhNFRZ7p0lUbZB+eg6VfikOjCRObxcVL
ZfG9lXaQWSYsaQ+on+kdzi2OT2OyDaLxy5A0ywfiAL5LdJf7n2dhG3c6Io+PaB4W
T2d80YpnrvwjAb9s5ZCzctG0mmpsf2/wgN0aRQa8Jk6XzZzTfpZ6LazQcVpZipaG
atpUU4AEfBB3gXNKzdNi3bl2Kvw2u7g1fwriCgAzzpNgdU5hNwKNjmhBYf9pbHJ9
DQqDaT8iA/JUut44TZCusY/6O37k0U3i4t47zztB3JNH8bBUhfPTJp0qFZjCnAra
AXfbSUU2QsyCwY7VCebs/blzgmig0q36O0llxmwtv4xbl3Ln+IqqG7OM+eeSZwP4
YFFWkNk2Q7blxXaBWvXv0jPGYnGQD1KOjZy56wcVPfGgImRnzsczloKDlXKeBf3W
A7+hyxmYPzvZ8bjgOHtZa5fEbhT8s7ZFw0nqmkF5+p9vkDFl4TvuJAFQ+PpxJaIh
nsbBUQk1S+JFw9/3Ntb7j608aoShtlsDEJZxJtAuY0IJObFKoEiLfFzOTguf4K3O
ur8c6O99FxlwWGfOdoOmFj6JaZXeF29oI4hHioW/LWoEY58hIH2M6AHThkv6xe/i
pZAYUFSoRfRi6PRojVGUsoCU1K2w6fZimSFVOTUFq3RTHLuvTHtz6IKdDhIpe0fO
YL6F7Zfxc0hujmuZb/KJ5B9ogWIhPFIm5NFqGeb7bcWmj9jFk9JGFYSMxo5VCWTQ
ZDGPEGQN2rTGLDPXfZzrWlK1VqhcRxssOlxnOmofvBykvGBvilXVG/I02wk2QfOw
C4GlNBbk5gTOj//X1/RrEgrsnO5ct1rw52XhEbO2W2bn/L5EkBfcQgF5XPzMlntu
2bvlnR/kqSwaUaUGzx+GCIXMh0AUWEQsVEZqWrJqyq0yQakxs39Z9z/qhEi1cwsu
oRCVwS7UmWI77F9oJqOeGhBOSrTOvv12Oj6NYrLnQLKrTTcYs0Xf/PqmdUOVPCY+
2vwLxh4IS1MeHq7rZDG7R8sLVPrr1eZzMO9PupPjc8YoyTLkG8L4v1Wt5KZg8e/E
YnwSeM3QUDYaVnQgkyhj0ow+dvLyyBDKDU+b5FnCiEzBoiEcgf1RCHA478LiEuMH
aF27smtHoiBeckE8c6idUZNOtlyiOrxgITaIa2w7ULnsDIpJaQd2t/bKoom9WnKo
kXWFqvMg6ZUArlOn/H47iaudimWaOE6Zx2bhUTG8+PWRlDwUB2uihNAO2QEdSH1p
DQ7CT2dph7QEwJNaus2cRdzeEPtCRvR+Q8PGMOSLo5616rqxpxhqTPJUMfiq7ulJ
QgLAyQplACUzWZ6zHdQNvqOmDaABbff1VXg/7fuGqZPQmDT53xwWM4MqSJjiq9kb
/WsGOwaRK/xe+fRhqHTACmiToGikup2x6oZLTMZwtQvU8BHPFnjomccl0Cf+kHZz
a3/K1/uEShbkhmq/ECHgVCeJVRAliKrqxJB8pSxifaI34eiiyTRr3XsrtXt6BqtN
xFtE2z/2jD17KzI6ucwbTJS0b1tTmhUFxH6W1wY3FDRqK1gxYuLFoPLe9upkzI8H
iC6MBFoFT7675Bwqma/x2Ys4AZ2oMyfrnOkVKN7SpUvJniOyPS3EiyIL4vc6MA/Y
j25Ah3cDsEOzOTCIfLs66bNRYVMI+OXDXAgmWuqyekprnzPcADmjyTLJEMTAsGgr
b+i0AK8b/BlKj3myiW6Pa142bSyLKGGvd02lAbbRUjzJeHg6UmT5RpRrRa6PH5We
BiyO4OgiqFuiSjc29iBbTmWRpC95qfPsRjBh9gxT+aOw7PA6ansllMq4gIWUO1vc
GU1MbPD3iozq3JgdNB0tRx8GyI8O+cqnmR49FqIhANiZUPzCw79WEL3rmrbtjm7u
JqY31bn4xDtAGJf5jgzHzG6l7et4vVgqvSnEWCIvE4Q008S0AF/rUGlM6/0ab6zZ
K8iObgVg19g15/+KliuRGyiHBpjb0mD7brYF3cfd+VKuEA0bj03Y4B5SDdx36lDU
HYOfTMRtlk0Xn/dljSCIhEo9ZqHKF1jiqsPsCdnN8egmlhP1iwFiiF6GiPZzkLuy
pX5KYgEQsw/+sRgnV8PfqNOq6AYW1WDbYnNOeqzjhpcSr5ziAKbwacfZuHTubD8B
Xwu7iByPgD4KwKzVW+kUOVJPQew/A3tKo04oEgYwRXckgQuQ6rTeGdbvDbQcWgRl
hEo/iPZWojHbqOtUWpU1EqbTczL03SocwXJ18NEhouM5syVOEVQfkzWWUOEhS9ht
mKioPCPnZz8vDuIfbzoR56Itv6+XKqaM9SI3zi88BrHQxYLm5DI5bQMgn+82N5LQ
Aiqb61wk9yAtVs1YTBdQ/VCiKJ6ft3wf8lc/Vk3xwhQHOSBRb4uO1Kz7ki/P8skc
XbdYsO1uEAwRuRbPN/eMOm42k2X/LjmMaOIgHdFZvMnpZkw8Xksq/9GmDmcAA4dL
lTkSd5Vr2JcEpzbkPLysojJm/NGdfBP9WFQ/b+FwXFDQY+5hsRsvXW32gM9LXLib
1kGUeLukEqo/Hv4TUwL0E9v3BsuKAGkNAvCyEgr7cNsP5ryvJ2lSUVB0M0xA2rGF
bVuHyrChxEFBDzJiC4WvxhKtIBJdEM2/xyOxA8Y+iCGprj7STizWee94Rk/nRRD8
1fVHrmScvBBbuRKkA+yciG74onHhWwTW9bL27xFNBpwlhS5izLXQKUKgIE3ae9Co
UTLl8OYsmIRTcATf0MXcxm7NYEQ505UNJsAONxTDDjW51AYM0FkKfGl8MTn6ngwv
LEYo5LyQxmyjw1tKPwEqsmdVXVX2aQub0UzwIQCQOb7mG56bo+Gp10zx0B00jt2W
wS8iKWTEYDps7e9a4Xg/pkz5IlnhCWa4xO32iVnSqWygg9xUtzeeQvjk0tP8jMiX
TaRPiluWsSLfpose9Aj7b18bWiz3BvqEo2W+KJduNYSsC3hJqveUAp+8+w8XAih9
qtHTspaJBFlKlCnqwCilYuiMXuOaoCMKlxPluvcLjOTqh0Y8k2h3zvyf7/eA2Xsn
MsY/KwijVDoo6715tt0KyyPRdcOvAerPv2ScE3B//oqcbxu1ZXcz2C3ocX9huboS
Dou3tUZtu8Yn4Y6Iwcee0dPOqyDeh4M/LR57bIXYdj/mkHOEjZcCKGiZjUxtm8ae
U5fiA7BAcvmwuzYsE2Du45IsK0VvLqbLka1S/9F36/vR5P2zqVzcdlkAkD6+q3y0
DmNs48O3k5/ObrFJlmrOVgaxU5FrdRdoXcdYcegnmDSejcSl+msUK87AGqVCEVlW
kzmm5qlALzy8Z96DZelbZdGY49vV+rVbX2bIrFQEqsRhGzKtj5YyKJk5efFlWQdT
1Fz8OVQKduT1bowv29Q7zSWfwXGRpM0ZLgc9a6lrQ8bJ/1qD5v43470zX0qHXcoE
wlHTA89S5aX+OHk/vAsZ0KrlMUCYA+wZ3/kZ86qYmEsmhOHh84azkLUs0/j8YFdZ
umPcD5ZrjINei/Kdz0vpNX4J4RMYzu7aJ3Gq+IXD1gqXG9RyNFNohN4nVeCDUHuU
hYJOskUNHXAMdn1a9+qH0jGj+sqmm8qy3cACmNpCFjyY3TMzmQGDIBRUPH80oQ90
BdS7cZxzquYpK/TXyZ6pnr6fA7gXJPHe6jBVR+RRXTTEFSUQ/vBGg7wvuFoWsr38
ISSwIdGtovfoYJcsBiVz3ZXjpUftjZRlNJiOPYWp1dRPRkbaqVl56lzR3MTC7PQk
kRD8VJo1JshwDMhXuHWfrW7EDWGok48x+8j3KYPrz4/FuO5yczjEwLyqfa0voQVV
kwXLYwRQIDjkxtcuhRAnZr/zagiiFtI2DUZQ7eJzTWRxteFV79RVcdK3l/h+PpF5
KsqTh2XI8lrMkzdeEH2MBrR6BQ/wNx1aEt0f9TFiChNt8swYHrS3KfU5OcSgIz79
4Q1bc660/9FZnF8sii7R3vsUYJo+m9hJyQ/asL3/M7epkt428iuGOVvU65yIGgR9
5xJXHE6Fg2gxruxVxKDPAQhWq+p7vCLKqHj3JQ3yGkWjwpGD5i2GGPvsF3aO204H
xNp7IN5g7RBPB40qbRRCUQ58C4k7hdbMPXOFjSGnuw7hUN25Pvww7mpuNFsTlzaw
zkRI0v3DjQFp+JCiiG0Viqkqgf5kl/UlQJffpiI0uL6Qx5m/gQ0rf0AO10g37hly
pZzFVSu8p+xPtP1VlqLWmSxSexBNDNaJrErHlehwrU1/ljW3xzFL829HplmTCEC7
diCw8ddW0PJGRHuG3nhaKel2708UeY4nf0/IT4hxExd56NYLUmJSwUPxuLffa7PX
io0eUvqU0vrHZE8ZATGOU1gZ8kvs7nb7UU2vZ6A13O2+mjVHoP6AQqiEdWqwQu7j
D2LgSmh/4ytUjlz5mbBs8afZrgCzwFER2/NVBOZpL6W2g4DkbPTW0IOwQVgDOj8U
g6+Vl+QmeuL4nMiJZFOy9pkEdhRbxW8xKPM4gVkJEye8TKXTT4sQOjgq0+vvDcKN
eVzX2YRMnLo7aLfR44sbIFjHJG39M2JlT7gDry1MyZ/EncxGSIATA7wmrM1vH8z3
xzKjIxGmv2mxpnl9wOo/oSWBWpaPswW3RJ8Qbo7U8SGVY/WGJqF2F9efLPxilJwu
oyEAOwPA4SoyREk/ScmCN+mFbrbYPmqyPcoIyOvgWmX6meWiq8LIrw/wZeH7/+Eo
SoDDbbE/jGGGt2BTUFrdS04TI6HpJB4eaakOkLgzuM3+mHnftXvC1g/S8vunblqK
8m1BsAfrV30SVjwpzH1qVQ1AbhLNkbBD1+BbTPhEEIY/VSty4bcvgIMEPEsx8nFO
chnL370nv6onFnhpNqTGhse56TgZKh0s/3YQBaH8PnNYQsDIHWuQpx8yKIBmpssT
gn2LV2nRyhhnvWrxpljK34UnDNdFDCU2lf4w3CeuWE/aFxORcG2ohffBWvGu4I3E
KswNHBf/kqtHfH+X3Dcu2TK25oyM8u1WJUjXtcsRPbq5YcAL9gDpgh+AMOKnFugD
spzP4ewAFFGFfpfxCef0Rt7M5DlzkSm4oe0DSsxsUXH2/r7cWgb4+TN+Mx1i0UVB
+ZacImXjg1IsSC38x5YquqNQN2GFNZTrINb0IVGQr0vEmWkvO+ztA7U/zhqT+Kgl
SnEna2lErniQSju01A3hcA+Es0WOK9iiKsy06SOx8X8730N7l/UAGbMVJ9SPk4de
8d2UrWtaHH3J+dpiVFbwc5qOQbGCQcjH0h437fUUSVZzubUJcqeGScHGe8Buho/H
rwYpNX6Fxh1PsWGRW4ZqXhkm8pNKlzCyz8WO/fUHNWDHxQXfyIJ4sDrajFvUSPwg
lzQbfo1NZaWcNjFVIBw/SHDlBypGOzqA5+WmDxR4Q3d/QtHOYNvx4pJywT0zIaf4
ZfC4pWreRPtiPBZ+dyXHnhz/bB7WvFkQ/UA5pzmJV0aXyxj9bvKar6QZsj8c0fmX
MYJ2tpAf6lDqOahacbfxpyKcSgyCLLKPIeAdVspnYvzrdWqIFPEVlF/er2N0vBR9
4b36f7d4DG4Weu7ZqsRNAkwe2FADoEgrW+IUddp61bt14Go8rmm6hU95HuwlNF1A
whkCv4BdCYZ7HYBSrfE8tRs6DY2tAFSiZqGD1/gXHTR/JuTxt49HTr/j9ZGbGMzS
L9caHxEIntE32ofkMr/zOWYaOhv84KpbLRGX2ypKhZ5yKpHsLNKBRNd+AxTWwpCm
wq7zfX0KzM2ajc5Ok+8TD6ub0Ig6OGbNR6wDFJYF0lh5PQuy21ABIM3mSmtcmx1L
448lUz0g/MLoop6rQEYfq8IziZU5XektzsIehoxWx/FSlkQTCtZ0kzPcd5awucWG
qQ8yDWpnLPRlSaUKwKfi1ruSlMsgvBkjUMhhxUfWIUHao7m0oTeI01kt6Tp2NwGN
zCrKnEGbIqiNmVtr+77pOOh96CZn17hfrpNn0JIcU8TrLeXMPPFIyMKL5bs9cuX5
JqMf76jNiSR/9Qry0VkjKS/Y8V2C5xA7FiDMefmBAMR17S1kCIrQWbKpwgO4fiDP
S6akcu3AKWbiqpiyrdPvc0Ihm754DVqpHbW7F2GvWNywNM3g9rdxbp4G9Q8eC3ya
R678xgTgYQJJxyM0xic0KQPyYEiim8D32bZA9Rwk5EVzeogsfd4Lu0pBaW5gRhM6
Vtd8meZvQW35vWc33x7QiBDdg6IJ1vhXEPr6VsCQLd0NvuS/x2sz8qWbZNINOwhj
GFHVQshItTUEXKMXqJJYT3qALBLws5DS3COCGkiE2gxKEUzwAjAa7G/M/+CUBzjJ
y2CV0KWgQvbpfC0+v0lW6hQbOQfiSVccHO8KIZlkKK8BF3fA3zDeQxlO6PDKq4BN
kJv1i08PZU8/MwMdXmcyqs/DxsKi3wEIAngCWHZv7shRzVQNVQDuexEQXMcRLT5j
RPfmPaUEWc66S17o/9kRTG6eXzq9JE0ed1Sb0CchQJy/ji4WYVayREXW/YdyYrlt
yteIhJF0mRc2wvL8q4+DhnPHfRA6UaHCklEXp9mKKJqDjAc5lsLMJoL1lDDKHRki
KFgfzsBE9mkcpy523vn8RMnXv/5AH8TwhG0dMOlkvjyxhnc/DrStynjiktX/E4Ge
H0hbQ8TzioADcxPXkoIyMmySlkvMmWZNXUNyworLbxCVOLpZlN00gwStQQzz4ftE
EMsNdPNfsdij5lDOx9zY9TjD8cvW+LloEoM7UdIYKAWK0gaRthrYR2GoTM8hC4kO
ZEZbO/SaE32ODxw+XTodqzlYd5VFwwgVbZ2cepOEPY0Kzn9Dc4YnfXl04BME0/bc
CyaVCHV15lcVWJPKQo13HDnXi7aF0ae6+2fQt1ov6mzpafPoVcz5QIBKuRHalyXU
U4G7R0Ika6dbFJdj8PaEk/BcIJVKQCzxi1wXt2RCBL3Cs1g99znucbYLqIiV+aLv
+PBNIulwK+trXjuylS67Rq+tOXT5yy1pIBpwc3H4mgDe8gwqBnddvjJlC/lXGKBo
jsl2q4EsW38htiSuW9mMg4981r3ELV1CZy+zL4kjuvwjl1K8xuS7cQ5c5CxGGGLn
UHyHoAtJFx8lWw1caz96CoPloJMHK4B4Smhk/D2E0BCpqMZeAZjauk6cPbSKbZAr
fafL39sdjstPVJdH6nCa2Ed9smXrwuSYRJvxHWyR17csXK85NnAPtOIQjU3E4J4E
ApW5ChWdJMbinoPFxrwAnhwq8CP2kFgfskH/FWFFjTFOHht8zdy939p4ak+Dfw1o
7tJSM5jtMwR4XuXAvyTbWpIEODj9weID98igjFd1L/L2M8CCKgOp+RfEyBpF3KPm
n4+9qOtNwGDXGyMmv+iVvpoW1djXmIB1G6/mUWNnU1R8u7xI454YDnGkTCQibdX3
cFAQMlai7eL0p7kA9J0Zzw3GS/T9iaqSDUNgoxN1TifSEAYr6Z6Un9uQUvWBk8O8
ceC3XpJ2+XmGx5A91FVll8MCBUkXI1+skFIHywZzxdfCu2dxIxtCAOuC2etYvDGS
dNq3n7aj2UXiISa8Xs119LCY7nepjTREgQ42E3qTLByv+K3yTWOd5Y4xVaDMP4dL
mZ8q77z+F/Ua7jCo2QkZWyL0ZpWEFOsYlxprGa3Us58E3eOebOrfwgTTicoZzEJo
r6AHqtZWrZhBCEl/rcpBnUmaBi2ITAZc/3KHdRZLfqyITdltbrzFTESbST/Kubrh
4C1WPCVWER6+pPXt0odQNLVRR4qodesaxD3cxe7hboDhCGup+si6S+oQbNLIdNZj
y58ViDhjDuXkA7Ylp+X9T6F78oK2HjVGBBBbUZKl77FIlRRk1jdmA66nnnocdifg
h1ug/gU73SNArzESpuehmOAO0WOivoHBAAxAAzpEzxYC7Vyib0+D6OLUxHXnTgyn
KLkaKnfvRpQsi30s5etB9Upj3W+tzzBT05UX2hyEfrMW2kF6QmrmLkvW015jhBhr
lBADXuWyY79mexjRe4R37NURvTACOfIXqsFgj09ZyArrhaq1njg94DU+0TzlGP6z
AFQL7GJrOGOCznXSU/TO0UBNXl4eNtZA0ScnEQwAu0SUcnmbLLQOViJhWBE7Yo8+
CfVu3/LI6f8p9nK8MXwJZD2rk/gkcDLjYUf8/l+Vqpjf4R/Jh6SUkaqvgSTIwuoz
9mSE5CuGi5sHlHDT0SXflOfTwm6hqTgiGbmAF1Be0t6IqubFdkV40drjgsqD9xeJ
2CZdT9Cnn1vmKu7nvhv2NgZvfw1avKV2IEzhtkQRpEyUXh77LKhQVo2FOPD7SbIA
69nmnE88ToTtIRzXBJtnLPu33swVKgP2dV8C93xrYjYzMpCr8WuDE9eMQW2YZNPx
4jxwlYDN5ci0Po0I+VDAl4CPubC6Y+0ujyB9XtVh9R4sXTPuhnFovp4jQUM2zFbM
Zr2koUVr6aJ/GpRF4/YT9PPlfXRkzuo55opkYW1RLv/EkfreOA2BDRd94/rCSQSg
YO/3CoRVwnraaRIJkGdg/Xmku9OvxY5pROSsGEScOUj06X6rfmMWBMnP9BAUKMrW
oUpZXENdk3Q8S6wt8aiSSndI5qQKkCyPiDLNQSSGePJtkjcTO70tERkX2ZHMNBPK
yB2OY4cmD+uJwkfLv8H4l0cpt7jKIvdKL2dciQmv4BamkJkSNV0ioCJ3iYt+KX5u
Lkom03AwS9M7h4QxcR/XwgagTw1ei3Ndgr75jOcQWxrU9CtzHjKVi0UmWgvoBHL2
dIA0k+2cS9UNdSVTBHzDFw28X1sG04DcplwVM8d1fjS6g6Wc8odLj2LGXlx5N5Qi
AK3I+N2IxXJIfW4M+XcLf9TL5sqfCYvel1iSKPk4sgQC+Z52taTp37H+PQng78sS
nnoVAQfpcrLXJMCL0VmMRdwqVfd5UM+65E811hDYdX0fDQyJ8bWIBGzSeSuV3s/f
MIKaub6NdhTdaZxts2v2j+GBZ93JTm/PjWsu+57Ck2l3EVswyUej1pP7HjLtZOdT
BWMry0prQc+OYG55nc/Lv+7s1nnih7/2oPARpUwj4CQHG0wYcMyhv68RM+JHrSFg
4724peAHUqnNDlPNrlQ6ppKI3Qqt0HejcN3gZNBLYy5AZIKO8StZ1+KQ+KadIQXd
j/wLnaGP18mh5TdlTaN3WLNIEC60opClx79Qi/ld6DpGl8wSlfIgQlskIq4emzJG
1/ycNIIqW0ERmXpa8ArCxTfIDVmmqBCe2OfTV4ywpnvFZgDvuDLzwRbjiARbwZP9
5wuTFTFhzFlDgdoELsBPWHvBjNf0S+69HMDI8qft8CdIeIJ+txaDzHCJm/dK1vIG
bwNMLZBTfDC0oeNhb4sbOEKwYsqND7fL154W6xjFyNgSb6S8rBF0ZBgUKAT9IpUL
6z2+9ZHyOAQ53BEHyKk2vILMccynJ4bG/Nx7EO2CNhGVwEgkP8b3yWzx4Egh80gc
oe9C97eoQFMyxmte36zYdXwnpMQezgi5p8wSaJlc6FcX4FGt+h9i8znx0qWUf4mg
LowqIUL4D94cR1Yl14z4RnAZmVzDQPcNXOATnZEUFY0xpC7kCywOb0kwoNlyMpU5
wDLc4vUFXIR4v740lmf7ELBYUSgDpRxKROeGPeGvVrbXAq3laOX6nPQsRX78AsVW
KSW+q702+Sb5EAl74s8lq+ubfmv02nnAyZMK5OdEYTlUeFGkxlDH4PVdf8j4Nsgf
poD5LZvsW0Ql5euTt+CTLgodSk3hMb/LW+btjFiUnFrUQRmcM2yrVs1LQP8JOKjI
SAZSB/i49FgtMLm71m9oIRrFpHUkr9RelDD/J+6d9aBkugSsrAsgi82cQGVPTzTP
Yp16nk5edGooIQbLzwxkr18/J5t5isEqyHiZaSsr9iFX4iDVBN23cYx8qzBVyG13
glzvnh2BbBBVXpPX99oBjdBtDtCIzO4ZdqJPr44VQK0JXpGuYKWj9WKqHdICOtzM
gqDDOCW3zfwFWuGdqJCUu3KJNkIIfqTHdwTZziIXIUle8kLjYSDyc8dDPV/QsLL+
1ILEerMW0t6N9tWR/1nubIMkk3HTxEubI6e48ywidTNCQVfStFpM7aqe6m0vi3Dw
Fxt9B8bVWctwPHnYQ/U1DH14efSnytTHjb4LjJ33ai3EHrLc3co6iOmhUQ0PRuMb
2gW/cO+Tj/S+pqI27oSLr8COIKBZFuv8kgFV7h+9Pwk3P3t3vk7Dg0BfjoteaWUi
M8MWUG7o2gGn5AC8MjTJ3LbM/JojX64tCaY+rTawi9rWT+/Yw4qy6zCF9zYxrwjH
f9L+4T549RNcVlMP7WNpGKCq8kZrCmzPk4203NQpY0lq5RHu7J0d+onbngFZXi59
U7pcD58pJCNdKvGxoSrFUZiy25fJZeuGqFB95f0rOT1YIJlrdfrluzgqkCQHEbxl
FyFrAVPBtnF7zoe9yq5Sn9lRB+Vy3nobimQKuYvvTfJ4uWdYcR2A0rmNUNA29zrE
ks9dCsyVZl2OUCe2L6O0EKgWC7vfkV77YTSzpcdDUV5DPebot2+FjDpRUHxnH2Lb
vce0v5jvin6NgJk7q8kJxSiKdtI2oV4MjCZ7tIgYRtlUWTvTpwME50d0fS1E6VJ/
63cXPxasZAlTUm7MQ7S2Kf8guI9dbJNNQD/HR7YXprkq5eJoqVRT64tXTW9uUAFV
n+qdqQVw/dOTabdR9fbfmlb43c6y7dv/QzGef/Q3sL3yfIvj93oJQCd0mZ7UdjkK
w/TNk4P/i3zJMd/rp/tuxswhIIxIc80R8FJFwGZuu9BI4TajhIz+FFmcbgi19Ipw
F7JIiWZ/bhFxGkePuC1dwCiFaHxM2xoohUBuyZH9/idN1cdpuvhlu1XA6yQ8vrSk
MvG7UjZUHU9Pqy5GTvsfXnpfoxu5ndVuq4QRWyBfWS3QHY/4Ie8x8ICDpdFA8XrW
YZy93Z/6Zednb2VFelN7Nc5+CxasL3oyjpMPOMznGk9vNNs0ySmdhr28L7yItSey
pdpzOshP9uMZ+9ihQ28luUEH8u4t0VpMN/7ZxbbLI7lRKufgHk/+2090q35uVDV7
K88SBNG5sBWmViafLCNVcfu2glA2zp5vD8pOwvbP+cU1O3LsanbJNvJSNoJaC3EG
N+t69gf+tXe0I1BvLxOuRxTmmDKAWY9lNWTDnP+fArVf7tB4Io4zfWJQ1JkA5kHc
RNyryf91g561rsZUZskLygZA806bxnydrGGHS+v7LD4=
`protect END_PROTECTED
