`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qr3ec55OItJPGBLu+WnYAZrxz6YWS0FxhYsYwuWwBt93osDrI9BEtDZY5KaB0D9J
gyrSByyZukEPUa6Z+GBZtqiPUN5Z6oo+G8zjfsWcNvBvGPN828EyaXx1GBED/m9y
oLaQTYYoizVVmKLiUQC4KzPSWwY6urZi5L9V5EXYKbk1UDaH4ovVcStcqnPuD5RH
iOVbFWhIczZYhj7k9U49CWggDbRrTG2TTXinHsDa/xt9YhH9iZG0P3cI4PvD2T/t
kFRyufIfizMYRVqCACONpGXIJ3g7eXb/VFHSWGc78PeBgoJb9iRztkTfTfOsUK7Y
D7I7kT5AU2KFFd/f2oYzvV6nrkbRdUpwUPlnZUUUyIbi8MGZ30z9a6qAlvtVPPB0
xspGK/4u67+fdjaG7s9/hyHmZdXT3K0aY4NXVvh6rGfWJcTXzpf6g0GIO4zE0yz9
YS08yEqkpbCcgBgnrWTeDg==
`protect END_PROTECTED
