`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V9hx20bkPdke1/BnrXR0kP9JHDj2M7Epo/k94V2fuSW6baCRlLQcyiGczX5+qoLC
pl4wNSt3nQ05NpIptvUU7iAvFvoZ6KkebYzgvixraRLCLu2ii4QPOW2T4ls6vsDa
9+AkKeKbndZpbiuPwxUGqo8pnw2hEtb87YE/4okn4RW8REpyL/Ixzm+DVAoXu9Mo
0809RKyp6nkab7zOjU4l1bIjfhsICMzgpXH1hLd8fJycgMII+FdxuuC0+++gJ/cT
JnOAdCdoSn1JioW10wrghhVQU6y/kjf/Egbs3Ugqp64oOVlYFad8el3QDfMCDZZi
JDUy+e+tf8Si6RAfjfEwDksENgP2890rK3DSKGt8GCQl7LP6J7WYfiKFpBFx/oXx
MpLsG0pu5fDcj9uPEBo/W8Lz6+RCrRScm8bb1C4GpjO7U5XzK8pYpi0mHmjoPTyS
lV0eNSBiWcMW7YxH1+TDXuJXlxFW/MFskYU0zcAyLyOH5snQwJA3U7B04aEHLppq
AGUaa7vjDYL4s9Dv8Cs5VyrNRPyXbZOPv4BTm7YhAdbEaIWgx+QuKvo3Tx2iezW7
2EWVCiq1QsUX2kUCkIUtNJz7J52CnQmgu/o2DjMiQp2RgZusfKuNvZRsOK1xSeLL
meB4E1K0GcGPisl0zdd9cZj5YCKU+BhAheAyZ1NMuDqvdJFPd6c5BdJXSzmSWASH
JbYnXbmgv4Sum/+Ze2I+KTEfi4uFIyttJlRUb8hT6mUZLignMhHRpHMXfnDCXftT
BJ96spWvO1GDmjOtJZOXl4kA6oTfIIVB2gmErcqX1vJIelXMqgHMYMca3BVAImwe
T9Gpz6Q/gKmXWCyacb//6MIOrjpkrmyuQoP802pB5F3aDj5aO2TjBiisGRhzGew2
`protect END_PROTECTED
