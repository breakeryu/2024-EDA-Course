`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50wPRh6XW8CboO1uMSqRvzC+G0omgpx2HKh866cepPuuDtJ3nmhMfuFD6+qTmLIt
8DQalk/dOBtZGIFHhqCCGUN/OTR2Tz7/hU6ermENkq4uVWd+E0bVH7j/kTnpflaO
kRyXtr7fGfmuQ/FIJCOiGq6rZGW0F6IuYygAjqNv9HhlYxfr68O0ySPyQFu25X+H
RXxOHgUbRNb0j2rp9+Tx4pDex+C8dp8KSKBdgAhZXztJta373jYqcJadT69dtuv1
+anWy4Fvfkv1AuM3H8Ll76F4P8YoaFJAAtL/02tN/ITE1evWRyDTXq+EeUZ/NXwP
cFA6WTielU5r1sj+PTH8axYyuPfnw6lM3SAEz1MztTsv0hVivuD+Xzu8/xfOkPoe
whcxL16lgNsyIZSW6fkXIoZ/viK7/qHsAfE48CRWzZwKuGFjLrvwyZokOEvg+mcZ
vOoC7spZbEncQRmO+qPXTxz6+xX13wpJi1tjeg3m+jt+X0hVXr+g5bzcKJpxAspb
F44pXzTnrLp9lOYVxiL+4nNWpym9YIULS9FdOBbBcehFWw1a9VclpiLH7WCvwJkj
lyg5FZWVvC8vbsZxyUJnJPah8eSmBGlBov6kvODmiN+rI2X77u9rOz3g0tFru9d/
Y8IxoPQN0Wp44YLtMG9id9DMgdfr/CN6uokMMnV00jCTm5r72WK0uv4c3hIdpBai
FoQ9kxBaMjRv7i6StPoTiwYFqI1u967auXeM/+8Vo0LN/U8VOrTkjPEDALc6gKgp
hBrYZMwjvkxhR+I0x0MOkVwX7M22MkTQYBZXuMypNfn2nKUM06GogtTqPBYntxFR
eP8N+76DtplLzJ3Q11v57Wu8HyZiOjD7TbSAVnjrohcEOQ2U8B32IYASSRU/PBIZ
/zgFHL1Q/r6BcfAHli8hXdhUVXud+SjxNTOF+iviEoT+6bXmvL4uAP5y2jqtCAwp
8Wwi2cZ5Np434oxgbQ/CaHYOBEXH0xbOBN19gWmHOzL9s5FgBdUVdTgN1WWJYjGt
vyAttxoeWqyVmp1V9WCqUV1Q9NHHXMrsmShrZrLiW/rYCxOjVjtAOkhA7jO6ZMQa
`protect END_PROTECTED
