`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGH+IL5xEtn1jPXhAVi6bk5FrTnT1Z7Qq8R2pXN4CGoVJ89MfhTddfi4D8LFaPz/
BcTFWASd9mQh10NAdrRld9O3CynL1wfYAyOzpOcZv0ONltId7nTmNpr+YsokHaJT
vd6XG/ni2f0xxFKViqRdQ5grcu/gY63Ia5ehK5mlPLwiir05X3SBGPXWtsfadlwC
AJoXcr0u80TEzslzswt5QyxPV7q2Q9ftdeBplYLaXTrtwmb+JAswExF8vIVP/QDM
ZnBuZjVQHbGTbbd/r7EM+H7cmBA+5elL1GUS/iE/IjIIUTQ8buGTlMvr6kaCEQkq
O4VgwttVFoRjLs2l8eDssQQi315gewbppIO2Co5+18mxpgSv3I0FpOV7ULKCnQT0
x3xnAOtkadbFGqvs7zrMI3PI0k8CVpgofR7zPKy+wd+v7QLl/S8EbLZQ2VTlRvxr
AA5t86a4uvRqhPuZlFJYz8Qz27uBNPDHvmi77ZMc3ywMsDG7pyXkSkR4AxpwyDBR
HMuyi4CjVRO0ou/CkU4YuyZNpD1QMDOjE7+/vUa4QWzsZ/S31yjkzUluKpHB7Dqs
xUExQEbktT8Nw3rhVDjZlMXFOx25z0wa0rK07k7rUOjfSHLKaG65bMsBQg80hl8t
zCphny9jVzk7t99N/LNLnbZfKT9b+ImM0l/oA4XPG3gg2oKcKZvZWlY4RPkpcRyS
CUeaHYgMJSwrBIJm5fsgJcsk1mwKHieOhBj1BiaH+69Ym1hpfoe2qWTsW+blDbu0
7bFYYufljCv8d1LsPoNxFApT8El1qCAmJvdYyJtHSbyqGiOL12emT0V8GgUBPKBY
TZhTwlrYocMyWJeXpkrnFSyUe9QDW+dUgGeuUP+j/HPPitR3aL0yZD8dFIVVYYBA
05sT0hi/rVgW+qg+e0ORIR9PKGqi8xXdBE1s9TUCM5/pCzRNIiN70XZjaIugBHuc
oaHx6aGdAmwLi6fBUk51iVFGs1RmfaJA0m0O/KGzh6tGhBK52ns63Ey5Cy/49J/q
oh7ztRk55HUTXPjjJFe7Xj8KUHXLUVrEDwpZ9Cm3JbJiFVlKJGxAoaRdPOYysKnA
CjWOcBEE/wSdd17x4Z2G9VR4vs8YpooaaGwuPBeeoiZvzwT1HmcfbB/dqHQ9GeOy
wbZ1+Kw8JvBIEMGcoNqEaYnfk0wZg+ynPZvH40tzH8PQM00b5Z3iYQc/lRL/X/aw
8c/8QfHOw9SpAqceYVnPIYKFtVt6KrFxSFjphfsb85lGGaDDckwGrhYTHZlAarZ8
VDV6/mppSdsqb7+jUZq5E9gkXFvOpluYDoN+Tuwy/MpBwwUMylKfEl9w8gLbpaiq
9WcRGhIE+0wdVW5QnyjJlnCPGHF4RRKAS+mJ5GaqMMmPDWaOf4E3OoG2XHYN3U4H
sgzX/lR0ahpOfidHowGvJ/CIB976l830f+4032MpyO+tKFjJ/jRukSV70+Tm6oo9
80FXvgLVC5G4r3IvcANkVsB7YwSncrau18wVfBO/DFEHpuGkImMeT1oZAnI2azyB
a8/8ha4glJNHgqml6JZ6BEwb2Ot0MtfnOt+E9KKwBvR0j1Iq06u5BQ/p/yecAMWC
eQQRm/7kdDH50XXA+s4No+Ext5XseRqktjNVQtkJ5XyghNQCdD1JPVMWk1YvZYwj
HDce5rmxonbBEW8EmYOHIHkOqCBC0G1c5sLBUwjlER6vdDiSyIbJ/PLqdWTp9jD2
mDrALGGoAGPtW/UQGSEOXoVWrwJQuSpV02A8Y9UIBI32bjfbgXhs+++qDP4XjWKC
Ljrrvy6YGNRirYTn/FHAXBO+5OR6t0J7vYiDg4SYybToYzg7wD0fRBiw3wDE86Gq
9h9txRD5rZoPf5y0nVXHteTA8afRQMudzDpCA8PgiJSMrYArHtzhrvIlaPqAXE/X
+BNp253CHcJCHGr3CxX8DGJOEwkUHGJRrmg78R+MzcrIJRaEHtcgInyTAjlGKNP3
iCelzpcxfTwbLjgI3cB9MLDFAJ8avTg9mXmvLlP9bFEKa9DqC9LxLxQ5fSCBbLrs
5np2tU1V0N814sS62BSPjm8QYe1A9wi5x2JWT9ptN7yLcguyYVxqSE454N1MnY/d
eiLZ5chv2m9fYvahiFgrE5PmfI4ZP8sTqrAXR7ZQ21p5E2+7Ye62Ly6G9DQik0jE
DBWcIAdDFBybPVJiWbHFluuv4Y+r7zXLCp++j4wZXrDxu7zIzR7vr4Wu5dIVIj8X
BwbNX4jboXQElXORw6nD9FHwadf08QxRknQYCOOBY1+qnyYYUObmhyXsZpNE/d6x
+jfF0N8/2cjysIvHcwEwEBXVRliXoqUHSiLteoXifkKffOank6Gi0i93B84Su4wt
okaU3nxuKLqP0+pVJ788fX6SSEG4jnjx3Mw8MPUfJpZPEYQxhk855QJrKBzh8Jea
n51vp80aaI8M/k5cQP6DLSbiUwnU5VitHv4AVNaHq3vJ29SnFceVF26qn5MKyqvs
rybbBMtAS6/Ji/X13XLnKRn3zzphthpyPsQddKHXY/tSSJiVoDBYfQSv1RCZvUJM
EpO59eKJZg5ZzQ8ZcVFuH7qKB5KuQrRT1Oicuk1lhD3kNuezlGjVY2CvE9osMp4t
4Wn7Ef164dT+xRucv8/CsZ4IMvQFTkb2pXdOHXl4WaN5+9eydB2RCpfJmB/eY1uK
qU36MVG8GfdmRmyGMd86s/7QMDyI/stTjW8gDCQEoPSZ4ZsKZJVAz1n25qeMuR+4
VuXWLsyZlewy4VfXRfPEl1OoTnEXIZ/Ivx7gEMREmlldX1ooZjoyYbFAwwmGC1Sz
chGCZucOrUBbkQ2/dFeYaoznni+IqB9M7nOv8sIJvhVlCEqFy4us01tewQ3p4ro5
IwIhyJdMbmrLSrrQC0oLzK3t8KQ9c8VGyQrYFQSsbLtDr5H0MzV3KyGCyC741YxA
j0558xMsWaUD4lL8HpHGPb2yiGIppnH8U4S9AaJjKkGBQUvk5H+b8cg/Cmf0Mj9f
FNxDiPP+9TSrgiie5F2NzBS/OF40sLQ2+uzC4WOQJnQkZvqBI0i6c28hxl2KM9A3
6e7d6jzqy9gwLRd8o89H4PTVT7n3A1xIRJFdUp4fdmO6ehBn7Y0bif45kDHnbHSt
ueP5k2iTQzeoSWwL5noX63gYRMNuVCQcy7QNGTWhdmXo60bCP5YKzuoCbgueIo0r
was/9cpN2h/khUbRjW/oqQDuVhm9yAHGB3sRd0U/OOZRJOtCcaxgc2CwN8I2JvhV
6rdjJMgiRDC7yQ+V0ePRV3FEWXBCeL9iDJQUXLaw9lo+srL5Mllxn7v6up5Ir5MO
9hfjNIAsu6JO8sFpi+YN1W/KvjYDYbx1xk7XIfCgdaSiLAKr+tYXXnZ7N+ELzvb7
KnhcZir/EtXVEL+9GsakOP4ahLPDlbKBddu363YfCMtXN33KBQ7MwF42oIG4EZb7
hPM6B4U20uZbyMNvnhCX7YSykvwtBb+W1bieaF9CoyNuXBGkTEBujCYhoyM+g8Gp
oJobL/gi6pVJyx9KGHxdFUuqx072hMkZAHnS0l8pMMMwqLolErgLNygFrSQf0GNk
+fR7AROnzd8Qv0imlD2fxuy24DhaCxcpLup5wIZ23ulqj0q7b6J70y0BTviPWfJZ
mJd+KJLR2nZZn/Hb6BWJNOrfYz9yR/nEbieZAN7JFEcMJF7T5gKLC1aU0+WBFqDk
1VeXPrMp4OZ+XmkQy29UiaLNiDZ6hONGYTC5ibq7s5fdHUG4s12WxYSQM1rDqKt2
qTRxvWLeaF5ppjxUqTkEb5ENoZvT0G6S64+58bquMSiXq/KjUeteEXObHOUKBotR
HiS5Vqv7vX8Rm1OVswbYcIR5xha0w8iZKq/2og3nnnZ8q7QLinw0y1rCbt8v4zVf
0uX1vLgeq7qvQlDTros1ySfDKTBFiilENd+13S1U/f9xGaSchxAiheTu0XdD7F83
rIlzA4hldbCDWXb1p6IXq+p/8EgAQFuvl6+9QDmQxzgOViIXHWSiefcgu5XB/kKl
34asUNK6HRaszlxo47uRVz7UFbhobyfxhbobOCUVcjLU2jG5MExAOXLZDWJoxey3
XCl36SkcuzT3P5J/MfBhQ0GMGpuYblH1UXT+dG9jhIfkcUGH9w+GCRJ17AQb5hy7
no1j6GWmaFsKFh5UL6z73ipC1v8JzJHTsYPljrpQUIWOfuGKT91lDT1BVXnUXLrq
DEgv4LFSe5xhOJovAG+/HO/4V3xhDNOM2BNOWMC0tCZXY/qj42arFXeQQvpOf1+z
UXLvDXLKEDuAayO+7Q5gCpGTC2XB152cukVrhEa+kudUZo0HC+pJ5EsI4bN9YChq
PzWI5zRkuP8776G4kZpgVuP1fQ4+xXp70ITwZv/1ZtL8KRRfUISvJs09A9UGyJjc
Y96p+fBeX2b+T6Ir7TqitINXvSij0/JH8TXN+OtxucQf2t2hXOZzomSuM2IZCfsP
mgsuiAANMfhx3JMO9cJotcrLYSyAXL6QhAyaMJoKdbxQL3J1Xjzh8+feBkNWSEOu
ySn6Ed/ueRS0gpwi/Tnjjnxeftu8HYP8/KNoLhSQQcpYtQkfoH0X8YunPXrvDOMl
AL2UQPCd0uAd1oTkm7RRcXfBr7HKWHm7Iv48ZoIOSegCNFkRa/2oEcrimvQDR8lH
gnG/544YyNElpOxTNC+XibjM/jX1IwXrSj7HzP2WkayGwpdaf0tJrCXDFe54mWro
rxndviw46REsBtc9enzcabatKlgpcSJF3B+avydKKujnamPK5LDjIa0SMyTPP2hX
WRtnm9Nhp0aH7Ihe0C6LIKQMvk98enFXbUE759vq6iwfZ1jMCO6fr/qss+z1GyQa
wLvSE8l+zjqKreQcrLpdk8JOkSF20+CaPv2SXCP8HspW9v0QT80w4/HicGNuawIz
TWERjKqeaV86tKxjTkRSrZhJSOyQ8kJXveDh54Txk0txvxiWzHkqFfd8C/TGuAR/
yIe5C8hcFJAeBnfAVGTGvhDBZFD4OZNZ6WWA8rJyaHijpKzEFdyZzjthBvFsaSC6
GqbZexDaRjqzYNiVgewsBLzQaIJ5GuvsHtipGw7L91rifNCyqTYvDYFGgErVpr3y
C9tRTj5x6xadtuDiQ2RiSWqdEoVwo88htpbgcBQyXYSaGSa3o3PDpDkCXei6sWeI
BbZ0/1aOA2TJLj685eQLUnFE1MhMXM1mtVJv/AXpyfiM+VUq/rrafArMsMbbbeCG
rK3N5Xd+Ep4Phw6G0W1EHBHxzQ+Fc78QbmtQtjiZ/sM/RTjdDk1zQYX9E6YEVksD
A/TvkeymMDL1BCjH8B8QJfPT4jB7kHchyrrKsl0yMyzQZJl0zyIUEHhD3/jn33m0
qomKvDGpnkiaEzESDO1jYNabbbjDxXFKKH/DddqUkUUugmJANnfWDo7dDqwexVlC
FovzL/hBF+R26JI4An5dKKJ5Qdtu7VrH52wamD0rC9yHs0u6X6CJROrE2BXneQci
3KA3+J/nNMzXiURPl3ZI+AOJXxUa0LtcoUEfSzSpW/+cUr2QQu1M31CUbEjYvEsh
Kyp78n9mT/lPhleTia7IaNpmErI27h5hDtOd2FLGddxD0QSwwEwp5D8Q+y7qXC4I
E2JSaYstGKW17iXnW5NSLturOZCDhAVZPaqIaAXOrueLraqoG0WFbBQ1Trxs8rck
G7L3SillU43b64FqkCi53nD00S1ngV0DyY8EFdq+en4V9CiZeAlSIGkFzA1bwm8o
difsMFYm1pvb/dygeT8LS/c6syO+IerB12v6zbC1TeYBucyXBESp50vuTPIDTuMD
9XtUt86e5bDLV3BtRnaBRAN9OriGOWAbEIdpGD3HPsoy2INPw5qksEl6csPRSbo4
JLv2plxcqLovm65C/hM56ZZoe1XTX1Bt7S/HQiSvNr569okr2eWEXGjXovUnQ94C
W/ffUU6u9CdXhjUtatetB7GHh78uSyy+6jSKu4qzz9Ekt74cMbGMCoGh9CUG+i9O
pR/NcWtQfeMHU7O+8FntwNVMX2n02tOaJ4N/j1padypNv0FS4GQfFtwLyBLJ744M
TYL4sl8wsKe2SJOsYjElCfTPpWcJK17afoMvHAL8MIN0Kd8RbbQgV0PeeEXQ9Ntx
afCdqkkTTWrgDimenmPp0wFNw9CSoyP63KQngDfSyBYGVtqRt63+ivmcsWMQe8Qm
6klnDDKQsxFx0W0HG/qzUvlw2NZE/nfl+lc3UubGTQ5WGZ9tKlKISRplYxWZ8U+M
TM/z9TlkdF82Bub5qog7LFzlqqGderzRrb5RA5zO3kXCYfyHBC+6FWqT1Fe8gMHD
fix+4e48BJJ86LYAmVtuj9FbIpYWmeTdZLphXQgqJKCdpVFv6rdeT4dJZ+36uyvy
FrG1fVi6gag48ER7FfXO8bCB3BN6HgvDYEGspHGlJHILz1GFwNq2J9k2M4aYygPB
26lQZmSutmYYrxAu43osPlIUcCuLZpuVnQQP4xhERoDZ1QIXbtd4NMAT7v39+Lkl
s22GU7DibHfGywdbLyHbu5pSd8mRjIbvkFz9AgVI/uLRL2skMx8J1DbBjoeQaNUE
dnrOPXJw40WBfqOYUTJD+IKAG2ZIi8/R61pMJ3b0I5RytVCe7KOVcGXfbyrF+ghD
aZX9jYBgo4MDUyoElcE9P+SP679C1Lo69P2qaWykDqPoNpwWC/tWmK4vNBZT6/2G
VmcTITt65L4M3VPxD+Q4yr4qQwio4+wQ/PJdcFWzWyvwOQoChT0ipM9aEqnAcp+g
cV+wZlf+o4PH2o6ZhMA0RqTITwEr4QxQj/9Q9GW9BxKBgmhwGOO6j+kC9q+LsIA2
86lA5iP6UONUx5wb11SOVElcMWglTpdPhif+/DHLa06hr0casy0j+u+QBr908Lov
ZoRkJT+RLkK49vabcOqSLHX3Fjv01XVTywwkeypogKbQtXnhG9v48h4D4ZopP79v
0BY1VYB+XpXbuC5jGi4/8t/S+CblTYRqCHil+vC2whRxmwhZ+Yz2Hofgvw8Ykgob
a1JOSBGiOM7fWcjBxiEyo/RXvyZI7jZP6tuIR91nurL8gIiDlsCpPDyZmTYzDWwd
a0DU/snN1YPDr/3JKzf6Q3CP2Ok/dysGAToRdJjonAS/QgpBv2AHl1MH8Ssxlr5w
W+JXVKXw2no4cNymOYzslltOxlMEdnrB0OvcvgAJ9eJE23JlbarT/pv/i/34d/JO
ld65pDk/SItEcZlSIQWjvfEfq0Jt64FvikFOgoXRDoO3NQtemc4BwwQo5AZ7CeHG
JRW2fwaY1ycySKSUwNc2sQAz2APGBuZfB9xPyMHisRwzHRsUI5ojTC9bWd0iUIGf
33xaamwGQWCT6xuOYAsvxDhq67RnSfUQ2wqdJSfXbHPze4q5Cdo2GCX7pM+h4dYK
WAK7T2cWQkwevONwSCLIxFeYKjfruyPUiqMe5I780eKiFJKbRwZfc0sMOYxyZ4JP
dYAurV5HtAsXQj7lUwTMO4HjTLXQnaNV5QEecSPRjCpBcdpApwZuKv5FsELrI2/L
gIYdO5TStP8JyjJLLRqWTFUfMHqEgssBp7pt67ojY2P/HA8RNPJpOY1nmyez1bna
EvfGio1I3zmoiC/XRfytdz/quLLtqeGp3wnCRmqsbL5YFjpIxO9E6N8PfldCjciB
vWpz9cHP+mZVSPrxQG2AOBCNr+Ip6VwMg7Ub5oW+mh72pqMmY7AIqoO7wbn/d//I
q2Ch0Dv5y66iGf9GPzw/zT9ikcd5EcZFeh9QndQHkOmZXDY0UPAXimZlNdFeipdA
PBkcDlg2Dk+JTlDXFNyj6aa/Z1Fadqf8NzEWds8/j8sHRdlsXGpuTgrnqS1lwZno
XWJs61Fea/2B4DnSg8e3bBLoeDbo54Ooa75Yoq8dBXXYLRLZ3KkdmVzbJm2Qa/KU
7u8tXbmSD1Dk4F+OOany/hDk3TMMcEn1VWQVvbfAtcBf/jh0tSY9qt1OZK6qYjKE
iGtb8eTGDwduC6QQSd9Hx2nqqOBa+u434v9xkNQdt+SC9zu7HM8CVotEmuKAAnDm
2MIcjfXN2JqNU/ojFqVvI+F0UzGsdeoUI9drcRFmIH4FZaW/VTNofbLRaJwwXlrv
kUtW3RWP/y8xTLSJVCiX7FVvSHpyWvey/Xg6lQIVFXRE/NreQ2yczD4uU+HKZbZ4
KiYciaii1pch3qU1KHgOgKyQvEQzAUx98RUXiLg/d7qfBB8Kqdo20MbIFDk2gGdM
Hl2nL6E5PuEMBScOD52j3GQrhUpqmxebq6Bkxr5fz6tHcnkqM7yLEergV46GNn05
eaUSD+8YJcu1BDtQ4QPJzLzmCdZexDBwfKocw+uFtNIVEe0uWu6PZ1gic4y5IsBT
1Sta8J/33ynoNT1ImNU8nhl8y6aPgxLCLGYjY2sJdscRRLhHV//OIbBVgAn7T9ZT
DHppBLNlUFmVoAR4LbmkO2Z2woZ5yiHkV3uNOgFnXptHj5kEeQxcbB2M76ymsW+2
wua47+9j3FOc+KXxBcbqPiwYaKcAAa0xelNmaOELcy52YfhSFQD2ZAP6vkY1N4lm
BRnUhld0kqGMfdsvfm7Q292wwiz+aZum0DP/V6NqjhV68/GiXovgK6Txu/0jYCfW
435Va5MJ4A2ESQ02+9D6ywZrLChrqWOiKqPQ2pyeQHWeTs4BlUwuOuBKSku97QgQ
RRVb2S8072xIbp58m5CrpdhP8mEhZT2gV+6+UyTrt5uq5SW4OHTMmy6ezZwgHWKG
YOLd/UxWGrkT/gsF3aSpv7lYoqAJ49ZdbrYIi4TwpAB9r3d8BYlYz5QHBTfMkeKF
oipfMGE9oWgKUXQthOvBRktB0bigJpLFKOp9Ain0BzGhGDhUTb6T4TLrLwbmF7Eg
tH4Ib+uAhjs3Uy0CwnMtdigtiVsjegtktnCgtl44tqq5os3l6tDLTaGXZdAv7wO+
8Pd1UoJKSFD73HvWYkmIl9IFH3xDCmjpfGejEx5cs9oPTclC6j9GVOsnBYYoVwr1
ZwVuictI2A0Ba9iGDGncjsm/4dYkrnYU7covN+j01dcKj0l2gcdePvrR61O9Xfmn
9uk+BM+joHroUXf+oNYcgtdxKtILv6u0YIEt/wCBmVH3/kvHvrSclAvR+ub1TArE
Gi3pKyE/ztLtThgb29i31S5N4488t922UlTzdd1SxMaSOAB4qD7vShWVimKlEjFe
A7ObmTj4xdSw8fnoRfPqvUR+LRuyD10qUhuNf9xq33J4vRHjkJcxDYKfpSkE6mpW
7rmbaBUbXx0MuaUPBIaRJ3K2MfxkaXPoXV6/9ccXphhlU5X9SoKrl4LmjwaJQ4DR
2sqbBIQcx1pXYrCCyiLEdHBsVpLi4feeF09oAwV7MD3AXlFkeZnaJXFtHbg05r0e
+xHAnNax5k3R8fZYbt1jWy68bx67/LQK+H4mVEgkNXg3D9jxXfqUwcmpxrELoCFQ
U/KhhG+emJAJNL81r22UvdFU0pXD8QVFwhQyeuTt4eeCZC3QOx9EEBiyv+VeBP+G
zAzndAEStpNru0dVjo2zyl53yyeTc1hs4uCpUcKzWy1s+beDJtiY+VI0heFGCh+Z
PYHUA+g6nMnhjZR+6CwMAL+i3eI+B7vps9KEd1yiMi+OVqNSLSf8P1zXS+XZUUja
6RYkv9J9h0/ZKav94+L6g/kkzc/55eHzRKkposwFyIydwc6ZCOmFjGqvTb3fxHeR
JqRWvXSQgAnxWPDkGYtolmjHucfOee0of30uob5sXqnjVsnXFsG479jg4ZwlASvh
a8rOaXKi+1OzJi6xIklUMVbia4UiAesUGYCX6u/9ZJUl25Wj8c0h2k5t0Z19LHOk
Xjk1L5miRQ3pbHwMaw3IdebOaXPgkIaI/uIbjUuz9OwB4kYtVXOIIY8ykNy039c0
7SYNXP/Kuv3GEMvDp+i/+SwvSbMxqXsZ0fG4qkJnf+JVkSTqXWRRgYTQiUCWZQfs
nEYtaONwyGroUYq0aCDotVKCyyUS/s1fBu8xl9wJcTxg3VYBY6gDG5g8hdN8PPSb
o4F6Ot70OjbVd20P8HdnF/d6lIRFSeFKP1QZXkIknS8cihQ4RQhSoWFar8zxqYy6
two9o9zcsa7h2JWEC9rsrPfz2O6zD9JqtAuKL0nkF+FOh0yQlKBszTgReWSrfShL
KcjF8TtbXEzDFLt+NfjOlEozE6NwPTXYpDCmfaQY2Bq3tqnF3i3IWdd+XkIL7lq+
SKjKMab5Aw09417ulYz5WdM4yZEhiB3Pcqh8a4wqgFqvu9ZB5nubC+/KAS+DCzgD
qyQIHjR8JgjYOKU7xhZIjvnnVTSYJiU0tLhrumvZ0z+Twm40vX2LaePqk49RxaUZ
j3AMeM3JeaSFo6b4p56AW/Wp6D10AqVPV+KtWrPxeYdYsS3EI2BBduGyThMt1FhY
YxzRUCue4SZdcNJyQ4uzOHdew7KxC6MBQuu/oRZDvY4Gpsgl1geaBBu+X9l/Xmql
wLFVOt2RcYPGpUwS9p3yIBpPE2zD74AW+IEMg/lUZ7zu9dalLvfg6EpaLlje2SLG
eOaucR9memvrDVso185QPEzRDLF9arQiJ0GBObhlWbQNE0Am+mpmzs6hfFirDB27
YlKUz1R3T5joh5OsEmo8Z8MOSc9ULQBnQmEtFeG5ZoJ9D1loW1qroy2ryi7CVig3
rkSoTOStOBWmMxqG46MFrYlvDdKj9N04hvagI0hApSoYrzzH6hLpRZpDrEDh2pT2
Eq9eN9bnQ5T26YoAM2Mww4DNGrZ8L5U1rt9wwIF3k6IiW4O3Ybw3e3u9U9CXdQ3H
w2XG/8n0Pyv0Tca5X1BWYavDqM/N4+VVFe74kzcAa8YibW5z6dvnfUo9gB0y/OGw
Xl/6gKhkCXyp3BKEoa2aVCZ9XAq+EUhlU18E+I9DvpjYiVns3n1ZIK9xtaPCY9t+
QrWwbnhZBizZe5my9J+UAxIXR0rfGimB+sqWBcWEGGJH6mCrgnOIIBiwtE5I/wih
j/kCRMgKy/v7cA7nm4VnehiY/jyj8kQN+T6PzQ66zN+JotPmfDNWkLr7wqtFPv3V
CG6yb0xKkjgfzaGdKNVn8grSnS00VOvp8jM7h9rOg1WnGIbvrM1mmICapHD1fS3M
lHbx0KbFxnG4uOFr4epJeNLs6xf4/kohVl8zqZlUpWQmtPVgP0knk40gpkrMTWMN
lIMPX8gDBHUM7+BQbHBpFlTtw4z//6TOGPlP7Zmk5cVunHurVAurVn9/O+/mw6Dp
AtUBRonRXgYlvQn7RyvrT3cUBtc26+8VDrXUerAsehFLkIHDb2k9Y7CGKujWD3FF
xErNjjTfprnCTG60Ozj11f3SSZggZCZzfuEUss/ErQseo+fj/KF6b/UhGhFc+FOJ
ktK20YplvmrTr8YgS3MYFmQoOxVYUHpgckfjIqfEFwTDJvvjJ04QHCvbEji0COZ4
+fSLNZywyn9izxWgMTCmahOKAWoW5nPWDLDNKTL6bFVvyV0nAk18XXnDTgmSh3cS
9raPi484zVqHyQmXgwgRIWFf/d4a9FXy8Kbo4LuwVS43kWhD9CZEPKSsJ0qf3Y68
GbR+WVZjOL8A03Z8g9fg9xUuWLBxJBgiCNx1LLJdK6g/l6GA+UzTFBHW/RpYNZix
pIqEk/XeQujpozRd7UfI3frz/D/E6xbhe5ZTzAqS6INkQ+QjNbfBXCqwnO0eHN9n
nOCX+paftYp2dicvn9TGD3ovmu889LBlXFpIUsqwuLBGnW3CWF4mBWpeG7zcSspQ
lufzG0U6PHEf9abJ62JfZWVG7GY7+qYcrDw1mmAcLnBNFyPqnyWdH52dyr4TXdWQ
Hh1oyPDM0G+gZD+83x6+lDbdo5CG/J2ee0WQqlfGiKiBvn/da2R+qKluBiPRMiL+
ez/7bZ12QmM7vFWYERZneP1bXkUhsNuth88DjE1Yzc02alEThdlVnIiFQO65qbFb
f9EZ29az/ynyT/XuiDtA0kMnDN7yvjgGUZD2lI/HlKu1lPtKLPZHZ7Fx7Lyzede6
AnUCvXo2cN0LD4KBtURd03NWvC1wZlgDjEF+y0kAX0DnR1kOGvRl2AQh46D7ByL7
Bq0joBn/BNwT4Epq9uHFbK+JFKt0P4U+FWzxSs8hCepsGZ5DyviTcfwwgBmRuBJ0
GtTLEuVO8dMk1CYe3PlU9hilxadoqkZ0VsRdQSk/SrqQzWfQlhJLBgRYaAeBxoID
ZavKL6KEbuf+/fhsOfo/yeAM5tEH0zQJmtsfYjqR0FoPmzl9bqPtmn1sbSKts8me
/e/JAqNpCTZ8Tu7OcyoCpvrgXbbJ7rO67IhDZF79MO+FW9K8VF+/l6u+/CyFZh3J
rKm+T16i9REG/TdETxnJDLyVAzG89FZTeayg4JGeCbv3GxOLVMN/1sMl9uP2XloQ
2cAnCFdf2JMty8lClKsSK/RBKJShuA2wr0uHG6W+EZEjEES8pllWiyRmxEci6GFZ
is04exNJimToC50CYTbkurvYS5b31ZtxDvIfSePzOpm9lgk49ZP1SGReBU4OR/yK
q8yPhFL0fJbSYV5a499uoHkMz9HRt31g4Ukx6UHDiXa+kgDPN2tUALjwfgElBGut
jX13Y6fE5aahgk/7cOCADPExCiPCjTOW7kbqrJDlkObf6L6QkO0dQpYd33HhmuJ9
4QsPvN+VLp0JHHUwHuH+InBR8LT66hUi7SPIbaMEuFTKq4bCG5DQ5xEKM9nXP9yI
23cW583k0elohj1MEBF+9UEe9Nt1oUgRU3B9Ewu3uYGq/KSX7GDa7YFfJFinycUC
H7j14+7v6afWqlf06lxyNJXhT6iSddfGyMJk3qFPFk2giJr6Ytf9nQLjA+A3v/Ix
Ug//oYw51HZFGzctfvSw3tvzdTeTXe973za2uBihaP+biNwPbTkLeQkl32Ze/m2S
fcv2WDkQv4lxaAAiXalW5QfoSlRLXZ5+gOvSXVoXwIv7JMoB+JzXKSecjPVDnYUt
cw2CCASOB+CKOrO3ZSnT5BKLQq+euNT5Z9Z/A2jE0JKYH79lqap0BUzAPLnUFQF5
TFxVB9g0d5ARiNlGmkb9W2oXBNmv5COAOZPhDx0iXmP0gblFjfKs0seCHcrc5F+s
Nv+QS7c2MowDdT2XQCD60ju7reg/F31QnNQwg0ouI0Sx83d180/JuH9U4/SSFsQg
JO0zT9OViEv6B7tdht7CQgRr4lCOY06eAuutI2A0VLo5KELIFdmvPRCf4tVD6ZwZ
1Jp7bZ+VxlCkRnl9nfhDk2YOXrqzJpTP2VTEKGkWfUpAHRVQy4XoGKj8DP9hHNts
n/3tlsJ1gHX8UtPqFWKpItRdekMTSU/W40akb9u5z3pBdEEGdklJ3AvFngTQ2eMB
ySuwTGS1WqWCK87zGA+mmk6jwGfWpSbcwq+b0S2BbtaqYKW1TpPLUuTnZAB5LfOU
XECzr0FGCGpKSPQkCCNSEqtUIU0eThLwJp+ImS8MnI5vep2vHxmQwneomIL5jgiK
CRB6DlRsL3X9OS+GxMWvV6Znn5qaZ8dtkHWYpiqaCa/aCXCk7+/29xVeg7r7TjTX
EilWcwoC/ngjDt9IFoKvhFmJZ9zLJvD5D0c/4mF2Kr9YUfyJkmJpUxoymUqH5+SR
XBlQGqKRwvAoC1by+HgHr3WlYdVUYYGzOv3MvtZ/zv7XYlBwHe678MI+5fi3VkSu
YPnYMZS4NOWMLfFKH9LiPoG4zASDxSpvZiwGOetWsMu+lAgWerkAYV6ghg/iSX5v
e9hu8F2ufuGjOEcq+Lo3r6ijYFwEzkpShnoQS0Dt8d4TT6zR9SgkFz3PeeWQnmIQ
v4XtmP4/0zjAlZxEZRWZtAELiPuecz8xXiLxlURp6iGui8yftWmASXxCpW7ptF31
KbtQO6pa3kaUZNi8y/xLYAs8PfZcJsOiStxgLkOnyFvpHVM/4rPmKO3Y1gZqeRO0
4f0Ssc0VTi1TFDyz7XSyuHcFcTOCSDthqy8YkYQBcTxXqy69Esx1SxWAkk0/MIoc
5xrD3leEfXqN2fkQp7JUHY3Z//2uPmpfCGF5Bss6+S8M2oC8Qh0yzyco9fw9plFy
2xPTXdW/rCpNhpIRvNjjnlPegwD6+VWtSFpDweIFj4g7sTKKXC97H/zwm15Mj9kc
ES4aRR9TKjm00hnx6A1HxJxBlWCVDxR4FXghix3QiHcmdRkRRQBzkoDCOUrXV5lm
rmJAfwyh4EWQuPG0QOiDWEfWtj/NOqKeUvzxiLNfDkwkeQEcvmrW0BAFr3zUyFzt
ZTcZV5qroUb3mAR+JQgLAdSLrMRD2fuzjZMwlcetPAKwSHQUPq8gMAmnwiTHfsjx
O8OIa3r/p8TEJseq7lgKFm7iPvMeBWOme+HK3zUMEIeePDz4gMW4pNbVoDcpz+PL
12Qh7EakHj584GPST9NG6uQ/8gXqHUey7UP+vYLTZ/rAyjejBwy0uhwRUFS4IajU
S57sE7DHLlO+e7F0TNbQGeB40lCDv/puPdzI2bXA7H/9dCRo1a+4TxeV5u8rj96Z
UC4N+SmIIJ3XSqV9aZ1vD23aJGt3zBYJHwXRAZ90z7/3YDCA0JrI5AAoie2viTBI
ep+0aBWAFoIqUhTYz1yHlMw2U2b6Sq4C1tFwE9nfOobb/aLKnnzVfp52knQkGyvU
HHuL1f+eVkKIROxyTV23uj0uM2zsCTjllBJ3yJ2IzlgKLFhlpv2hJVkRc/0VnRrS
Dy3nnGu9LVYh8UZ/SdFstPBxT7FnCIAIzY7OZfPgdp0V5fYrcoDdQ4JAFuIzDQdu
9S3nHeP8VSb7EeZVlfCiyesWId7aAo05eSHnCfVcRU3MxG6kAh9Xg0DYETMTG2a0
HihBUu0x59o0/ZezJqOZVNwad2PY/437KK+0yoLXan3dircLwK+EAQjLbiye4fyJ
yVcMZfKSiEJKwxyk8vlUCB+zhvANxQYTC12pI8gmLI6a19JdFUe630Uez4HpaDe0
bsXDOcvRzcuiFZcZeZr9PiTi5RWfWzOQzf4OzKWNN32DQF2jHqtHoksrKurL+NwI
JVG+9IH6MeqXb5XElomCMoPFhT0Ca04cmsrGmJncm0IQMsboI0P5afATvVuFFUPa
QNp94aOMuMfEWPXvG99jHOZ56GlMrryT0nZYx6k50WpB/fiCDugQSwAr3d5xwfpt
EIYd2F/NuNEbldISdDJU9lVxtKi62t6wDiX0pqmPk+RP9rX2XBUE8UsB13TK9jbH
/435gEDR/vqCGnMMy8CWhZlWM0ExW1Ly2XpuTY30ExiAnhqF+XrnMra8qHsKjIIg
zf01xV1NGbhP6th6XrEy1pZsSb/fdcc4Eo+x28TWeMSwIuKKV3KfQ1DAKSXliRSw
JXYjvrVCg0UvcrN3acll2Kc9hyZW4aW9SKvBjJBA3qvDBTNCmCjXKm6OxYRjRerL
berSU1BLsrsWE6/L1Yzm6Kn2kYvMqoRx1eCLU7TJ00j+/bipd7eNHlaeN0OYDt2G
098Zi7JdVssVPYErwZcC5BmnaKCIjy6My20mOhkreychYkOd8pL+aZ4s3uvjGrTJ
aDUL004JlRQypsfAOCcLnJS3iLzXZyAYipCMtP173TcEM+hMlUi0ls+Yn5lBD5Wd
6O9Hir/qpF4itnWrOayVJD6UCpQzzvmEsLSxbQh0LC4FlE13D+sMF1E3kRk9CWQJ
p9RrBUqOt7hlYw1sSiIFigFLoVOQ/yxxxJnzcG7uBi5JZBf32ZPpS5VGpFfhpLdL
6KX6FNGTu/hzwjuDjajopN22thhdNpoHZx0pVs5esK98KxmMCJDnCOsldXRNZmyZ
jsJ7iDSTLhAMSLWEqGAseVfhsOU0rpXpmofZevnWTmKNT4tfehk8Hi/GkB1qW6dm
tWMJdOu7uDDj9Z/y/QF2KHfv+j8/rtR5sOkh0gIuCpuZZVxk62eOr8DhcHH+7qeq
Z+Hbr1QpX/p63w7lOlRBn22Z/bXqN349eRZKo0qyeTa39+jH1P8CYiUkRfbwsWHw
xrasWkgfbuAbDUvz0W9REkIeeZXPhfcd2tOZNW3ZBcTPkqHn9j4uoNlvI+1rPFSS
uXMT6FELpVZDKFKL0muEGUfWY5L8fT7QaQ4jOriwJi/y/aTHZ30Bog7LIYumhOfX
0JeOU4+Ll5gMcun/gFj8YqD+pxxIs05pqgHTeq23SLvtkX7qaRdbjr66ZX7Ie9FR
KsAXp0VZHQKRvHMlM8C8J6ZV2nJdVIgWw8I84eIJqwmZmV5DkOZ8eDA4XSdffp1c
LIW6D9v1U6ur7RXkSGV3+5X5WClrN6EpG0qMWRAUEf3zIOilwV1ly9cfaI+vaW+r
gNU1IefJB16WzPhwvqBJdsO/PZUkr4ZWn+iGXp/ndG+8qggBWPdwPYcd62or9zzE
1N8hc2d7+zAvbjhw3BQDptfhOufRv6OzlCKJcC6TDlkcme1N8Oxhjv57MAjdsvxX
CQMVUdb+keAwbRUFNRdD/G7jSvT7gw9w1XRTXwBgkHdItFq79nRzeymib5XANf33
VjyKiXSDhhG/hcb1VMligo+zdFds3bzjGWlM3/HcwQKwCm1GmgbMs5w1zAm3DIhF
IgBrFwn9OYIt6qXtDBZ3G6UBFMZ38rC8N8bM//56HlUC3LDnT23hHndDAdDmVfIO
5i7SQelJKYJXNow57K23szaOiYpb++ghuBmbdy3NLrlnPt5CsC1e6BTS+QdQcCvb
G4Iagr3dnjhtTm936qiaFfkGXn5JUm5ZUjpSwDykFjnH78Rrl3K5h2FjRbTYVrv5
NP43r+yhylcWu1rYZCQLv799KUILZg0Ebc8Wm6ZbkIzJYqSMgG0zlQEoH4R4Tll1
HWmjeVTcXLWsR6di/r4OREkso0EObAqcIW49dArWJl7xZLL4AigvPpCAy1zoqdMu
HAdKXByuTtJPc3MxysbhFb2ofGSiK1oCou+hBLnZt+INE7D30o67MltSVdOsEhEx
x9NTDaW7/vuRzBTYBVqOZzysoNXz2Ef6rzIuJsSmVxqCn3SE77HsAxHA4zzM1c+o
z1JMUDUYKjr19vuJtIotTU5nNywVWGCZdESLEWmTAGi7g5G9Mun/sCT7s/401FIL
AKvt9am0fxSznuAVHWwLidCh1unc1D/gpCcf39yFS0JlNP0cq4evav2vP/pqjICP
fxgnqqpuEZnamQq0XublsviodQ4a+HCXkcG1WRocmI4FTWMeC5Wy3O+bKYa/8bEd
TdoW2P3SDiAXSs8KQa5agtVHgo93MXI0JZ4x5Gw3wLgdaG9hik26pyslMarhrEFI
ps4PVxuKpO3ceXpKc1hVJxtP5qh0qH5sM2O69/R7gZd1j6RTmPbH9X9QX/SYMYqX
QEYbJUy6XO14y5g0k16ivl98B+nIf76Dq58twg/NL0Zg3WRqugwkLFRa7EA2Pkhn
L3qcQ+rNTopPKmUpuDOQGP3iqB/5D8OUMHHmqVJQyDb2g7uZKDoDMgLHyEhCOBcp
ZkuI4ak1Aa2xsZxsrtA0zr3mOJvfkl9UDYlzRFb4RpruhrWXxU3oDFu8nBCach7J
YXtRsE+Ex3QrXgl1+qTA9zBA7ykmeN+QBvve2qTZ8MzIPJKucKQ8PEMOl6A2QKyO
a+T4vqpiJZB0bo3zm1n0ugywIXUQH0myX1g/ZSGsPpvGY3xkTy0vq9weIpmU+H4i
qXXzN6gVZFe5qfmPnvu7cS9kb9vOJa7GXsRqgJJLXHrCHJqx4GteyrnbWK2Kuml6
RWkz8+zf/6Fm7zodyb8C8FDt2rofIe/WBStdf0MYFX7zdAUvbhOyyqpMgnuDCKNd
EP2uPBLd620TElFWQyebToxl5wwrqlvKtCTfowqZ+JlCcokC7In4Y7CP1COpsXbX
WR89PDZLQsydf+6rAZY+HTOczVvaK9Kp4lUa/kGOLXZ4teBiYxqW/WVVJIBq5Maj
5aCpfkJdlOCfAEeoysuNIdyMyZIPin8O47S7d+ECQZl5d9uyewu/qWpR5/ZAAh3T
Q7VN28ob5HG9hUj7ajPwzJnwbyUT4bV2Hdyi9gpzQq9o5rdjO1aZC0K7moSn7S9N
9rhdaovzb4y2b+7lxUeaGodxeFCMS44KxhtfHeCqICfwfA9tSy0a18BKdBbwHXnD
qRf2iedCNGyWc9ckx/NNNf2PqUlOiwaS00ZgTDHCtueSh4IOon2BAzR6w6kN9yYQ
W2Dk6FGs7xN7tyv7DhoLWuPQOkdp/2YaM+QUBaGNwUE+KS+BQqzcXZbzSHDovIFy
IxLkcvW8mGYC4Nn9Zx3ibVTrg1SsaDpwHa51FzPpTrqmBARfkUtlqkc2GA8YC8aQ
JGJ+JsRcObJLjyZMT/Dd+DdtGOhSGfIgNWynwY/pYA4NIFPB9Pn3TjUNnXTajEEy
fYedY0dHDstwFsa+O1X6WAD6H3SrW0EXppC1PoXqr8hXHVdx6rtVWRnj30vkuJZY
FsGpLec1Puqs3yRFWcr5Ri4jy6G0hTBBtRSydVpChI0LAaNhZY4fuOIqM5fzQKhe
QmBoE9ECFSUZjt893k6ryzRgy52F2qNVu5jU53Jne/IoQQjMDEW9Yo1/2wpIm6rd
p30t9BECdwex7j8ZimFa7ljHh3XX5zsmlf5yjaSQxLnynRx1mHv4jmGLWnoZU/n4
MlOiMSZF81XogzOivXX9fH8kzAAlmT1mWpDBWm6Q8cWyxeIquplAHzvZNjend/91
LbPIHf1+CHeX3Aqe1GsQePH0/z/PiNjydMBEU8hqF8HICE1clv/w69Q/u5Cjl3Qv
5I+uGy3JMD09l6xDT/HPDY3IOozpIyIRyKmL2qK6TnUFhvq01mhfDmp5EOgBk3lo
PdSg84Qha4bUcUzaMOgfZbxxbEZWKtmjb8yighBbKJZwMdFLfju8rNyl4xB3Q2IS
XLTe2vY4d0TqmGjWUF6GF10LZzqbFgtuQrGGv2J4qogOt1ojfdJFo+kscrM013BU
VdP7On7USBc6Usm2vcXa2177WYOCK5qYvm9/RvPkcBmqIr/YoPpLDsOclEcTZ6yX
qWSvgVqb2D4BQZHE2TcqQYYuHA6nJ5n9voqaoiEAOUGVpCpRnJCrReOyMG4+6Ag0
Cl/xI9qFV+yfElmUsnS+8F/wv6Y0JIgbz9MgP38Y9Z5d7Onq5bMIytzqOd4UIKBC
WRkmaMRnYk7SCeJp0ynr86Gx4jYh9ucJycu2QWNLt6PXuzY2oCVPijEZMh+QcDdY
k0zestSwYZP6CA3jJJWBbFlcSbqkjz3zNX5JfuPITMd1x7/dr1eiEU08n1eZihdU
k+Rr5yFVN8fBEqRo+OrvWvnjXyWKPfjgheAMbseogQMF923VSxBz7AwdAtlafIiB
cLS+hoV5M2I6+v+XUnCr48fy/TLOUda8wt4+H+hll4CI3McaTCiuI5xP7I6xhoMq
OSo1XmeKlz4qOoxBKkaMftNONLS/u2imIgXcKW8zmlcX9RGuAM4aKplxl0cXW6ky
Y5dYMdvaDj3juL5TPvDS5mUPl82u4PnzvudXRFSHRIGWvYJsb1nCejUA/yJCOxXC
mIBzdEU2V2avfQtTNc8ZkXNPc5eef0ZWvJNjVstdjnTnZIQ2eJTZYbhH/+8SubxD
JEoj1icPFgM6UnJHriBZlK9uyAidhQ4FPCXWUkFewKNZyKvpD+JUQjmOtRb32rcD
lBh304EzROVtCxjqkGbqMI3D9Ock5Qw9FRaek6E1FmYQp8peu7SKpHL7om0EEBV9
cetD2KtQ+qQFFOq4kebsb2lF3Dyg0FrYx5WvEH2n3+lXhC1cmhOpmLO57p52HNxz
0G5WQC4m89U5bUi0jh/bTexDJ9T9KWNprlEMbak8SXL/XXBqDeuygmTHRcubLw7t
OcrFzcPc1mLWA3lumXQwevzEvgALNXw16ML+Ywxp4ZCU93nYGyiyICl6ErkFgCi/
+MnZOEXd097DNZr9Zdf5TDpZq62IUvIQw6Ra8c14KBHVU1pYSymJohiqg6j05/PM
RnDijYPiexVyU1TXUvJqySxl6ZoWSX2d2mVgxKwNoNzEHrrOmJ+xlk0VzjMJZb6F
0m5CzW5o0BN7Uw6Lk6/PnfGneEU2GT8IRcQiK+Wjzptafer6uPRooXP+h0z+lMSb
Gs3EXREa9wBnp2e918XOxnF06st/MVWw0Ja9A0aqZlw+Xw8SyXG77eVgy2XOeR/m
3rGviLx3U5hB/hrrOdprVMD5uDuKDjZIuKJexnp8KwwSz9yMHliun9m1xUnmxmQ5
+JwXClsz0uwbmqVPrB6F0ZDBAdiphJkH3jTfNBl5HaJm9iYVcogMbiLoZ1W9yVLs
AZuB829/b/CaAeJYNV/vB5V7ggruqMgdo1uoMr4QLN73MyUrOZqXn54RP1YMZqxY
xyoID5YFPqH8I1QBP57DbocnfpmrstriwiPtE8RQCW/ylZIDM7V8xjA5fDZIeShN
gRGFJ6X7Nf/ayjLsv+CgUUEOItoSJq8XHdRieBUQgN6IMuM7D7eEEmCTj7UhUgw+
Ap/m+W+VzzZJ5IB8UwVNZ66QwJPWASaASv1UwpJfscLaXBel54wUxwqc5FEApf7/
RbqxoVyAUcgi7iLmVxzzq5sViPRYXlZ7wB/HKdxcnRC6+Zpax67jWrxpuSn7Lb03
2uyChoSFdSAhn8P+xMzYWoDitRfLLSgiI3GTniHRUW8zzPUjiW2zMlwM+6DsOyny
Xo5t7nYtfSGRI2ngQakFmuZ7i/D/CLLRP8k7WY7s7JzfEIJwSZHFICeYqSFjaUSI
zBPf3/+9h24KJMsPBOsA6xfMn4erN9+yiXIZUYWpk/h5vOtq+KRx575vaPLtniJT
kOyuYCg+BxAna95Xr5MJTIlwMujW+6dahJKZSdCfHEjuz2aMAkBJqtbwsHApKvGP
1yRhAyMSqackxy9GFZikJT5cO5mRLLOdcshbv9lrhu2J7zRhJlkJE8Blqf5LKFu6
eMeSNDnYM4rYj1tMgr09nwH/LMaO3gswPsgXwvAvKcP/NMFDDDh78QeSTjepHxC5
xcGuHK5/pDjHBuux7wZU04XDTTLQhwmKLTeOA+suTKD/kOT12E2I1NBBWUF85Ft2
vlQgArGy9LWJqWKeHy7lA7P9UV54jLpkJV0iMX4/cvl2o8pBRV1gQUMMs4isWST/
PJQOlEgfDtoPzFd7MoVpU3I22qnN8j7GTgJY/tj1EN6n7S/Z1Ly9O6mq9JmBVn0m
pN85AFdtxl0dBUqjDAabDbCrck0FI+ndJp+zwihs6kDhQP+a2QS42FIWOdUWWHxN
1wT+0Tw+VioQFkPlakQPsYUHbxUROybw8ElkpJ9pOBilQZxMwGFpcy6N/7bUqYvP
iIyUlDBt2oWKuK2grkZ2W9qRW83ozeLGPwFnR3+kFSjtwZyYy9DeOkxog7P6l3gA
riE26z3ZYAYYIyPPApa+A7tcXtlk1sUAPEAcC/SbDRoYBK/7orA7go7c28/lkiTB
TPmpAW8c1Li7gjui+8e+Dkiq+FE9HXiOoPl+Bc6edeoh6pdXpyE53G5N2uxiMCxA
DdaFUQyG/TDfV/fXgPquMvisoRAvMhah50P7Ayt4o8O67MYZKqqGv4Cyd8nl2CmT
cAzzfiog/QJ42Mw7c6F/fikRNw8xZdCgllhp7C8iqMV5DcCmTKrlq7/1K8HFJs9d
Hjf1G1x5flBXm3LWQBJ8Gx81vYLIJkBYaVDFdeH72Ieu4GVoMN9r5sJqwTCd+Qkz
c2ULNyWWQwh/a2SPsARwydtWPceqiZ1IVylxB0pUxFs2Hu6BUf5U6evFbuh76xpL
WVrLeUAeAj4E9x5U8a7Kh7GRyhBWEe65YOE/l+GEvu8g3Mm6MU5DEjKng917Y317
zcPHBdsvjkYxPKRKLTFU0Q3jiJfbHDHkeCMgwGCt538OuMoD/wvh7HtkL1VukLh4
00nJBm8BsqL6w4W1oiextI61tyrqV1PSqUdvG/qDGRt0uRh4KdQZqUh2LXnbHUXA
IQWk+82XBW6xWTh50edy2gljRS1O0fm7uMYCQ+YPN9F0rw1R2KwplmHJpKI8XNXa
9FLLkIhTM3bJ1l9Fc/P/j6GnofioPpaHFF51oT/dk3zxNgqgPabeyxr4HPig+YJk
515YPs6ITbMF0YS43Ty4CMPeYOvUK/pq1/PYSBuFaTjN3Bh9o7UHfK+wak+ZMDH5
RTSizyBjxuBsdF4peYGtYJS4B18kfsnkR5BCaVAfRdVTg/RG4zXqpWk5JVMY75HQ
HSQSGCyGkoiJ3BnntpylrxoQPDxaAusksBlG5hJdk6a/pk0zJUbZ9hH2DBgmuNj6
q/OYPxI6Id3b53h/R2TPHDPYmE15S/2m4A9GwCtrrw0k2plgp3Q4tsNzEiHGR0us
f3Dr9TLJ/oERpFhUqqoV+EaiDoYBx2XxhIfLY8OwZCzw3cXHdsKyM9m76fImJAhm
QtkFrro66srgiMDjVC5oPLxdiQGGWk7UAojET8/wvr+aEEpoWMXKO43SyOlb+m3T
Ojh/8tE4Gg1VJ9dBrSPl+euOAPzEuTAn+OCAdiXWFEbdWc9l1RKSdeMp0HkqCzhG
5KAiroYey+CRQqaQiOto1eMNA8j3QziICbEathC392zSK5zHORqy8jbdrmeBlNYM
naCpGiBq7LZfsGKx/fmEpvyAo6+OSYtEls3COilFgSiaJvwOX7E7ivV3Bz07G018
GFj7OhfM5mAEu1UcwoWAw+bwVn+amJ8j2o270D4lsc5reETEdw/852OarIOlkccs
Fgvqqy8IV4w4K4PNggLG5b+EuFCuDv+bCgxAcQcsuhGBTNhtoKgBIp01tdOih0Q2
EVDS03Lp8ONBuR3Y/W3Z3qjALih40VAK+VZMOBVYeOWyc66n3u/q4WQeavSeIfI0
q95GY1v/ltctkMdBoKEmO0YpWO3x5OSUikHo+LrxYjViVsS7GPPCpuSxW4eY6Io/
+K6HWixYEt057NDSapzLDMXus3XIXn8XOlyURxrxviNL/MSIuJ12DK8KdirkxIqh
cR2hP+m3gTdM+k7XlQ1tYOXPUl6t102TLe/+FUeE0Sxhfoaqsc9nwi5niVcJ7gvh
aQDgk6mn8XL7zyfrFX5Siys2l0tuuT8L+Yh3h1kg0nMIxHCCsIO4nmHpQ/YPRcky
iWg1uZ2pteSTIMcusBj5DXI1frw4Qnm7g/hIFfpvSE8YvWLTqUU/wNg7TvLOOswu
vYYORpi/85g8ON/p/pYvwZOdmRIuJwD100IpJuUPWECA7yWdTvsDKTYKWSPOlESM
CkaOUR+4qbGcUSaIem2V/wEcUotZzwqXRMaTHwHpO1oZbMqTqmufUcR+xV4sy8Jg
wolzvVq+Hn1AjnYabVGrcgMIyyzCqor8gYyuk2ZjXRQWArFFfaPuNscSVAwIZMLW
CXkdlME2DzSysbqt/iMJ2PsxZcLiEq08Fhsz82MiGpyF46golw7hPE1J619tfnPL
rx+jDYJS4HrIEBH9+ppcy8a8Bm/JBXEmgjmW87QXDoQb+7NXtwB4a3nAq9JBqAk8
sQWePWlr1BhQLcujAjuYtEizpF4Ixp6Dtf4pn17OZJUzzR5XzhSJCkbSqXWJJwGN
FMeC3hCBfJczvMmujNELFK2rZLzVs6hsj921R2Hv8gbvm009WGILrlQqvFrU6cs6
c/BXBkQhHuwVlCPT7jcp7A7DWzOwu7qxHS99h86V30wM2P22o/JQlRbSfZDx+SJb
g/uaQ7AlIYqTGUKTGplMmKGawuilXAlE/9SbCEczCcr56HynX+uAsk9iDsU+TL1L
7DlYrz4aGakOCZ0f1HES0lj2VMnjM9CPGGRLAqKOY78I979+Xij9MJZQ96B+plH+
HzIsCK8O7VC9uqItipvQWJT2uyC5yBfzC1i1XjX3jh+iED2hW6elY7ecOLqdqv8t
Yec0fxX+GLCRdgvJ7mDgjA9kjLG50YGbenneMPrhG+49OepD3NHgSz86RGpf0Gf1
+xMCYvR5LX3VNti/pPVH1RNz8OJIE65zjvyNOQUmTz69hCXi2l85+ZuivZf69I02
vF7G9nBJ+cJAdiFzK0pTlXLf5LNqwmw/TS7CL4VaCqBaUaXnVebjE9j8Cc/inftL
M/rOAot67YicZHAN67bDvTuyY/J1/awMsRcqZQ5K9mYb8XExK4pM+gHu61dYSct4
f+C3A9PLtAszcNRejPAcMNfhdTtNkqKPkTxxGt/5CFE8hFqacIYklVVHQdKP2mDT
PzO7aOsLwJzdj0iLVofJG9pe+15vSgwZGtShzFvt5i1vhlo6gRmcK/e78ha9L01O
ChfXOfXu2ZCijmGYZiTNWyZsYcYIwe3CjM3vpvhDxglzqbd36gUP3Tl7591lTGrv
UIUVJvl7W7sbl0py+0AjikwGK8qogNyaL6DWro1B39oe2X856++DTOdZJVNJzRyr
gnw1MzHOS+KpT5ZULLAXhIW9ZRTaw2NuTzdn7F/7eXzfK9E/pneo2sucJ39/R+DK
12K2kt4Nxtx+JImgc5H2QQVN7Y86P+vBPUeqC+bdikBr43+J98Jk4kvZhEQZ0N5V
gMwtfjW9l7YeN6zA/msJ56rQUer5K2I6IVd3lTF5uUvUbjr3USsgl7b34EJWUWE5
BszpHLW5Z2di0VjzRvlnaHoLXnpsUUs1188iUrBLO0tm1p/e4crqpvMIeCCuq77e
SzJ78lCUZ26vJ11Fa15ie0dRzOwreNFPG5H84IlOBEQ+6AZNW1DQ5gcHz2Gg30W9
4/pXRVM4KxUA6TBsydOUm6+7w+Yvh6I17Gm8wm6LCcfOCfwSGjM74JdLw6JWCbT3
6aSwnMGph2fzwhcIp+ebL12q2xVfY6lb/e2sID2vkqgrd6e1uz0sdwKmmPGYdUIv
O9BEd+17yqktAU6JqRCbXJoIuUca4a/RQggmSlA9p2ncJkzjy1zsOioFw2fbAPWY
EMHxr7cR8O8uatw52Qh9fubykN5NnUyj+x+BcDg7ziiLDBQGlRJWZohdlP3hZazU
fQrz4ZJjgoWkilZlBP3XqSEwh/IqTWGrST2d9yOW/nSq/RY69rC0CW9Xs14YyOMX
Kyq8/08Enr0QVXVpr4wHXDQuiU1Ef/oUjRdC7U87sb2RuGnyfbXJRnOQ8lfPbHYe
fyJQUJVJUkMjiVe3F9CZ5BpCYPyC9FxDbF7rLmUvkrA3P201X/wcoo4D+ouFj6RT
XcxzXVGVDinjvUfRJuKdARNK8Vnbvuuu5fMubxSWeGlFqQWFusTL05ZA32UyzHfN
rjKPnm9pe5uyfVeRO12pd7VuQYAWlb6XiBaPR8pc5L7qYOkII/XVoX5mU7eJDzLF
WpcbL5UQs6QVnz67fuT9EBvsSAqzOCsn9q7j6eti1n67PVpk9n8ZokrpKUfTCYRV
Nt35hSDtAnoEtnuQAn1CWaawOymyVOVx3lKRj1bKjV4yCULNQdaxVIQL1+OzMMTk
s9qGkY4Q0BPqy5HC31MeqLjI8W5j56cduDVsiwRMDB1MrD+l3cqDVncf9q1t6MIK
g4X+Iz4pXG3MckFx1YMTFAJ1CeNllyli95GeAm9Nqk894ZsPulS0YfmCzY8/zx3N
1wRRAve/ezdEPfgAus/OM5dxBUXSIS71+rWPbMMzrkFYz6SYns3h7wKmL4hv8s6e
cfyM2Vxr55GHcu+9qDbtTInWecKS8gkHmxk/fKBSCQITdjkqXoxD52/zjbaZpV92
O5+DOvPxYVekivfBdHThG9LM/5Bu7y8uJmHX0bxxl3/SNAKMvzvkLioLzkaoYU9H
rZD9uX8jhHLtgpXewQTrExJhCvHsdclE267k5XuMzn8BSmWBNFeiMZtkBWg4HLzA
iyDorU7B7yvPUnXetPRyBD50yT092oJojp36B9fOtKH3TN08HO1oiXY4sbqhBurw
HtttHeomucckQtEbmAJgGmEmHi/NCK1yZuJZ/YOTSGnPGCk0WcQkDR/f5bu/JNwq
hpAj5lFMsEeLhm0JC2ENGu51F8cg5qewNZwt9w/D2KN+F74Lnl7v8tMBOfLiE5+z
ztTrRMPKRBfExgglli0O9XT3gE634v5V1/Ff1fpQlvbnRzmD22O3E14xsXCf0IUK
llmAmeRmINbXkqRmis/owAVjned1+pBzjgqhWkSWBy5rhlmc0OgC7BJMR7tnUcJm
Ekzpus0WWPlB5Uuc1YscHlD8TH3aBL8ebJQvb16xJQkPXLEZWD3PfP9B7wBW+FLq
wwXji7L4uIhaoTQFt7D7tzOQ7QcA+M7J6c/PguhydLX1usOM4boLkKGdcE6zMNNT
kwzeONG2axCGSOLOdLJSr86XzIXArdhB4dA9WplqBvEjZpfvmt1E0Oev1/zXEng1
ZOdUW3r/RJY1ilposdhCmF5Lnqp8cUF5cNk3+iGnOztrZVMfK+9OlY1KOC+kcSfX
tdixXlY1iU7WwTt91xF3sVlNyqAjmemVFROdKgYyB8NaSpIURaVhwi9uCAC9r+Xr
i5VoBVZn4a+5RmXk+BEomdolVImFb3cxKfBksKLTUcEuiF0mjZ+wq8g2V2MDXcod
rJBXTy3vw1ahO4R/HnJ7oGwoMsPAmcHOC5xVaf5ITrm+9/hAY+8AOvaxoyKlBUg8
K3bG1A0daI4u+gNduEO9eEgV2T7Mwwe2vwzLDBtRRfTDk8Nt1LV0YjHl3ZGP9xOw
cxuP5NIXsgk51G6Mu3n5kY00uQ6N8e1YTCqxxv61iKUM0ZuM/KFZCu8doasEARo9
z8n7P6lWBijlga7LDvx/Jh7kf71TViZqy8RAbFPpR6/k3C0iuYtQ6B/GzleUdLEA
oCyDm2DdiHbVaMbDrSG6ISIMEFQygORXa1lZDqzUwUK9AclG8upZZLF35QMozoeP
5jEERWv8ue+LAfwgY6EWUUIJwG6st7D1jWCFPIGtFuQ+3qcUPpKMwr0T/zzAjMqK
gaYkcN6z9xr4xVIYmKyD2IlG7qgIPLQUV2D+Pz5BjHKumRNx7gOLHzArzZ76LAyO
d7FvPZL76jVjZu7QnB/O49QF3kAIzDek4n7fzmUl1u3BbU9WVrjPoQDNvCaJ7oHk
2zVvAls7PMVQdq2Mjr9eqvtLyMfKh/jZ+ca1BxkfzsR/WFb00hJeEJmPixLoOWOo
/cwj6OzTFjI/q6+CB5OqLL6BcYSdw0vP5pOQSkNf/4fJ4x1iUE7/sOddWLCMV3w4
XREdFPPxfdMIuPJz6Pkv9VPPu9V+FR4DF8PZXBDmDOaopfevUjwCCsj/bavZfBRB
XlInmUevW3DC1bWzAmkMATXyTmHbjr3LgOvym4aKf/M3omvVcfQDJTQcNHyoVsCb
M4ghAXSsKz3gaZ7XBQaAqGnAz1glJOscWc4VcGcOh1dtrmsKJ0gZWES9GjLZUBVl
W4ua2vJngcwTLZ2SgJ7EWtujy83ypZivIUHgO5k2zEqy2sXAKBmwpy5ra5GeuxDZ
vuvWp+B409I+/5VbRhnh5c+1HPA/RHhu+O0qc3gMuJyH3F1rhiPpRccHstuBvn1R
XC1xHBCjGrQBmi5/KOvvEjXkWKASBPfZxjjJs7VbWqmuwdJI6uIguhmQiylQL49P
Bvdzw/x5qfaY9GjW+4xlDBg79RmbleSVxggzcm5YzL7s/usgpKtZrJzzMNbR2x/+
nS8yPZSoPEBhAuq4IeHEt31yU/96rvAHTPIOH2C+6KaMdpsgPrVGV+lfBw8mriAx
+CPWuKGW8FYUfvOuqSJp9rqa4rkZZaVjVDrZywJ9UsOyktQmonCtP/PKldE3slPr
jsDoeP+J+l7Iup6YFrql67UqpwLsST3uJ5wNBDYXMS4k+nIFRxxCmaNVmz2NQLls
F80dFE3O1XFFZlbbAhSp74evOc8G+llHuXanu7YE1zKZ+IOfh9TSkEnQnETDeyO0
o17/CPdLkHF9H9T0zkreEAEONpUqmjuX4MDJ3dXZmsBAf/jnEYn7ZwMLxs2oKky/
ykHCib5XAojnO4gOGxrJvMgn5HyPCK9s+qBomVsNsM09IwBCQeqbK/gk+u6Zp6IA
xRcHGUuclYXm0nDo7hKp8yKbo6xW0eDT07vsuOSYG1sLAf/cgqRPuUiAVL592vNj
hv/lbIv2KnbodVnvvHdrg5ynDGHdERaBbIYjn0DStvZAbcTp4ufvXc94gFmJ9V0K
AMkK53xKVjQt9Ij0w5tdw9x7+hmGQhdFSR3G8IO6hPJOHZiQmaDB5CCt8wfcbzg+
+pwnbn6yFPnQ+DjN2y3CWGWwNkVUx0con6P8XKZNaK1p9Hfag+Gtn4VKC6+sk5ix
qygcND0VKri0N5KOUPWoCx2BkVfLp5kbydiOiUCPTM7qDqQWflg14txlkIYjLcK2
ekGpAkEc6I/phLtgplrlZ18YYFFirah6MP7AUVF29bF95+niWlO0nADGIWB9ONi9
Dnkyi0S8AHU3XDnSwkTv3pl55/E50d/1g1pL/Tcqd+Nx7ZjN/7J/wG0WnpqYbjbP
xp42Up+x++1wr0KwsyoITYIloKurqaRtXvnoWgSL7hjGOqXvO2m/BdqhilJLzHMN
exbhcfAocPnXdTVVwHTAUPEzBSsfaQJfqxJbq/o5M/bjnTG/dLkHw0tzlf+G3Fup
6eXmSeyr99TqMDVxdf3cMVqLQxgHBQabj1qX4yVPA0ALS4wx1bTPufuUBGSSvyHZ
upXOy3BFBuepO5kcotPTJlw1qHIYSPdznXyKc5vxWWiVZtiHgjl7JVWkOYIRcdLn
DdU7HQf9TPrO/4PvuX6n4uwgunctiZWU0VYcj8odRHP6wP2hzzu0XZnBmcOzD+sA
0KRuWmszfsOWrmrytgWIyxMIln2+EtW6YBPNcDN09icgmltMLbyODAYD8lmvktxE
qQdqCLYkV1eZcSu8aVxXysTR97nTAOxEwCzhgTQnbjZG94hlJnKINnXE3E4mJ6gv
CbDbFcAyZl4gqAdvl6On7F2TsXtPQ+qo9mz0kkM267oKfv3lBsYATNACxYCimn9m
XY4A7r5a4IcxIUeiWpKggewvTKMTPQWQMPzmHohPTrU7mlpfBtJdMrXycbh2gdYi
g35wfGRe+d5taqcHQVaMu17FeP78n4+7Qqb/t4DlBOOk8cwcgoA/yogjmOw/6Lra
W3Z6QiN/uYihHKLx0bHCqdvoOMMgTRTPOcxUg/Syi0pXewEojAHmok456wtBWVJC
txwKXCAHBoFSgrN08hTYAC50h4PbKrAnJymfNrY6qkQH0t8mk7CxY8cW2h6DGcpH
lwTphubzOcBtCB6bq3BmbUBNtjTrLilq8kSv5cMhmsmAbMhlUxxhraNCguW0j2M3
eI4s6jrPiFh+8h9VZQ2WQ3Q6u3DqCxuP8swUHija+cnlyFlYJ0PLJ0FaYajKZh/o
MJQgpiEdEuaaaleM6X3VzdqHtEywYQslCvsWs+keeoqTRWrbg+4WgFNrFhBB83ST
QsCqg0NBuoFxxq0Tt/DrhJUu/gjVckD3pAA+zU6HtXN2u96IJcbv9tC5PJCjW/4/
MbwgiXw6X9CtvSUNJGYSkZj9CQCBy/ZAIVR4xxAkOah5/kRwfnvJzmA4ZkjeCPsv
iUB9a+18ztJ9jLcfYbJzIJka0udpCdJst0z9JfpV8q/Cso1S2Ip3ndfjAN8DkaDU
TXxNueK+xMu9LShKoh500om6rFOuRyflxuMDqX1jrjiybD9NcNyc4l/afSE3/aIU
dtc+OSI29Wj8VfZtOYk5y/XQ3iXXdTJmKhxC4GBeU2Tg9ZTp4fEv6vwa2W2+K3EN
0LgTEkEwQaDEzzzF19NznJVsnkD5nz0DPn1ISmv97LkulY+UsPIdomR0h5K7AT/z
DKP4+bDjQ+0gdtaL9x0xsN+8lMpLW8+P2wxm4hrz4BPlMLebGi728yF3MOYMlbx1
fDgOk2FUUUOhhlBv6HQXVtjVELGyzMSj27+FzEMMTXdYbs4ydXNhCXxjwVhGFdFZ
SJ/31UJeuK3r3PaQPNeM6kem2r2MtsF0/ZKyBhWeUDAY9tBGBJjKBwUgIGZ1bPVK
VL7tgDfvlicWVkCnRISaiLD9z12iXj9i/qGdAMOuc+o3VTRgTE7CYP6898Ry2d0e
KlTcD5eDYDF1fUGlSDZ24vAv2VWlmys2R4ZM1GDPY0zZso8ufQAw0Z1iVbSUqPGd
RlgFOoiyCJ3bxy6XDuwQ3TGrHKApLSEZyW6kDkfdcl3i9V7opAba5Fw7uZB8l/K4
wShDueSyb9K1rKjPrszAgWRkAMqGWHIw+0zVdfbIxXNlB77SZNUoxcOabq4ICMZf
Vymmvz+2Nw4SG9xTn5Oc8sHsd8ondOpB7mtvWJtt+JlWTDvYKLbqul4mm1/hhUNF
Vd6/DwKZEzMKTRtb0Zt3BPoa/GUky1LTwpOqvrAs8zAZLVokVaBvCQvyKbDM+gGb
N0uyqvHkrYgkYq9nasaIcbiOFvPuWDGXWtGXOwV/XZhMnMTa2n8xxUqEM/M+k0Vc
UgLfmvv3RgOuL8QeyTBarzbVf7RjPtdGCh8M/rM2mqQwXlEaa8rS5k7P0LPsr2kc
UjlknL5pG78gcdBDryuue0tbxPu8L9apf8+XjyQP4/ytWaaH9WsjDAYOZ8jke78D
3Gq71oCuITon9gQN9NlNCU0GMJZiM2XYh5lMWVjzMkT3En5Cb4wps5zJY6wf1PNF
ypDsZRnxb6wW7zY6F+92Rzr6QcKsxJGurr9lPeYrhTbNrCzwbyRHKjRojVybLCiH
p0k4qrof7jVMbGUd6iObTEow1YVP7zAIB9b72b7U8uitHcV8/jo1mC58xLs+pMRN
HtCekfPIgsfj/zKPg683gvW75otLK9Blc/FJq0kIlFHQHIT70AKi3RdjoGmbTr93
5fPJ36McWYPPDYcZF9Yb8Eo7rfGxfZwQt9M8oZbBYg1yJLuVTi9UQA3iEHhTJjmX
JuspYB6CPhqJ7lyQ1AlukMZ9LC4iW/zoAvfNSS0fKoBLmhWJjo+L/2fWM/5IdXx5
iqb/zY7Ht9k19LLXERRPkG73Ivom0373cSWAfKbVxq0G5kjBASSosk4OF3MKpTAx
2ImH165oH4ssSfx2v7VSmXoqLNGWoPdWqmb98bYaAItzx7gn/li+3Obj8UID+1Dc
vQH4JmpvfZkQPKQqvUymcQqNMo0Uq+CMAkLW7vQKj/5zJDEiR6MDME2JH6Vg+AJW
F9sxdK0raYlQo9uEd0ZOU0DyD82W5Ar+bRIHG4A5mOBKRmtaEoundTtte+tclIez
gYaGGpgWPzrPJpEhKD3sOumMC/+mNq4WvOpA03jxUEKIbU1S1iR4gqW/dfTQBBzh
++yvU9YTMc2P7+bW0zjKT7vOz3pN2IJYB/YkUVsqIAjdfQtqrUXrBDUYPurc0APX
4SWi72Uo1oSAPObrkwhHM0KVwijNhFzRgBLpNQpzD+7J8mcrzNUzDkyRWCRbRsgy
CERzaaEHbi8IgbJZT73DNYX/jPUk+356aqaweLck0z+NFEbtk4KJxDXXUNU/Lkoz
6N4o0KuUVE2Zt0h9q8FT8+1MNNVS/GAyWe/ne3xRNXhNv6mY1d2SmTHM6g097z95
V6jqGLSi2evurBWRNHFOHlCb4brWpmAvF3frdAl/wOlj/81GuQEzsxERnapHBT9s
/RdZu+uc2swUwv7hUolyKkm40XOU/Z4Em/+lySloO0eoWiUWuFMXc9CP2dBspHPk
ZvQOlWOBY9k7JLS3z84Jy8tOmp5e2zgzwFBFje/40xrrLbKHuzIHa0KGtloOr0lP
Lsmq4na2/1fdmlqCNsU2XRbC7hDgNe7UhmwYgXwuVAlvAPSkxRVfTuLlwdyf37p/
oZ6BkHw3XbMn0HFs0Z9UAJHfJCbaDfeFHBmC/N3tyMioDMnl5nsFOMTMnPBvZMav
M+OXNutT333pbh96mS9JAY48Hf/FdcUcyEx4UruM5cQmxz+vwxPZxJCsoSOWKPhH
S4X1FvWJ9wSn3oA5KaCdU4QaK6bwZ5T5e6XUuzGDWqegEamaqi9q7D64AopgkqBI
vTzfRM4m7q2VO3kW7wqSuJIapMj2cmk2Xn6Ksy/SB6U4K3cxvSSFRi9Ndjg55N1J
dln8sx+ICU7+zU1l0JVBxnPxkOWgiBnrieDCTArJHgA2+My+yHOih7l5hPZK8nH4
0iasbI2FtGuxOQwrUqzfcBSTHYO+iMfffVXErc8eyWG7BwUEeSDh/cDs0w2T9he/
EvTdNR2OT1D7jOwmRYisAq1Io4r8BEKLHckcQAkwLpcV5psGeBP56EyYPA+xhXmL
JAlyqO/8V7Dy3TuGluWZV8vIxuQQACQ1pn+leLVPmSIpg+9j6ieeopLanX9K5vWw
mFTuaYgzuQoUKFDOaUtqyiJZbBsdmBNFJVhVw+qK2TkyQg9bOX9IO5evSmQH5agL
YxktXGobdpD3OIbPnjUdcjOpxIDqOAaF/ROdgwtWWwYsU4URBIUBIIUFGgqAQ9Sg
Wep1+tG8mRpTFpgQR0sdgSgJhErtogOowb1peUKz1RuCLLfgY+R3Z0CTggSY+ToQ
Kl12fTi+mmh/cao4hdepATEiKJmNSXSuqAXCH+ydmatiB8tiU8nUo4p6AJJaboTw
+6kSqFSZweYeskXALYbC7VKKZyMorbWaotW1SBif9C9C41TtvYDKvqTxfITI4OSq
iUIy61N3rUkRJeUg85xqQNIj+zouh+6LAQx/hXAXDx9eJFHxDcpKcN8jFfub5x9w
vVs2yZsIelDVKLGkih74Gk7Z5R3DEgiA3sac8nQ58IsZkD+9hd9IMdr7ToXekW3Q
DFL/LNDYPo+WIc2CkWC/K2ydllP5exHVMBfoYFBSr/tg3V6xro5UVbLm+lBD+Eaj
9UiNzSalajT4T27L6sUcBnkyW9ks34EM7Iw5iqv8NC3nztBZP0n7zB0QZj7iyOsz
TlCOXn7s7VuWEe1V4k501nfJQF6VQywX45oe2tUKqFIE4Fgkbbce5YOGtIkn8v9r
rKV7i2vCALJH6/9wRO4i9EqU88V1h1xs1KPz7RgGIpzhZ4T/s4ifhH+haT1/2ERt
6tl36X3+azmnPrRgL0e+4jJYo/vD0ECsgw5lvqhYPAbDMsQVMh5+fYyd8zzjwkmk
eiPle7TyUsVGQMCKFVUk+0+KvR77Au6OFaW7N83dOc8FXLNi78+TxcYfg88ZTtzC
ZM6QfLxA9l/xDqzX/Ma2WeVkIWPqwuTZnhXvlKDnfu26wMJZGVnMZeRnEz+F2tJh
jkGbkrhytK4GusdLb/HB3Yimle8HfDchWJr0FE45xMMxraF38O962WYG0gPdd80C
EJBdqN5+9ueZcULQMZLuixkZ6PcKuoJL7ttItNMl25UVxRSiawoC2pJDCaCTJi9+
oNYMHd0tWdePPK3VXemlo4ZoxtkjXjVIhKSyrClcyFrTiktzPCV10/hB8Jf0iViJ
rs3mJSvCaserFHZXXbZndwNLRCIn1Wh3ty5tSlPnxdSRxjmQTh7UALPZ6S68/Ugu
+bXgneEWtTlQso4OJJCfCCVXwDPv9NwCf0zjhwo9TtvOxApFRLvA7xrijjyOsyCk
BgZ2reQF+GD0DcGDV2aYvanHoYKFOuS+o++lYPgX98MNAQdKWpdw73eYS1FFNDoh
KGuf83kmpFV49DDSDz30OZQ5AUqc6z3QwNuxxbiCdvoIs1D2PKlPSCq5L0IextPj
HVk6u3gBNSY8J1JtCIlORavsyUPq4GYRAukgyl3SPidRydaoal0FjjqTc7OI1RWw
YIKeFPCfpQvQHeY1K7SQJun2ZdxycIMn7rdVCXK9RMmMbmT4ayYgYHarW3FbA7RA
tgf6pH87ggACSaSt9t8DEysm1tq8c3nfZpHPktDMQlZjcwywcK8DcECQaUXdHM1R
/D6fjbFEANKcSvRaL3PQe1gAr2IM1bkp89mdxB57KDEaHuHdg/bPx2rY6toRd4pC
3rzE9+pL7N2PUSZWC4taSwSmdRqGrQq7SHa0Qh955Y3qW/PFqt8+0Sh1pvmOc9YS
Ux3ws9eIxfbnTiZKJh0oRGurTLF5HKRppNfHvs0opRFPwFKd18GnYX5kOgZ0H2bx
ZA9fwF4FzjNXxGV5nAg1bMVttNkQ+MgGNmLtKmLE0SUkn9SPoRaOlfwt6qly3PCG
d1FiyTD5m2b4I/sxbZ8ybynwPTpWK/lxzfvVnnErV6itTMYkkwNMuxyASccD/OO4
3HM+3SMsyNlKdX4yrtm1XEdjmo53NeLhIIwGgCB6xWiQrwXx3mW6ehIRALE0cEyX
2i52hBLm0I38oJlZFR3aW2pFX+eO9qHWHVT563+VnvHPujrk6r7pM957KT3xIXIo
pHh3LPYS6pxthSOJWUVbPev//8FbjRlGHep79/8tPjiwmdca9KmTz64+c/UQsqwB
5S/US8ptP1kSF52UxvaGZUhvm9T99Wxk/rOT8VTlAMoW3xs4XTiTwaaXoUbTcz+v
FU/lHRtdmjQv3/gkSTMOZZsUpXVeftwzwnzb5v/x9Y9TFnE3C5riiyl1PydrFSpm
cQT7sUVf7z0m1ZvVQjI5qkGoH9Re2kFEz9+8kS0QWA1Wxvkegkjyl4jURP4bIytn
oqBnDuODm3bQrEVPSjWLpCC4sOT+eU17/ZYzalPYQI+BaoWbjz1zkzf8HR1FMuq5
KEXj4PMfJORMqCKND63vrjxub1UzUawDl2FR+jcNrLATFKc9IaIH4umivEtxQF4/
az/Gd/fZiTH9X5Kpuox5mT07dlZjwcA9SwAhY72EZx+0cB18kllRRtHE7jBD9yM0
4mRFkzMUdKw148LYkHyBp7eslIxfPGlV9R36M5hqdRihJ4HDvGWqvXHJhjcwr2il
oTTBkkSczJGpdEO1tmcXBsvJNg74TLQc6fvGYHPzKsxdpU0t8Z2Ma/KL9WxVPGok
lwSR/Gf352Y6P1C+IN5teKs7PQC9t3kRk238XniDBOJgQBkH80KU56HiSgWtaLt4
I/lSYe795yCB6/DX1lF9V6STpE3JI3MDbd7Dl6w86px6uRwFSuRg2J7TEdAbvHnj
1Mqst3f/uGJGplxzgPl0UqAJ3r74yt0amT3VVw6iwF03E1XmRlkdWU+HjXQ3lg3x
9G5/7Mpg1FNtvZGHhXHuo2BmAv9/BRGmRBL89kGkyN4pVtHRCf/RBJ0wIeT5kguQ
pNoMuirPiVFJmCtkvIx+nO65oNKv8e8EsVlcQW8zcFUXwfKCPcp1FViuwmXkMfNn
v7BpaVQ/BKJAfOETvVRF9IcIZq7kSOaH6G/GeFss+gpwkINklwp+n5vGNW0Rcn3U
/Q2jVSCLa6sibwMAgXx7zPbE/JWkgfIHta3/aera5ZWZuPlqUBjhoTKH2mvZ6A56
PVcyONlxa3bHklV4WNd1lRd8N0KjYxgU62MqBelwmelJvfsN4jhYQqpj5o5SHvkO
tkgVnjQWNlAmc4bC9pfhTBZWGZoQvzvISvzoPKWDncTv4HB12nKKZTL9DghdVM9n
XCyOqci2nAZtKkeP4gFmORKqqse2opNq63ycE443mOeq2JA+UU+obVAAvgqHtEg/
5dBcS/zsE9237OClipy3wssL4S00Sc9StpG4AfBuNjV7/Mbou4eNJewsWYcNy2TS
tY/PlGWkr396d+i+WSlBVl6PtHVHMERXQ8yUqdnFzJihFgH4R+7tUz8B6cZaLXUw
8fwoX0pimtQtKDZUfJrzWXFMCrTXThlKTWuw6aYDq4dX1pdZ37SsxNxk8u1honcQ
vGpHycdffQq+JJsR7ylxHqTzEGyd8bP1T/Q2XHQJKT66yy9y3gGxoCnXLgGDqHYH
zQkQOnrHaJw39qNiDoNIp0qYofcEvRdhMafz53CEEjVwrll8AeftJTi9OcDIZx1z
356bWo+mdP1LEPhjrkrG6BU25Aq/QmJ48GZ1d8h6CH85hOK2FWnbVPIgiQEvFAI9
idOiMS1jmZUdiEez2zzd9RGfjKpTRBkhMVk6NuCayzK9RT3BnFixK28UHC8EIlvl
ZBeXIslKmDn6lKT7RzCujfxcibaCabGtpiBFn2rCSpKRCOZork81+Ucdoqbxtkz+
zaYXwWc9cc2QMJeelaei8P0gV/C2bTbl1XCNZUuTJRAPIPa5/cKH/3xW5ba+Wc/y
UHqRZmeTX97cQwGsjPw/QYsp+Pn7w6PwE2xcAJXRQGIcodk/4+OqR8OJadN1F4rk
/mglW9ryeGS9dFAMqqQKZj1KXMQCH2WMMdIkh6htjHXpROnlPtN9ot9O+AZkM5Cj
udc5fHI2RJfTT7k/Vpy7cwu09KDE9shDIWEPc5z2bURQkyh2uLCz8Qv6Kjb7nuDY
k4na91qQkDCmJfrkRv5dTjs7LUeqXlDKReNYwwqO5dWY36nnmKUTrtg7OTb5ayjk
irVPpxanfh2+kmqzc1DND3REqDj1A+pxgJmtDufuESEecgbrXX1Es5O7xQUu5U6u
09frdfZC1wwvqYOfbQ8UsMZvUfs4oMd5sKECuLEdCrbcQzEhph+EFvvJOQZ8cQZt
CU4e6AIUgx6suO7HKEskAM6zoNMEVFiHAP/KmG1BDXJT7WDevLVr810ZAZk4r3lZ
SrZgxZ/y/0bi91My/KG8/TBsGcr6X4+Mtde1jQhVfvpTiP1sNtgvlsxrcXD5qLTL
CKBaHt7VGddfulyh8h3O1+Fd0CLXBxRPcXjJ/0M6xgrEqcftD7KdvjcNn6UZZIuM
U5MJuDJ+1NW+CwuDZtPPmPMtoYKAoxnzXvvyKTxIn84hQfaaqN4Tw/5IIvbBWlU+
hu3FnhB5WjCW2C7QFdm5U5NH4yt3MxIOdJTzsFwB9h/iS7/wYVeM7cbYcBiUpMmt
/Wcfxvxs6kzAArIH98eUYfomscf2kyuqNXW7sEWEWK2A9mgWXAqT8f/qV1bzBelT
0lbSa2yOYduioNXyu1I1OU4kZJ/WSiqhdOJ7aRpmkNzHSCP6Vg0YO/MwEi/oEXeH
Cg9qsfhdzhWbeQtvTkXXhQ0c5qz10Vj9xa1hgnsq3zxULJ5gcsshACvJXbtIviE4
fXjpBrW8P/gMy5NLONCGNCv3wM3nd4ZmggCjBdkHm0hm3J1nW4urspJ36jjsSHlr
oK+cxCrKjNcnAgFhM8qphhk2DmCqxJLFkJOVmYlKqDixeVoASDN8vTzzAZMaUftL
5TJvZ0MEQS4Vi0KUmKhgscUUtaL4LjAdB6zYn5IhDD9IUazUDdd2VzHM/mPEaGjl
60DF/AWKeGHHJDh0usMTU3pG+vz8AXMPTlqf9qqUr2TqoSR2pzmcAhVGgKJqLs2q
vIXRL2Du90yC5rMa4yfKcCbF/hsRhqjUMZu35UfQeCzxBRMpd/s1Mqx4jZS6OgUn
Xkm+gtc1wwUiEuJtlri/PtW9GfbA3MpYaIEtBIum3BI2aeNDGdpBNrQwv3B0qbG3
OCh8vyXdvN7V2g+zAjCTa6r+Vy4qok5ZvcjUJSNUNRdsWPdmU15nrh2XI6wJyf+7
Epkrh1zDji6JtATLzwP05edzVCCAYoN6s2oBTyJXgYIIGTZiRbnw1qfVWS8lJCo0
xzYrILKDuJjC4zQP524KS6KbKXhOs/ejdoHAllW2d/8rWu+7b7ySwUV8ULCNfjHh
SmgChydK0Vx/QBEsVCkdgB0ogMCOCNQSWZ5265zTBCVKqvjpp4TRP2WP6bYHqq10
eCOJM8i0jk9XZh4oA0BnEGVlcMHMZtQhrEDWzAeMleRzdVxZJkgdcfVy6jB/MCDT
W/S5xEo7fC4q5idWG4wnFCxrxDXqoExkFk+zXl5PuCEpbyAudEgZNLVEfDGr0X5p
i2Id4RuXFMVvjXITyRMRyvLHsakzi/WXbvuJMOCjLEi0Jb0216Vx7VxD42+O6Ri1
FsseHxJJxWeqElfDYmUxlikhkG7sJGi/7scMswme7bDlIAewA3Ugfx18PcUOeZze
osca3bIMboNVEcXSp7bHWn6DSvQt2i3rddMFnhZFrSV7TQs9UtLm+WNkfclBvFCl
vmQatjPX2Ar/cnymPzKEtJSRHzDDLA4+JP+zm7cH531gVX1Sfm7/BZcrruQLzray
hxQEnz2TvlLKyPKcxJMrSVxt5wKqcHdBbsotUbIqD+DT6qxErtFRaYziwLq5eHmm
Eu0nSmqpywU0MULuf25DkqnIvxzKrUtD0lIhhqKb9A7P/qgAWCq3zesibYVOmDPR
V+Jfsl39TTADX4Z6T+KOpMLe2W827atYhop/ZOZ2Y3uNLVVNUBUiHU8f0URzzy07
alHLOILFMepSeVRjP8NR7439rX6YToCOVd+kv/Hi9Tne/mH1K937S/Zf0TfbwBMV
wTvweUVpGdrc+K//MEjLAhyTm6ffQ6dG48gpQB4egrWFK/9nv7Pvb5E3ZyU/dpCX
NvC6/lA0uw05369i6jZMpl8Pz2tcpO0kzXIu28+qKCCO1gQt6LHGb3L8HlA+jCz7
/d/R+GEiZd7z5VelU1Y0cNpbsg/Ug0UbdKHZBx/sOhCa5x/Lx0CSUyOJT9O4fTIO
rd2HCkGKGJ0XBKGQg0XXV2V1iyWsO8ZMWGg9AL2YvR7GjsqA5AKB7vWhDIWkW5yk
N3hX+zXjynia+9PbDcmnohaSucE1D+CuU5njLildscsAchXOz08RDLDlrNZLPkyr
PyD9hNLLnliSzSdtVQjcw502k4qyNt5eULnp1WNC8XhzUZA3xIfiSF8a6puFEisY
BGlz8eyo1bauObOH2I1yU9SlG/5L24zTcqBHdScrXqmvEG6+0urYijySVmLg4tYR
60z3GY0A7CEjTMl+McHFE6p4Y7GChl5VN6piDyb41u50XFnKLvxQ744cl2hCk8kH
Yy94jsyvlaj7KHoFyrYM7GloLNYNAXqYbOv6PafBdovvI8YTr1i47b+MI/H2YuEF
ZcfytnxtiKxt84JHasDPr2HRrvGw61TQmpsdnan5oH4VsRLa4XCOa1aEiOvvgCOS
mcPqa50CLKmPwyl8DFm3PQdX8y7hdcl5KLfaFYHxq9S8Cast+o4Vo+SjMivEk5ys
Hm0066gpUeBcTVFqO8L49ro4xYIMpcW+hAXjKhZF6oDHyOUvqPbqr/eFvv7lJyKo
AwgYJG1RoyEh5MamoBgRjk6FXnPkX5NoSbbxYpLGAAx5BV7JlXWrc6nR59392EVZ
lmFSjwaBL4h9OFGAuPcg72Ea8/VZmDsYt0b1BDbBkI1Hx4TW4cvJl0Y054aPFO4O
6eRBNY7jzqprEwP0phv9KfjsblTjSUpDmmOKFLr7CETzdIgnJDDGMA85mapYnKSF
+4FisB0nulSO7myDKqaUXHRruVuZZ6dRDMJtndlEo8EFgXNyAtLTH1+VNPfGPwsq
feeek3St0mdQZEvCMLv+w/N/SWMwwVWMN33N7JJdH/e7lBtmxFgxxrJZNO63pSs0
u5TpRIe9jrOlz7zt6/nczzyKqqUfMP7eQ+pkVyB3x5MfHBUEUSBwELuzN2W+BJeS
WBj7v3jGUYz1M7/vHuoISTzsvVGDuq2nZRBreWmIweqOrFRQIP/aAlb0/MW/L2DU
KAjh4GuqHTRwNWXCgUP57yD0BnORsNbF7uMAEqBKEMSlSEJTQS8LUNkQ0GIqM/XX
OAkijfYSsmTTvpmmFEEZNUeBkEdknIKpERcJR93q18dAT2zSMguDdnESCUKuI6Mw
boH3Rg9TFIXOoAEGAi5GNt7lwp6gZWPyP8IymPh0RRlgiw07isrem4mst7lRfPq0
ee65k5uqhrOeM94gmK7Xk1dDv9QPtxgVHxlp8ZDOJZ0tOTS+FpdC0pcA9XVzTbav
p0SpbgHyU/FEyt1KOiO2dWLKlFJuC4nJan72Qn8752Y9kweBtNHHj8rJPFTXRkQq
U2/yMX4u4EIMDmlm37P/sHGmcRBd4isujvQNSi0S0LeBNXwtsrl9sJXm3vtUVGXT
GxwD3R7ItKy8FV7j6cTmDupE4iCJ1VLPXwEpeU02MYDUKGFRX0Z0pWZc6ogoH9oe
OTQvtQMq78oguojNn0EudTH8r31VYrrHZj2ppc8fqwGtJI/HK95D3mQWWJGf6Qoe
hNMGwpzZY2mu2Sp/jC5wDUeApZw7Vl12Hfb4EbdnK8x3RpoFVie4taaFHgmIBGC5
C7UkIKc34VTmdDVCDv32KeZl8fYrMQntUWfhOAdsMUYEyIlwk5qOPhMn0DHAd/jr
ZD2oKuLScfrQeLQDERhf2cU4P3PFQb4ap1scO31+xKRO06MIzsAs0uxdGK7m9ck+
ORzoPv8ogKU+DgpTy21WZn0HF8aqTM7x1dndI9lDzmqAWFd3zRrYdsOGoswl0zGn
LDyRaWCJfEh0hpgrXhsJ5kEDelje8ys8IPse1rRN8XDXl+6SmoMf7pkcsxPSm6mL
tj0NZxfoeRqFxTmg84yKNUlq3aeOVB3U1uW+qsIBoCVPsA21S52ro1fAJ/+PxLky
7giZDtmMV3ZgTdj8/PaabCDKft8oELML9qo3YmkxmBXCuu8PPGMUMO+6iBKSI7Fa
DMR9CF9EDGYnU7cD0wE4A1yt3DRLJzuoNHvGoppKYI2JJ+HKEOgZhW++O1K54PGI
vndyX4omGyusrezT0Qn8OhDlcLVmkyQvhBAOVqTpmoGzcNYSaDpZScBTN+Z9r3hy
kxvsaMl1nJYXcKYTnOkJa7iBEKPa8p6DMDyWkCFywTkQex6BwoAt5uQkIv2lg5Af
2rH77ipVi9QUv04ZyjllSHUC1zC4EOO5I55hfA9nvNm8CUqv63agvp5MhL6bFfjh
rxf9ZPQHAjAOiob4zHlWrVF3ahhTyqqNVv6QB2L9mEPV5gcRAe4Ca/q8J1RpQCm7
cbwchoCOi8NSrPtsvGkrAqYA4GrjkNWrbl1k9dQUrf+IvYX55MfFV1mOyiF85WGP
kSQfq1LnhtaYbAKVbUSVxgw6gT8CbuuuiUzxYKd10QhpWC88JPhf/cnq4VoLy2BH
894Q7dT0kAcqNVCcVQdpcoH5s56/ANYgkMdWzodLAyNtNlxNKOmXxBEt4ekLPAHo
1jthRaYkcCayvPHSQpk0AzKWIYBieSaqMjCK7her5qHeRFEb/tLeqrdBerltsAOq
BXRVC8uJXEICzzzl9qfxF1YsXtVHHr02ym2v3qs8AWlI3em1VFErGYqVG4lONFOm
SaFV8IQdVFDZtsqLjM9mEHr4J0tziGaKyBjmHIHANwtmQmSRsLtiPOZP3ZObRrND
aPJ+QXlF1KpkZUXdc76AyB6zB/6ET74Fc46jeTxSCmjb6a2bF5CbR8tAfUbp6QI1
aHrxQE9rJXC6rnS5rngHz49iGTcNo91LRMQ6dF14jcGSr8iuChQX5kPAG5GmPrA2
LAZto3MjsHxMtVQMcebr4kriPoSmngy7mdZZI0TQLzR4XOLbZWD1l2XJYwRqBbhV
AzPtWfMNFVOMPce14a/YFPJZN3zBNajKIGgEO+h793KRzkToq1sWq+Hs+gVmXIbM
MU1SAJgp08AARGn8ZBvztuo4rl3xjWMlsahjOVT53StuhbN5ajCAdIyB+pc4+0cm
Kh8yxJAPJUiQshk6n82vVwkUDyYsfqsNU0jLRzBCJ0DDTvVUPpdBXNxrVR68Watp
4+ZvDx2l0/dTpHYUF5RZG/3DHsziBq3juSNwz6twcR/b2Ad+wbMgmnkkXLrp4JLK
U8pYs/8d/C+lChTNvR/gT/yW7xHUN7UyO7NHJYhIlxGbo+yP7uv+EK9rMsp4HrOT
W4PY+Jc5ss17N+5fFsoBStG5UW11y+Asf16IDL3G4v+VzRb/VKmHHxCE6NTeeGA8
tuG5/vSV3cGBrEo4Nler1hbqzVK0HWhob2IEs9+PRAkcpUjgpLFrVFErjLtn5Jl4
DQvOksyugMubyok+kiY+CqEM72yqmgaZQpKKc4xKtWWBFTRab/wh0IgWFOXT0Ff6
fHTDgk8RO+LYkEJSIW2Z8WbVKX9uXUy4dep0A7nezWe3oTxgPwCGu+KkR4xEs/Ko
wpaIDADOkxyy6yo+qo3KYm9zjygzDwCqBqY/j5UNWwiEeL0/Aikj5qhRoYWkwjcH
Xlp+wmoQcl02TNqbdpS0wNFj4aiuTyHNoRIhm5Q1c4TJkTcJPa52Z3K2O+IkK5nP
zy1ZnyAm/Tm7hsI330V1mB1DX8VJHRQggk1OZc646CuEKtY0E/Jm1BRbkKXR4f3y
EX0h5ZdvwVyhw3sX0owpVGFygS442gYlKChdLLLwvd+Qn3WrI6PtoVzxTPSV4WqD
2/l7piwYMYSUafL88yTjv2gmB3eiUR6sjX2a9rtwDgCkVF6jPtsh4MWYYk8Jky7n
Gj6imGCReUrXJd9VsBX4Ey74RWWPV4BTgyv88ZRC5vvDd6o3VyGzhIQy2WbLYdi/
k68M32J+tWog46xKu+ho1rKEy01jopleMwu5H81xCPzV9xX5MK+S37tYBHDDZwQj
eqE8/awRkGNU6npqL0GdrDSnok5lI4tTuzZBMTpUF/zpbnsX+Tz0xVcWD5FWkwcA
gKxrrUlaeCkO4sdMT6k0cMfH61tKSP/bd6/JKwuxp8b/bLAf/RnmHhVLcMmZIJ3X
VNgMjl0fGymgMF2udmpzEyFTkk9VpHQEpWtuTQk4ybFz2LcUZY7Xx56ErjSO9a7T
xCI3+nefo24QH2B320evKeSPp6z8eHE19NZ7Ai7e8odfQza0g6oXhMtgMKdwGW+R
0aCF3Kv2qaGU3zco6Ng3H0xd+0xkM6WLE8y8LqAH3+8G7+EkSU51dJ2SDaahnSh/
9U0RNK0hZosszuITt6tTygC/Pq8F6SEMKot0C7+HfCzfX3Nv2OPJ/LQlk2tVC6ir
j5VcRn6ZpBCmQZB1LbS0yIZy9Dtwdywy2OgAgR89EmR8fdCn5CBLxIivnY+hJYHw
qGYUKJctf3pGqcA8vIZC5uZbugMX85u1fWDIfohclS4UE+74t37HP+C+CwkpkzoV
cqxx9yEsBtJXdaGOag+OTiJEWk7MeO9PX6ZgWYwKZSnvaZbC4uNWr0NjdfscsEtq
KuhRSu3k7S89HEBIw62SJQkJZOwekGEQ7hKkicVgmUIyBIOdPDzIRYJ7jL6hV3ry
Fi4g3+TU9iVeZbxmMbm52ONGPK3pJtA9s6W0DgKoyOWqmtYWDbAY061d23B6DbzC
n8Dt/RqGTIfCfoIiBHNV4mqZOlPwMjiobH8Po1xai/mYy7m0IhcN5VIdfinYYli+
5nIOBylXzE/MMPwTBWOwqjUeMFzS0qTgcgxR7XxBQ/vcKIxMW0dyN1/PM2/4nkx+
TzcXCjjShJgeX05dtkiq5zwBqim7ch2NsYvK+lHPQzYSu4F/8k3ldSFezlFzFJio
VK5ql52a+H5Xdk5D02Af4P9OJtjmuberHhgkYkmSyL6swHngQ8ROOYjh9rDC5KlZ
EsNOvd5ebV9y9bbVeI0watDnKRLnItqMdyFS5bljtWmb+a26Dk15XdK+DNuk7PkY
06ePE+BO0C1F5jxvTbSDoStOtqYgHm56Bm9aFGC60ndh33OPkulzgPUXvn/NOUOQ
ahFdUr0njornJRsptIKW8qvQlKqX+z33ZQ6SrpYksgZOG0aJrF1A282mevShCEVK
ykfxrp7pDz/CYIN2cJYiAtVXX9NWXHNl2CPN7lSTiCDGvfRSxp+1FmnQsqBghsur
n54xCtwD2WisEyondU1ptBOLh/qZhfrPtlU8y43z51oyQyX81EqWQ5OoWN6kPXz9
7LSdnGS4icabB3SPHmTZRoJOf0MBsyzH3IxRo236sSGqacQOiD6/3pHLQDIvQQL1
su2Eph/Cy8/LVoDZN3Vj6B1+4UpJIGLlzzPw0JHEZjKr51v3I375vTCP1y39J0R0
o7Y8zfkAcPCG3fjr8J0AcFNCtSeA/c0SqwvCq5EC0Nyh7aysCkHEiEVJBT11UmTX
3qBmidvUSJwf3dLdyst3Ld9BlfVGpiMfQOM2WNRzCPfd0P8tGTPxqYodvTrzXyp4
p7p3CrVt10C1ZNfhdS6foBR3AR5G9h7/MthvIHuvgNfmttfldgN/OaKMBGl7vATl
MBf+dkg8MFbh8fJ0yOBxYZUFLKqqmCow1yloDjFRNkVF5tgapDKkOvYmdKbdeXF8
A4oWv5ol7IBH7t4h90zAmSr/hS7mS+YOtQZkLrj0c1AcQ4aFRc4RrnuQVpicgqGn
WivfjtfsQmsGN4nZAE3obVWSNqwNJVRjqxxvUDNdbOQzktcUToGTvj0ukGcTdO97
QUXRpvAC4kawA4T18kEKlHFCJRYZyBJLmFGQd01FFBABgfKuA32xrPdYQQ9QSpQY
C3w8Gqo9Nv35Mrzjaeqzwkan6ab15uUCgwRXmOHJ0MmBx/qXcF9vBtJIsWDD2Gnu
yqje7lyXG/1ycQCGg6FIKF604N/jjhoXJ8DSAmgVLgGWH/JM1OXRcOxuOywSKuFQ
ahN8UC9Lv6ExjescXf8QWGcNIjxg2LqXwp+Ep+uqGNq9MFfNNEdkY7vh7YGuEv2z
+9Qm8qAIuBK/6e3IoaYijheUuTeIPsnKExVhYUGfnwD0UY7RPPwpDVWVJzJIvGe7
WMcGk5RfCYFWMTJ/ZWO94qxZBc2Q+z3uFtPjrO1YCxhDZ8flsxfzldMhU6i5F6Q9
5qWpxQE1oNoTXxU4qtgeaQoXrQJ7AwJy4wTM5uxYPbkjhcukVf11f0eIojMXF8hp
GAD9fDqCGREFHZjWgLKfOXO38kpbLZrrQGdntRBVXv7v012c6hfcHSWlmjz+0f80
G7kYYTdb5YbWz4oXDSYER4S/uWsrRoFklo7J0lizEkPpvzn6goYxbV2h+e1gKTAJ
Fo3K6ty9G020HudcI4B54jdQ7B7NZO+I3fQ1ulI6ssnqomoMI1VlMd0NqAZEsiwq
W6PQq5vesk2rwfFI9IcOqIAt2cYUnRbtwL0AJukqInST7lgHt/LsQYgmvmlSOFoX
388du3MrEHZLylop9akOSIHR30ZBSJrX/deTMT3rhOcn51yU0Mf7qoYJyTfghr3+
S/OROnTHGHYpLY0EHj3QY/utVfxerhHXKa+yMhtmspm2HkmxB9UMMebH699aA8Fa
l8XhvTcH8lejVt4XvoUl2DvnfyEKe0+tj/lyThrIAzMMAU0UgDL1EbcyXqn/3GPF
6pD9mP/TTSUkly8vIn1DQVQZtaoCJRWW38Z4rvL6ER58ELjnQdUxtHzV8/uhrcsD
L+xt/IsrXw/vi97KptUhCf2Pm326fzx2CVt4fQT/d8d8yvRp1FB1ssFvIQs+GedZ
41lmpQYmiJ//vbMYu2t/jTC35XbkSEOG9wS2orU5CQPqbCVbCiMz5/4NR3RGn452
wjU83M4HcQQMVkLmGjzZXbFzuzNW2YTYKB9WOu6SGXpxG3pCXrbXHw0ItsvOKuuN
+DDEm0MHZPoiYWnHrK7lCBkzNtr0evhYW8pXmsgI14ha11IsK91jZJNoy+4o4Ar6
uayqjDnbrck22smkDgJ8oiKzHoUWl3216K552jaVzD5Ts4ewuH35EU6TLo25uODC
rvozTVU6fs0n/ihVue5ZkRQr1yIkCK+z4dheu23eAFLECt6UbfQSW88Kxrvt1d37
rDkX6YJ7rnzFzJooTLqD5OkmXbM3hdO55EyTQzx8Wetan89srOkUgL+IXHzpqbnt
ZBv9o81dIg/FFCQY6FLKI6ACohAfOsbJyj/jiZuqlP7lxSjglowc1fQ8oGcKziHU
+U8DT4uMyBB+KlD9R9sQVVt2HD8/+eXZORkARcDAIvH0KGsJz2ljcjsmeQGvwzds
lvD+IXw+R1M050N1jXBZe3VsYw5P2JilJhX9haMe8OkUmdBEZWV4hEzyIsLhgXYy
AVngoTzipYmRPCL9AiaTd62weA2qTZw9t3HH4dunMgZVJn1L8t6qExUQcOlBVi4V
LMND/Q03IskL+zKMdsUCG66Ql5iKtSeYo0kF7uYyD88QCCLakYaRcBIeMjTLrSNN
4JGqf04RHF1OZH44HgkCvx2jLWa7Nvfledw2Pf9y64dP54BDNSWwcTBaoRDkzmC4
OtLIVJ6G8gt2Fq7T1v9AMaO9KhHr21/Da/t2mtSSTJ+7aMuWQTu4QbBXU79cUIW0
Z/fLFJMdrluRzfhmzM1DAzB9fl4o7Siew7In40e2FOdOP0GBO0fd3+Wfeia8W8rO
rCs/Bmq0GPj89jIyfIgSDoFQzMbG29K63ZL0xsXTO2EKv4Oi5IL8WVt9Je7T16bf
nc0wSS5rnyS38Mj9d5bRPCsiKBYnFlBbra/3BVJFvG66wjyTYEumcr7jLZJXhnPq
MuH4sCxcsCUpvrcgk2UMeZVOfj9PPu2gz/Xemm2LPbtLmydLS0Z9TGKcIBoWxnuR
ktnA1azhqDpIX+hpL1BodF6gRRCxvVLgxY2VwPjF0IWzXbE9UqO3hZO6tTDoIotx
Eke9q4PjtDg3J4hH1xWbP7BEmUkEf6lOmeYdOU0rpCmRXTt7bWwNZmYnJcNieNbr
+r421miJ7O/QEzPrHUscje3CemWIg8iPJwbZGjEp8RybXA8fBCVCJpx5c+yCyzP3
KkR1TvE/f8hIDTIsB2+K5MSETRG1uLJHAC6tx+q9h/sTjEcUxiXLuy5fzbP0w8qU
StKlH39q9G8FKPwx/AF+TcUnpL/yaO66M9AflF4dzcCOqxopqeOHCbXSOZyqAkJ+
/yBtUxu+Ss8xU/lZZ4g2Vocd5lhJvIIb3rLL27jiXjLBkRNyxhPEC5/udD/T6mkt
PvdaBl5IDZelkeo0xY0twb3oxsL8zFVicTvFdjqW9DgRSajyQ8LYHdfxQheGqhpk
xN/SgdMC6NLgoZFgdAIFNGpQyTdDvB5NNYJiBxLD7HcpLY037sHXfP49IBTEU0nN
nmNuybmU4Aye4KAw0u6j/n0aJrEHrmgitu3j+fhrFppEbPToIzI0ov0ZfXAFqeEA
LiABVhLfKeY+jDIihZsL1agw8jvuWl/NQzoBrfwi/D93pYDqjHDzal7aB5+q/j0f
jWFw21Eb0HNrKTVghjBoRcZwegROwsG1oQFCO5WPAJ2Ene4PhYlqpYIeT7PT9pkT
fm9sjeluqJtdqHbEFyK89jspYPqYaD9/TZib+mNEIoKIin7tALGJwzCoA5r2VrUP
KIqSO1OPhW4td6LZo2SowIHXOCyVdPItQrF5GhiJevssERZTYX7ZBTzgwMIHHj5L
czmhMi24gRqlU7ZjT+JqoOKCnUT8CL62aTteMYDeeE3jMA++Bz12ga5A3O+pBlED
uzXuRVBDNSc1CIzPe56PexwvyKpYd34HWc77NnzV3gC7yf5PPs95nVOMtWETM4pl
bs/UT1SPcLyv4EGMSTyxOEKn7zHEmfGvg48fPxGelRo2pMVAwcMHkoXa0H0XjVdl
x6cR66DxO5Cx/HyI67qZtLOO3r+svRnuW+2T11BG4x1jDt3DU6rMW2jqQvZP6RbA
s3ezCYGSgx3eRuPoXnTW0ZrAX4AiTchzXVOS07ezeCdFuRlICRn1VBYKwzm6+c/w
nG9ywAOiG6Gk1jH9Rd51j9REBL8TnKZZZRN3ItgvQMRvgZspypoWMkF7PZ/IhQrc
BJUFl/DWUU8/lWAXga3sLZo9UiQndbnxPKrTgyYZPRKiX5BTAN9mzqPtn5Jwc3G0
XET4tZoBJAUOMfsH/S6byCIx52J+gLdjFClUzB17/u7Cz02anGyRfHYEryPIR6UX
bEde4n3T5N+boGSP8vLlMs1f3c337nXaNpzU8XPcuv8nzFSVNER/Ht/fHBBm+BDX
bey0RLTCbQKb6k2OCYJ+rjQw9L1aJMIglsVysukFvEH6V9wD+3UUL3w0G46lFqzN
mRW4IZBVgPEoNfSuP2NoxNVuE4SuBjhg781QrS0RTI23qsv5UmQ5MrfnXg6iHd2+
DyeUp5E+d4WoQ7ckxBRl86alijJCAuZGZW4XcyLi0z7gpffFGTv5nDxkQ9qMtZ1r
+bW3X17tbsqWfExUIX33CfT+/7ruLqrgccOPQXUkeVdgb95Uu8hjq+MNypYinzK5
kZol/l3rbrI3DBrwbViHtJTeGUFnCnYRNYp/KtxsG6kIPvaFu/iCh3cSMsvk0AOb
7TkFfifpKiCp5a/91U0yxKBg+2x9VUL5IBbXmsJy/bHFd1HwqLtP+0mctX8cHleh
IvF8b2foBBQYmrHhjwEsjPXxMErGissqZor+jzPQppcSb+GXkgj98vB4OKPPdnfG
FKDgBiNqeGpLIP/sP5OmjdW6852zGCaDzzSNZC6RalYt/zAwJUwdk6lRmRwpwJuW
cs+/UlHZkdPLVuV/IonbZeSRwd+KWQr98QeVDnqTe1TQbVUippDYiVUIlm6xNkFE
JKPaHeEaVuL+u7l662gVgTT8dWd7+nXSxQE68ovaC8N+vWxTPFi/O+XfHEjac/iw
AL3zzsqIYVan1AjyU3zgaCev6StmNl7Y6Thr20zv+YwPlT4tOdE0DD4OYT10QYwi
K+44Ui9hdSMugXUjy/fgZCoT4Nx8dCMhMJsGt6T0MqxHASum2C4fSQlRac+HYC4X
s+GNe55rxra0iSNwmVYmX2v020Dn3bEYLGkdFDVP2rB6KC5GKflxa6L6xBaD/for
Oa0nYsMrrQUQk7M38gbODuQ4s2x7FCzvWj3ka4wg53prsWETf0jn6DZsDFXVHDJy
uTJOglOgF9MXLVAA8dyYIoSjERvIY85dFzzgboOZ31WQra78ddERfml1DlmeaaKu
Rzugfksa9h59lsg1VM/GHenYfHPAWxfyQ3B4dwkzTDPO2xaX5b4ArWeIJrIzKMC5
UaxtXhiEFoQFDLT+b/9lLIQSyA8tmL5wE4Gye7cw/Mu4hNZTES0dIk92mSGApRPk
waUvW3H8EMENB4L/8vDqcqYjeeHuNVDQVLk3rrnMOjXKZWKhpsZHLCWJ07QIPPzr
8sXfEa0GcQHyD7p68eCOeRjGp/jA0/E7c3Ooe06OTw0P2dTLD2zJNm0LUW0aqlkk
RG25eMRvB833WpJO2JE5kaXMQmsYhHfNiKZlNvNkBVej1h86BPITa59tHvPlzjGK
IZb5+M5IouJH8Iu1zM4wbabwWj6xXiDQKQZCb0N8LuJ6AuSwbJ0TWw4EtqozbYVf
gluwh4KSEBaCG0qAUxhtS3T/2egJ9zCDb4L/HkJzUsHa8TgALHMGmG8IBoNAsMIe
FJqMpVdDA8gZnig7Bdm7Y6qacQ+CZjEb9JlLUy5kuei1yL7cg4SKqwht0KFz5dgL
czJV91yOhhOinAw9132y5/S2rDjxOqnvZAyXYyo4hr9hBI6/GHThn3SCarTp1EPY
XEti5hhH6PeiW57OKJZxnxRt5TMjx3gLNCN2HG9DarEPPMm6k71uvyAJq32NsWvs
yqN89UuHMFcTdCik7OvD7U31PUxlfMNXR95iWCwYkD94SeZ6EV038aKAJKoZ+YGb
pvHIijaHuWZ7xaJzt4DlOAEG1PguH50E+v+rgkFca7tG1OjeTUWGUB36i54jfV2J
Y7xhaKx5aNRDQL9BLqPyuPuIHFjUHoyl8HSQxoz7e1FKLLywWBEP/iBcXKYJrloR
k6tRMwry1Nu7K6HGrvhrDx/8LalSTOWOUzA7VwZHvh3v+zgBdreph5gTq68QmNmt
8tfjfLqh9dI0CjbM43aNq/I+bSDXEy4F1177f0vEv4Ou2T+9+qvV9uAGwi+vl20o
VpimlFkVTqlX21bNqzJ43IDM1sIl0/ipLMpdY2GkyPl5mGdLhUQUnvW/GjPZvX32
8qu27xJM0kkwliM51cdlBQB84lyZCegAJvLlzwd0puZFuwdpstrWJJzEhWO6RcAs
MVhQh8UVpsubrR255Z5oBKZniGls47hfpIdJPN+ecTfxpX3GGG7PAncLDZXUnLIx
FxhojM3PlvUJJO5+5o/w9AhdM8l30fyRVibFX9DBh1LOZe0nnyCJ4DtMdO+NWTIv
jZ7qyiWdFLS/XL7K+99EsIJTqx0kZqR2oYFbBf/U4fwMKCMrDz3/G8MR6VmJc/gu
+5kb6d4IfrrRnEh5qRkw1/Zss9kZ3eYBx//ufzJT9MNrkhnxBvH2VyIVdO6b7Hpo
Y7vBqkEqpMQsR28gRld2uXP1UkphQKmyJl3FE/q5vvkU/CO2MC25AUyQamDvyEyY
e34cgIfePZy/jiscfcZf67MnZ904J7U8YSxVnJ6f9im+AaRBFBn62uPvFTGIyDxk
txqicH5wVMhOI3TeCOHgLWuJUaJf2QM2QDEfJvxmhgpX7cichDQDIYraT5SQHcFX
gYxjY1gRVH60YbaCGHoo3FQFuQ5wRh2f2tVGLsvQ77x9QA07gmv1JAm6FgtY3pmc
ZjlpVm2GwwFTZ1Kr91xmlRpgYW/jyj6I2MzQEH7Slb4+M54wkFMmXQ1dsgGiH7rO
GonTSMMR/5Lhf/d5Hi0bp+Z2p0LPYGLdcg01SqG9xZIuCSISb8LgiXO4TBt58FEd
hntvPf0EpXiWIPI6GkClJlLCwBwkXwLEuw0IsgVHde2GhhqBJ5SKuZwgKOCELzHG
ZOZohquSndNbn/eI4ufGuQgYHX0mWRhcjWJbagHpkSFrGVohYKZebDZg1BHhhbxR
lqj4NWcNJTjdSmh7P1TIX0/7GJEW3ZA8I6+PgrkDx7hR9yzlP/sVCfYnuoE6NZaT
TadOxdsHW10/beRantS4IKSLjDhrulQD1BJorrktjMlXDkIvRW8nnlIlza+UwguQ
8P/u15K0Lsdspe5Icxg+ndP1JFUqF14+yUkLowNopDIr4yFQxLocehzZa2z6lP77
OutyGIX6/yDoGqBmp55fFENAroS63+uSjIqIBrxpsvmYd259432OS3OdyLLmVSTg
6Arcnwmo5/PV+/vDxafJiTRwcGix6WiQ7RiG1WK3hZZlAbx3OcnMOfOJZp5i5bNQ
r88NFEQrU6pr95YwBjHlzI47OMoxp3biNqbACyJRAxuGiZ4PzuEotuNihQWzQDR5
hs70FYmqJa7LKJNBQzTMdkDFsL+wJJ97nVsu44ZcovDeLqDmCqnDoy0eEBHl/IJV
jNwcqMu78Q9p7KK4dR8Npa9wr27ZTbng9GvAtJ3l3O15bd5aKF4rxRAjnueyYZJ6
gqkAThjSoPhhnTfFTn10rKhXdGCq+zaqnEdkDjglOKlo/bLJZAnYgW7wjkEufV+h
e9OgKn6BotdbSccpN6mGzk3AhzdNUrkFu8BbJKiIZ06fDnWN3hdsEnsY82MJuIq6
XJIP/e9+zHIKWBUFOZQ/1/8fNh2FvM4k1I2wak99Mwp7kKV0mM44VoKi4T6A3OdB
VR7ErEOBKYgDrHR3T8czcE1QmxJTt5A+jTdNCs+NPaLqffvO3WTjUe8vD3wgI+iy
+O8RMZ9m+BrjhXw/y8BsQB3Y7VfnT2wiDrc4XJ+qfiTPWozdWysqjJewr3cLuGaz
4ZGr0GbzH4S2KPwnb4wB8ia2JayR0DJNCO3lSyjD3yhUGFtzURardKyEmuFwOw58
o4V3886dndxPdoDLy8iHOLQlQebBlMnl5XyKSCJVJq37/bNWMtMmmQJJGJ5pOvd2
3vz82pEmVcHxXTLz6ZwGfmGtZAMnlem/cbCO8DypjMU3qeqG51Svf7VOoJD71MR8
vi/hSt66BS5l1lbcYgEsiw9LTmwNwVbf2RY+5p8O4lZQLM9Ah0dz/bABGHFlqVkj
YfOg89ULiHBRBztW1a7f9qyU/VoWIQHyxqICNJ131poid/5VWOgqn/6cMISkdHln
M93ZUja83M36PPcVXbLjI6hmjNMvkfVyW7NjNVKrnHZJO5RIHEl724ack9OpJ7fv
5Gn53xet8b2/W/wicvg6nTnQUjwDqYq0EalQCvOCDWOEC5Yd4RHEFHv/XuBRdY01
hDbWlajIMKgiMYaXZ3pqxEjhPGmg/2Xd8wFNwy2LzsbFhhN3T3T2hJPhcWsWJ8Vq
iDtHymbjDAvZ3UA5A6hSf6u6vBVtqdQTB90dM5rERgHzbdE40fWL4rqsVncAx5R6
Lz/+w58l8b7lsDuV4+Dl/lOe6nGdLFG/eNebuNvAvCZ/yTZNtrdM//p36oQDUlqi
FsEtNgIHR9fHVTEY/PBd4e0sKTat+KUGQGqMMtE5me5cQtSoQJDUZ0HGIbzo0iH6
FbwMXNze/d08KzdpSFRN6ovWp6zxPxVrZViePi+5UcMeNCDWBGvSm/NpFkggoziE
FEtBgrkIcgcPgdhBySQAHpirP/hBFIEE2dYcvpQ8EAcKSvARnR27v0RHWUrxitzL
OE1N2o1XB4aPgHC5n0xkNelVX2s6wTCqCR1sF68Yle7pHpgSlLCHwijCdQRBJplS
Qcsk6IkcdSsuNXV48jEeY3+OUmFjTBXq8YXnGw3i0uakONOTj9nmVyGE+/UkmFSZ
4Tf3F2ceqPOZmFxhKkv4dTWCXv+PzJBIgphkIbdWyPtoh9lb/xbjyz3TvS3ezb0a
DY8QfocxICgZoEBWwKWxnzywW3DKr3ddj2ouaUzSKxClcb3+F7cByiT6sJR1RvcL
/yW++9Xb2d8eT5VvABIacqqegwUEF1qvkkiYifgAhoMsXUYwTdBq2/yot5jPltDD
tMZ5UHurX5vA2bpWyhiXucDhXsINqxSOOErQ4TIknkNwYEhuk2MRJq177hJqroM3
U2r8DDLB6+/AFc471A4nVZ8RumNerkaQeNAR+/Eh9ir63dMu40DN+8hFBexk2P73
9McXSd2cBkw1aDC+bqKLM6OgGd/nfviL9cucNmMz/5Ylmal2VNZEqAA0uqv/pZjc
je3olN0FR+vece9ch6DlocrEBqM3NxpLdYaf1qNhPT1tIrIobnpcPUNyNgNLPhyk
6MKjh9RqCt+xjIZfAF28Wcn8s5lxPK/4y3u5CD9iFrPrTxMAZb0vW3xkXzLfIpEH
7IfaOf6R7GsLNCoRN3GyIgyTFlQk6vvwxx8sn7Smq8N4Rg6sj8eMzwtldUypDQIm
wkWrgHnAM6lmUTqK0dHLHc8PAuHXPyganFaeMJkUz2R9vmY38b4xiu8WakKDuvQz
3bdhJCKNhtzS5YGSGuGlNE8PmWP4UtQtWe5lwuHNWcqA/3tHLDbYQVAeSasIzmSl
8qe5a+Mie4Lu+9PD3P3ZWr/6FOfAKMXrDdNGZgWRflNTgdHeiiCQmRIQXudZYAkK
odgoV/l7u0chp1seY+iVVaKY+cMwCsdJaR57Vx+8fV5dS82l4h3OP4Mw6P3ZcGUm
uUhpI0jR6YC17jtOY7W9Eb+8pLea1vqYgraT7lx2VvyOwYhbZtXv7ddAo1/wQjI6
45xqbAbXyFFR6umOoq8YDN/H0+AXIb6PFm2JO5MUppEReG2S5QBF0TWmhhS+CtF8
U9pSrqT8i9RnIQbd4TiiN+IAR3ANqCbi9Bf8RBoni8MbHl0p9IR+emFHUvFWLmVz
Als9KAvPE3DKRvZ9Zbcq2KPA3l9j339X/gO9QTcRpJneMUIaOrDN36Ae01E2flSj
55ujI7IQ7rosvpPUWX7gUx091G7CQFxVxsE76+aHttDpZPnl8b+YeeFFAq12qCXu
3N7IOUYcFPP6bEMCGh2EWkNgpfH4RQ52ucEGYbw43atrEGNdQX/W6oRKYPiYhZ5/
Ka1W+tSFB9DOoln7N3bK6lZ5HdbYGVbi4qk7OU74ZUYsV+PmJwFGkgUu+/2kVKe5
MrOmB/J1b+L0ZVScWxL9HKlnebNoTYZsn22B5RPI2jOQS4ydsrcaCG7W7Ahf0Y+P
UsIh8mlAPRkdtBtyGvL1buU3vZ0T4b/JkB6xwD4UNQfy2tRwWYhDPD+J4F8jbVY9
eJbF4wQDBIN1QB7p4nqWGS24BVoYg4O8OGQEgSyj+0vTQ6qUn0fcyYAJOW0JXvvR
0NcUbCsudhvGa2KYa6/DqSOS4rjHpWfSmOQ6TMvWKTb66z5xGQ3GSR/fGCe+6AlH
xbvUMUXuzlGU/8Cs8GbsmOBnK5JxqVPuWIlCdZlzSBc347tnWKtL91FYncWqPrgO
9tAY/zZAAX+SbD25OxExlIirBCdXzdkq1IE+KCV+LJcHFm5ryF6XucURq2T8Ljjp
d76LvAYdz4TJsAmdJ3iS96nzHhUgSG5XL0BZlw0OxcbW9ABUbeGZUjLv7nxlfxzW
9VVbueA4z2cg3LL568MpNo9zpH7r7wmgQU3sMVN0Yhnh466fbA8dFie1uwiLjRkH
DV1kLChkej0ASqH3Oh9enHcG7QapVxpHMMwgrDudcVDAHBYjBOFyGfmjJqKs6ilL
YW/o1/kRaHN2ECOCx909v5Kb0vhYvVK4se8WXN/wOraI0Rd4UMEmB/D8ywjOYHlv
Amy+Xy35jN5CHEaNgfXUHnE6uH0tsW2gvV/IXCgMUhFTFH3YpW/d/YMKLdgbcJu0
McziVGVb/ErRQaE06Tg7zEKsBPDH3Rqy15HSJBlPBud8kvi0EsU+VDMFHC0aKDMx
OMW5yrGFjULhQr7qvg0AVZqe8RCfOnvhkkWJt1sxwGM9Cgw65IrtAVJdbLW9ER7a
bfvaV4zr4TBUP0AmjF8tQnTMVJf6jaBZrThaGlDj6FSLXQnK+/wjXDxjhSX9X9ML
D7YTNWWAU2zYRTlBzYyEVpNFHHBaPi2oVdR/YAlVZO6mN4Cylsv+rgq0ATd4T18/
2zvC1Ps2LFvdHqeY+Nuyrv+RW9QhOhYDo7oDL74d7sZ073lnyWF/RVfZfNxKp7cV
VYo8zWPDfMOAIkePlah2MGWPLGTZwIcKcGQ+nyesm2c5YvFgpHtKpUj5BPwhCKVY
K4A1iSakTTrte3TloKDrUf4YQ86UbXKBXloeTjK2MDhu58mErfoPOMW5TUNv6vlK
z0YQCvQgd7DDON639qxV3OLGmEHq57/E5HlydCFR26HWtamvY8h7c/pjoc1eGSIp
oZ4WyVlM3YXf77rpf+Lv9A7oIlS/coyVgqpFGk48IsUDjl7Wvtu7qZHtnVc/mdfX
E+S1TDp/1yVggZWWL719BqnNHv2OFP/9ZZ2n3TAdBFJeiyEBLEdM4onwvR64aQRY
VB8aYNg8tu8g+SxS1mtnrTQZneKCUmrEgSYKjmJHlqCdw9tx7OyAOmP4bJxzCOh5
T44IqrKfMqx3geLRCfMRc6NATuxMzN/EFn1b5GzSbT9CRCDNB8/yIMG42deGqKfS
kklxpsyetSRQwGDppnsNhX4lrX19GXxgZIgCWAqdzic7sBGcQRNdVL3vnydwHR6N
P+Ae+OZoyOn/dP3rw5oSqzj9IwhPGdQlmIm5VFeu4sDda2eYCdJ7Bnso+MvLgPED
ZIbIyl4ZC15pgeQBO8t/BniEVH24TXnVMiXynPYKZxVoOGrpYQaMMMavyF/iRo45
oz0LUvSakIIx7OaNW1WrFeY93yeqOsYY6CdEsun8UKg+hrDW4HkSF8fcSgCmpWPZ
9577W9pgrY4sA8MfaxMFFI4tTvLo1C7bdslh3AWqklizSkgnmeaso4oj7nkF+9ig
xAPatcKwZHf09jj8F+16dVA/941yHpvwVnjcquxTSTONe1t9Oua9piL3goP8V7qd
n8PykbRdw41SdbUEZMdpXx6sCJ0GGlIR3baiVJcPqEyH/9Fpiuin4DcDhwUKs6Pw
M3miyd9wiQEQOsDWPZ5TV8Ne5wqbvWqw/QM+4L0RHwT/Eoxmq+lQcacBhk90lKu1
kUuEyiTmOiMO2HwRNXc528Ommchb11OvqAcj5SPruonKNgGC0Q8vc8mRi/9Iyxri
G6qtvqKWVByLJRsvKj0dvmD4hM8+yBEBvKYbtr34xk0zqUcKIpAN8KN5mx8glquX
dSQwcmfIXlXh82b8eT9bFatmbsfLqlg0XMPJmA89A8mhXfpimXqTwYAsK7S8koBP
TJaHYa4X5UOJ1HwGvYiDlkW6NevIPKCZc6X3BZzKmZ2iP+TR5JJwaVYkPvW37ZxU
20yOz75xpGTeZhH4z38XcFscrtyqkufJnCelVgZ7u3pa89qDJaeWdDAtDtOPW359
O7oSFKQbneC4XIeZjX/fj9ocOzhcIqpZZm4LJNIgXXmWa4YVtbzC2LCn0OY8DwMJ
v60uZPnEJh4It4vHmVtU+r6cBrdFUmoR5F2YMcjJsth82S8kLzae4Il8OlRHbmBo
CUDyio+SS3gzrWzcHtwzUfMW77+CBu9QcEOasY+5v2kPRsyiC9WlFe5/66FyQK5o
cyNAnQTCaWjZGR9BlcdpUFS6dcRAuRDoQSEhKnz3yp4yKrJ6EtUCky4cAQd615Ob
9qOwCAoI2SAAnoFS4yPnCOIXJIyWphTrWqaJQ23lUvcGdF/8gn5fPQ6smx4n+XCB
h2ViSSa7q4Jh5ALEu+31ML8cqVcOPbpzhVwjYzmRc28xDBuo5WIcs3izBusLDr3m
2tKaMnpLgiJlZUYkAccf5VWVkAxEFAR4d+JsElO0aPiiXwWgJ8CFJuDjUxpNi/qH
XSbzFfPvUVfdDkLUv34upofdEBNqn/wXziIvr0uTA8EcpTJcQcIN1L1IwrqK4dWx
1P5zWqTjaqUex9xZDZYqmKmT6ad5Nb8JxOCxInmd60sst0vI7J2knmKPBEMK3Qsp
7gy5xjDqXRktUMQzGOiWFnBhRzI7gTQllW63LZfH2mvXimcQqMnasDDjkF4/fCfz
sFXJgfYr9enP0WOimOLJWwTMIKg/E/sV2B/Hy8TTIdgen3gl7vzBLIKpjrbCAqcm
koJtUbNDRgzzx7cu0pk+1+C3uzqZGQmqTeQmXpqRWIX0VtP1U5n2WetU6UzzX9je
ZyPcBtCoWA7uXvwPZwrK6gDspPylMEc/WgGcT/PqHJiv6TogQrMIGB3o9CNGgKlV
Ju/UEsTK0u1QO0zwkOLUL70xgwsAhphMRVsGMuC3FPwCDM7T0JnYub08eiqPoH5/
ewWqylMqW8TlP7Yr/65iaK52zM1RNyJzuQP6j7tQlAxNulsGzh0fFt6XVAYS0o7c
/3jREWLPnbu6fNdA5fjalIY3f6RVE5KAWh2NTBZ6YrzReu5J3VixMYP8J/oAOM/I
s9c2hLmcKOm3yup7aR6Owpo6zvPSYN8wKflvZNVSfpNKBzOWi1iUIOU3874vec/g
36Tgn4mEQN3SdCFPfw9QXAEJYF9+grLZ79WEb2UZLgzlUWyhw/eqQgW7ugOLysrR
Y9HwGYq0OoVGA35ZjQW58ZkG6yolwsaRXNZgCYiEkMf2mJUrZ2aXv2tpon9uruMn
BVdl1k6MTEXboVzc46V9J96iPM9aerfI5UKYEb3XXm4Bdq0/FIX50fcqRCBj1z6i
WgJx3e87PWz969gtMJ9iw02CiVWFeg0PJbwGJpGPLSybAb2N7AaHC48mNXW9omt0
x+vxTMitzPTdX7bc+caHlLhNYwNivMIN2p6ws/x4ENe+3B5IpBDJaEcx5ZI6l8la
Hgi4oCpCewJtwx0jLJWrzK+C2/D/q6Vb2Rk2vYMsDCS51FjVos9YabkYdSafDZ+0
nl11T+TkyS6Q+YWOiNFtMoxKeGspEuieb/QgwCYD9upjZNLeH6AO47TpCvQHWlhp
Zp+QuWrjkGUObmbueg5u/m9phVZGJQR+cgDN4xfpGNmpx1JFZQFz6cX1bBR2zWKN
cFc7BQTMJG8l59YprYlEJDlj87MRYPKiTrNxXf5qxqdCih4ThCrgQVuTjqbhEhMJ
qDMAnXeX6qjyRIHedO7UcdF2fu8k0jd2Krm4hIoEuetCDpLUB3OHOAES81aQHMT8
NaznNzzgwPTtc6FB2Iour3KgYmK4HU+eTQRmPJguidppubnGYE2RNubcnCyqbrF+
TDLhclUT4YUsufaijDIuhYLiqn0EFbO9M9osXht3Ao5GDSHQzf+lN2/fVJeVVsq7
YLhKw/sB76AocdhRznXFmLkFfJJ6GSAe53bq2DeDKNGUxLVKYFS9Ig0iEzbdhk1G
ATup0iP7JmZWQtqIy6RWFtdY6uqFhdJivoTHBgGhPUTc/mDwvzrPuHCghioEzt/Y
K0xZlj27yrIg05Q8kYRkxWzkJjb5ZQcDAxfCB8cY1yQQ3oqvIubJieosJRUbydgk
C5l/M1wGI6/iyTRdIqS1Qq8+ezMV8kqWIXyHEcPcg8lmiUpTzIvhu3lL9SlsqTYR
3Xtd5FwbrrXsBuQcfGXNwUEeZWGOnH1Cj6XYNrVyY5RV+cUcfG7DKxkkNA2iwcsW
jeAa3/U+xchdg65jFUdXBCMQmKks7vljevNXmyJIV8xUNwV43K2Q0IK49xzyo+od
K9KGI5UR13+V1+jjCb9GtE1LJAi7DAKmAeZHp9bA1jDU1VoSm9xDU+XL3OrF64RJ
xpO814Nv8s6jlmDePyUV/kIMHQYfiOh0GIj2AxfRu1qW8KE9vW5NHue+oaTE4rA+
W+hoE+IMDrUK8QVfcUq/sjhiyw1Cmu6svGjytjlL6N6vMg9q2DBm5bPjh0JW89O6
nspWndArli/bO0cF/gA4qERrrtLyBHKNG0+VOIbIvMZdasGKnDwgsrHMrrTWKKc9
c1sXukNNynr+ImNb4weLRu1W10LM5zhCaVNUJ8TXQDvDKeVov9cFyJoyhP1zz/ni
kKJoqOQRvRpJXtuO2/6n55YhnFLkNZVCCdIJz8+xO3fTvpzspXGd6hBmIyQEI6a4
RJ0Pp7nAJa2A3WbFjLEtthjfUIxRtSYHLq23IVEu2X4bVsOsHtAd55tNCI7WYA2G
PWfrFCi+8fKSZSGZC7O9PhEgPX4aHisvsoHbYwI8wZtNyzr1+fLC1IQlJNRYiV/j
Cor6+AgsDSJ/JZtf3gO+OxhgjZaEFODYXWczxNDt2nB265XNnORzHTF1gUYm+N4U
+H19BMVRAXMh6kgm8jZA5buzSbg09K6adxCFsmynuytwvbNQq1kgKjAUaWnuGWmy
CWlrXxll7VanMXE5ZHShvkigrEklJvac6/9iTf5RQZMm0FNtmgLW92SyrvgUPTCx
fjvYwSUEbc2bgG5JAmkaKqrO0Rwh/IcOX5EyATe5fEnZhjnztm1os5yJSpIEikmO
bA3rZ1b8xDky8WE+jbvxlSqzgDFUzkyRmw8tTKFjsCduWzzhp3Pgh1n2RVOBTATi
9tUSC228oprAuq5QsT/id1TfDs2d7WczwNS6duyxWHMd3JSlEzW+/sA6lfQPo8i1
TgEjFITGJ6EmoEjnfELtTjGqtpsymnGgQT1AdmkxTt9D/lWPWUH2fb2/tthmv/sq
kD4U5JP0wBfRd4XnnVyB+woeNNI1S5I6PFnbmDr/KZhx5Ee6dO6T4DITjDW7IpVX
SgjTrGSRF40hC8X1w0uM0TN21xtWgk8gpUtH+wxOrHP1mbav6bK/0llqgRRQB/pQ
fhEA3RqTfK9db/inQXZmCnK5w8eTiVN0WEwPJ1KlNuCtnXT1UnMOz+DksplhXp8o
sKqUj/F/DTAsAg75uftmfkuko4Wt+EWtl4g1HRuKK4Y7gfaoN/ADW6mY43R5ERJf
EQ5IpRoKV/L66UmkuKlaZmHz/nfeu0yIbYFh0wg6GDGg2AREAPETmcbP/QfrHNRt
GKVo1aYDNJ3UXYWc8ZZATA+YKKT5mHWf+DtfO8JDhI6d1O6ujCgSAPiEb+Z0RC8A
rF5BbwQitM1hxeX9v7GyicGUSxeGjXWNG/oIBsYlsY5IVSEsgH63N0CJB1aRRBRm
hKByiCmzYuseu5qCTZ3+2b6nT6bmk7aF/BLS/9aTaAf6mE5U985oVXaNMLHuyydG
wCCGU94azRdD/d3HDtf6ZZnlg5AIyz0W45S2F4Ip82TaNad6fd/wfYjigX7thRq6
upK1S22VIEhtkISF7Z4zd9gWh8q06Pggo+LTgZH6FUAwVN9pYDlVZbElSH4/Zd30
nEQaCqTPeOdJUDYQU+gmC9k6j3lrFKc7R1coLsWTin4A9UBTa3plHyLcnp4GuAh4
166v0qlxCUAn3MpjsmVHUY7nJkDuE3a/itbmKMycg6/ETTZPNrp0PvkluAybzVea
cyV7f1IaUxn9tb5AJ8iSnpqRJVoDjJP3wocHZ/8WmCFvAyad6loxeKZtv5hVN9YP
+jcHr2QMGU4iRnu+na4oDKnzMIiIiiQynJOc/7dQtGQtlJIg5m8UZOUDwYqmzWaN
8ZBrbfAySGOswBNDMCtcv9eofGkUZSH3xsnh4sS3iwE5DKnsw9KNMzjqIRrq+PaC
MYHWlSxZ3bvtZyypxHDstOFqG4aecZkfEX8hZOA0wgoDS7vg9ryiLvNYpCH/4D/Y
Fs0fIFyVNQUSOK2h/2N1P0E6SF8qtaY4UXwMnbyjLcrWcqBzZ9S3KEDcUjoqcV7I
cR1xK27+AIXmk4I3gp2XPIKAyfIpeubxxmoscFEhOq2y2dOYXEOkHb7vgDtbEGhk
eK1NN4XXo62o57pdR+D2yCwOrm5rqhVo/50lflPy81jBLaLvGxn9pWheUGE3lX2W
JcKV6gYc6Q5AVS7dtg7yqwe4zrMab8xHixbE/dHpX2xiQ5i/3PnhaglajMgjJmCC
0ZvwaJdBe/bSQbP5m7gBeBb6ezLfwLyBLLim0dztCos2Hxm9A9XCRREgzehk8b/l
ILJHUwtivfFCZbVcm8livDPoZv8/uxlK2ESUR/zohtW49FK1j0WLzyFlcDTZqqxU
md8pC7SIfi3+pYDot+kyVjc0alvvog3RvUJ3BVNsq7AdavGXtyNpGG+Cx4RDzYyV
Wvhhupk9/TIHoN+3snL6T+R97Hf4YKSpsde4mEXpJF5Km6tntfTs8KVVK1t3I3jT
YLF8O61LN2rtdkUQ1bXb0dYnNiBoPpoxs72cWCuApLLUPr9apofjyWfxOfS+Uc0J
8XqFwCuBTfaZJhT2g1mYZ6pFUXlK5jKR7FeiK4d+Qxj9bgDoaXVh4A+VFMuyCxKq
4omNv2WEzxscGt30L1VrinalJ9fF7JkoEoFxNMN2JS1RMWAuoPQfFmTJcFpHirmy
nEelsHk8PniLMhSCqiQFI744XmMtdctb74IrCgsVbToT3aJGlZ0QeacEdtYPDoYW
O9xX6i8DcT52ebXWY57lsbXtdXRjAUgbenLqu3SanNM1KdeeNYyH1MbxxjPGu/XF
0SXEx1wrYxgZnO6H3mm/0xMPjakjxV12cOr0t5QSFq9MQZwv4VZkA1zvMAfUrzSr
Tn6r09b8J+DaPx3htPXoAKHqeHa24JhSVq3j4EbQn8GlHzt968frqH0YktINjCHJ
SMlOzDg8+Rm9T0gP/31L/5Ny+3EGpM9NsH8g1tUI8XyQeqFZTqe+hJO8GxPjwntF
IMnWnLvgw5Ai2xZ6YfjsOyly7/3Taz9jeEIBlADKgQUOvUzYcgANZbOZ+KA15dls
LNojHr1vPBPt3j5eAQChJlFCmucf8PNXbWH7NAksUnAh19dMrToISAZUM75aftaD
/VyKg47/zXwrPRcmwW4m/e2PwlLQ0aftyvq5kLoFXw7Afb9KMqfJSUxEbfyFLZpw
q1McTXVyfeJvonXRRPBQcAHCpAbm3W19OvrtcrQfM/wiBHaAcwnyKXfWsWpivIZp
jJiMn0jtbhCiAh09CHtFf4DD94YETCA1XR+0MG9p7r2AVlc/ULsSf6bIPtpEx/cD
6UQJRuQ3j2jSTfRl4EhHOmHPVkoLEK7n2U3D5sMAz+3Qv+UTpr6b0IwaEvGoNyy1
JhrlXitlyaWgFLuyve1qzTarJ/AASjPWvn05vaddh2qO3PdgVyp9wWdA6JE0+TkX
zJA4PsZRRFqvBE8t9HWXAHS6yVYtS1he5ZWyljuR8lWOUuRbaK4x61Bt/XFvIJ87
bLk/GN9NOGRSVzGYo0ROOZHnoiSsLh3hi55TzckYIEXDwWKWuBstu91KbUwFYwqV
lhS6n3VHUJebSd3bMFpn1EO7Stkc0kZdvgobZlWsl8n4ddn446VdlOLobKYWWMG6
Wy5eHKPLjd2yICi2l4U2sKvMlJvG80nUKLEzI9si57ToC5cwyCR9LMlfXzRw/iPr
d0pDzaLE+niIRVqkes8NoxVtHPMWBXnB00oEWN2LQXsbaiXOhbgsP2kUcqjSKxYb
ztJDnRsrWVFvgnaBZ21crgvTkfzdEpPK8sci883vh75uiNVpbpg07PkFwJ1Xp3Zs
2nwt3UMgBsvDf/NKr03fawqK9WRMAX4dm36c/XcxjuLkJS/tQjb+NGU34+WxZsZZ
AqrTkRrArCbGfUbiEBGUQh/XW1Wxd7vIkJvSDn+uj6LAXOOAnPBvcSqdMAnErNI6
K3AQTNQ2OUj+8LnaXR+bvKdPIzHMCPW61zZ8QzKalPTF5aMKWk9+qFxn/M1XR+eT
WHENAyCaCAmsWrGYcH/wogWgS81oEVBbeYqRd3L1cBRjzI4U0husToxCD3XYaV1Q
vBhha4sWW4FGSZ7ZPqBmv6L8F2NNoAiTLd9+ULDboU8bxl8stiW01BLG7yooAEOs
amcpkAuBMtbx1Eoag0efGTDr63idWXUU5ds+7w4Ym8mimO3K8kRseJOL6yX3llJE
WwTV559prvSOtugOJ8vct1bbNaInG8VGYMxs+XiF8GjHJ41OEkWsGEYZVKoKETfx
bAxHff0TQU1SXKR6Rit/+HafnG84wm0sal8Jz7X8JF2mplVsH8AUIgISDC3fIvzx
0g7C7aLMqL/WEwBFHCmziTQOuah9iAZDzD3zw8g4MwG7iNA8SzalZgIn2f7HObUv
v2nUc82AjBMi6NK3u0vCGPjIQYB4r2i/r6NIXE73VXXqfyjJiMDQUWgOrpobjNE9
SMkqYyp1h4yCHGIJoUbw9JKDsON/AvgNdw3iSuRyWumG3SHuCS7gTSqmq628rIAy
l7IgDf3vADvY9ygzXhxqTWPmme6PFn2p6Uj1XHJamnf5DIybu02VuSwg6S/tK9/H
tw8H2adv6XoEoJCLraABykwu7O7k4wyQLghPs81kPJlF7hz5aPtF7iIdZy8tiqXA
fp3GBBHkQrfDJlY7uUeu6NKjru7XfkxytId6jWdu0EYcDmFoCKZ88MB0xSdUDzCk
TIaP1UxVMVy1GpUw7/h6ZLQdbjoylqOEpNhodMmpVPeb1WzL/7Mxhq88bAO+oYVi
n5KME4cHFdjDVqSeY4Z7L9uYSG/d4vFzVbZJVUIDwc5M2piAS/TTqqf+h2JljwEk
9oAUQ1tO48Zkij7UPhZcuYSkg8cmevPzug6W5ImMdIGEHje0JeL0/JeVIwvY+3fP
TlzR8KLmuAE/lJV/aCevhI9xSB2cLWDX0NMnEFKgu5Ogc4vzjCdYE6F1PuHgdzg5
0ybcnDP3RODhlR3xEEcxRc1AzxpWgwg5JaWDdA2OgHqLty88P2/FjlUzo362QUzf
bGTwHcWXTu4GQ8lova0PK6zjx5s0bSmkdqJJRRd6c2XDD3gEMjBxvnM35dOzYcnx
JFIXfX/Q/aYdNhOwVI2cWAa6Jfp3cCSc/1XRps7QzXuFmELe8BOF5O6TKNDLVgEb
WThQitP2yLsVA86USxbRB/pB3IqlaZIa5esmmJXGMQY2wGl2lEmxEf0+ZpeEG1k8
kiTiyeodNK62aJAPBYVMLwJzlBsvM28I2DMO7rTQK7ah5FAdKWVzIO7cO/YKdx8O
rp18jY4uIF/D3guCyoMiObkbgNnH8hU6ogBt7xvk2WADGF4C9Wx8/epC4HDVAA8d
lFFEnELKgjZIh19ijB2NHyffpevwBJ9m7MKlEw+VkJL6PB+QJQTCnLIT5OewlBWF
KCG1Huw/7w1aE15Akjz3jymXVkuIFXdFMJqAo/LiOo/0trjMYEeSzQS/e7bu0+AL
jUsCbUR6XNsewbgqoyaMXmGoXaBJQu5WPnBBPgpwIA6w+DsAxjzm5RbQWNA7tqMH
z6aSoJxJM6SrvTcPUZy8dG2JkTbthZ1hczfypAefHMAE/L6cGXwFRo9HIa40UYjt
IARPvxPY6eAaBW+GpaYHTo1/l6lABfukcboC3guQPqjSu/aES1Wi//epKP3DIlXO
fXOsprfoD5P+zpZiAPdZHkrH6sPGY+KMC3S7b919pG6Umm0DD2wgr+RpxYhyRFdj
rNIKrPFEg9pn2X0ns366IKvpUkqHrJRtCH2qY2EUFGCUb64rKHupkyE2ZOww74lk
rkZGS0AmaIpVXB6Et2yyr9efDe0iUSxzoWFrkJw4vgYM8Nk9M9R37jLG7CHokmPM
/2yTV7qaaBdjVhBx8zxkIIaqkAqTvpxa4aUUh4yFV/h9lDwx8xEkVeX3O+hgFHe5
ie7pHfCH7AZ0sQrL2ooutmqyVCf6hiACLm+Yom9peBZqgkDLVm3m3NatJO01I94o
/MjVtzRLoSqgpcMWy3WBfXGhRKBEdEVTdfI1aFOD5AfJ3m9zMHIZQH/uDcbKAXu4
UVsNty8XBeA3pjqeEz2fgt/vZ81KJJm6BxZNFKpxuOyedjjbjTq8PAGVSWF7YDvC
BEiK3mMjsoBLh1NKNJmUfMw5+DAezuhccCW0aJ1WklgHyKeinNMqFoHJRGdktxeO
AdWsYiRhy2iEEtmQzrExPt0wVxR1gSqzr0eEV2yaADcRhiNybXoDnH2s949Ab7Ej
OM/1tODa2/JvFxi/NuaGy0ELnBoqnupAEB+x0fx/WTA5zJpRJmNcSMJkntNCd9Kw
fMSZRaMfxbxK/jNgam5TwI9Jvsao0juhdH2kChsvfT6oMzLIhVqrcLMTJvSZiKam
E6I579P98S+pIAqB2ipZ/PpjbgDwCT31W8rebg8jb3spY9KOfBBDi2GR3UTQtY8P
E4cbLLsNv4fcDA3AniJDjUHOcFehFZ2YDqJIDGfIAW7e7biA0Y9KkB8tE5ufDjPs
TLLMdtlUUjMh5eryHEt3nYyrII/I2fRgJUEZWr1gj9vpAaXZdxBUnJTC/17kYkAx
uyLS9e2GGP3QbGnfMyC2XRbDvpJMIEIFd+hqcES9znobxPrZp1P+/rLe87pkc1Gq
E8cL+8BjsSgmz9vjhLVAhzkKil/5GEbqNxoWGd6F/xRP0xuMijlyUw1R4cHpRHkV
FhU/P1WDr4+Qh//7JF+UbxdyQkarVlau4oPpo74QtGRwDvBUA4N5302zeHEApqiD
AVypYiqY3rVYlyvK50rN7M1NANBYY+EBfKnLPSMX/5iLYJdL79IhPyC7XtmSqUCm
YycAXXCXAp/z7a9TuaWmuyZESuyckbPIIDSa1pr3VqDMmVygyfc5WEElkcEBw9+i
It16qYyr3kH+alwdh0P0+eM2SGAMA6+KJoG6d9/l1FEx78fJlp1+Z69TNlIV1lnu
GTSWt8csP/ydP1KJC77k/zt8c3CXcEMybQ131she1vya0cUAL85YiR2C0AhPjz9q
+OFiOHd0aCakFbZue1E1lPuc5W30U5R4KHy1bohyAWowDi1lrtiir+fcLNd3OjbN
Qe6QUg2++w3p7kN+9DIpeRCKbASMwpXf089XAzbpw4M54OA8s9n3HJoofKhct/xh
jMpfm8GPVxHjmTubBMkpPC8gIwgU/H7LSL6Gm6aLQDwmfvXsUfSVRyF5u6PpZj9G
eMdh4rHUr07UOgommKgweKhmJ651arLvLJB0LOL/3IS7oDyxDgIpLc76onfWLVKz
ofxVXU+ltrOPCx080U+0vNBz1sWgqEZGwLoW0n3bUM9D6Kp78EZ4tojvQw39rwRn
OLBNb6hYx24P2yO6Wk+Y8oC5tohSkXYnMdd82Yd5ISI51bRc7qx3AQh3xCuRxcFP
upV08sKAXAkYF/MukBSuZF9C/JmN9cbaudLyRyYBXnt5N31wYHau6Uln4R6vn1vp
hTkxCWIHm5w15+6n/8aKHLC2lYYzJl0ITfDLF9/oX2sUojRToETH+EFBTA7FjrPB
o7/p9UMIET5UTiOTv/dRo66MfRllIBa4+bNtjPz0oE/mOc373Y9b0/I5nSKoejY7
d07dOKCf6OXSN0E8+PpG02tuXz/ayUUuFcp6RFkDBHT1/9912z2oMWZgkSURpUh6
BPpG8rxvFXvPW0E+8Ru2oBGGY9GDyNkMq66K/1/9yKHWZ2x/ISkmboIiVIRaH5sg
/BXqMCIHVALR+eejZsZS+T3BuJX3J44xkvB3K+5EYLAUOQdIT8TxqfarjCJlzgB8
2voPp6I21pBI330zufFi7+dhiGz2FUg+ildr7woTeejBEr63CU00gYo7Io4RXFDN
9uGN7iMSqIKDkRw8DMxSP5WGUWk3zWvZx8Sd7dh+1Rfu8s3mmInzioJePeGlo0Vn
gxlpdkqDldtmqdt5R0nKzaAx4iAOzBZVK3FsuPGT/uqtxuH9qCTUcCOZzLBQ70LZ
ylV24h/asHwgiDife4G+dEMpQJxBtF8VUrbAYS8sHsR9RkLcBCJZ8m6qITXnLy82
5751F3us0kb+WA2R+LZv65PHDvxOJuSzYQlv2/v+9JKz1Zzq8yo22kHGn9HcVB0Q
nZzkcp9FJhipqe2pxeRk2OyxALpPY3m317ouzZGW3l7fz+gik+TBuS9NXa08HSLy
0sHtHsq2ab3SSYQacoCS9TZ+xmLFmrusJj+7dN7aRtsE432SaEN47kvC6XmcA6b+
ZFC0yHEOC8COj4Cow2rGKE0pxiUsPvHfjB9jeX8ki3Iv2neUsxkuSf9jrxErFX2t
xUpUI3W8HRzIAXjM28es9TYDizKpvvTiDR0AjWXB7sB0o19TBmeJ35H/QxUjUe+3
bigMZwuJ7EGWcHr7GPvyaTXoXzXlJbdZPK6vpWzpFrLWWznVmOhWAni8hyiPkW+0
iKHVJXza6etct3GnStIuA6s6iHAQ62p8krp8ePEcxL8UOfpfWdsxS7Wd6LLVr9cT
yQIIOsAf3tcvszOQ526bWX1opYJhQgMqXURQXSTYhtnhmvfp/BRUb6tsGDlvzyS5
D4p2rhnEr6JjPD0tUo0nJMqtmB5nhNFvs9AO/U6YceJH2ok+LdLeTs5G4GlXC+DF
29QVm/ICDPApUgtnrrOT9Y3CO11K43IjzvofRyztzIBLyL5f9XlqqPusJlpvmCuf
qMWxv4VOnbnAukBvENJAzD4/M/5qTatUzMFGqA1xzVrXBqzN08LdYuxU3IsZzcRN
XKzC52v9jVmvMxqUfqQSDqo1rKHq4/ZgTRTwBccLHI41ISn2Y3qgSlO6nYjJx1Ln
1VvGsQPY0nwDaHRL5o3o3VUN7KNCo5gVBKIk9C3Y1/YC6swaETO1aSu/xWw9M83/
ASK/HisnHITx1o5Hqi3uLkbobUvpXQsUVxg250j+50aLZS8ZNRH6X7i2NJ49Q2pf
smtUWnZBKjEM5a0nWUQKX22vPRzwBQLCRKdcM0u/riksVwCFpNOrX74WDXzgmpnG
BMqr8ccFeor7DF7doNzbCenSgBEUIO+GJjrqFXLbtVtH3LM3NWBfbsDg0+w5KMEI
2pIvnGKD3vamOqwqTHRUNflJ6gzcCiGsZ/tx5pyBatf6N4MQzRx2ez1y3NcKmY3b
WDC9VPbghne1bTSaiV6yX6v+6NZShZ6tZIlqX1L/8vKPU6Jt4/Zwm6VXtf0p/s3Q
tbjjd4ehYOSbCHIvDeHR3ElyMDxTtgP8O3X+TKCLabX/QA13FG/Cqv4HdMMKXpiG
DFGk4b9zs6TkdtxEM/UhJJPe5EgG06DMx5Ym3K5COQIDkf2/ITlHUufVmZ1p0KM+
IkJPU/pGLDt7DCgxCAFAKhpC7ohNGPrxhD309RzJNjRdl7FOxhCpfj+P5c47u8Hz
iNsS+E5VSnv1+WS/3al1JPIBTz/XuOEJEonAG2U9WtxJ/Nz9Jlm04xuS2TkonXLQ
DwSkE4Y5KEGz3DDkCvgeWgleDsp8ao0RVEq89qRLOhLW1jOvsuDJk29Vya+eGvrQ
BY3p/bxhOSwnZXRNjF3Atmmaoh35AU3WUK00ld8a7wh3CbNjFtXbfN+f5JjfxEY5
h7dzlK8mGybpOgGEH5xpat9H6JFkvt8p1YgDPSEIji0ffadeFWo1JJTpxWc4hJlK
YqRXavCUcUIsgUboK45lwvtFiw+UOIz/NvTPL/stJcss9OuevvisrymlwWDy9ZTL
tRHzysXmRenG6Gwk1pSQsVLbCsQQlUJCJu7J2behuTsk/4CJJmq0YzYG9NhpD0lT
9Iyxu/1cQOejYCG+f4tBw9GbqF+IiEVfxT7YN01tZYj4NADh/Jt80h9BjLNAQaz2
wVWB5JEvwhtZ7gSFg1aqh2N0fpp1txPPbKOcw/Qjcqa7mLC+YlxRdxToibAtJizk
bt2RICqzXVLFevHYwtu5GMso27oIV9fh4uztd3Dfq/gHdZkXDEkrmQ+ituBMnW4K
29nhnu7ZAVrTm+shqVmekKwwHkt36289PlatGBvvBrx8QHv32xuwyswKpiJeY/dA
iY/epwVUiWxjInQAvxq5W1/gVX8ws5vBKojF/IsSBvWeKtaF+66YlnbhvaDIp3K+
oM+4YOaP1p1fyoOiy/easp5RjGKCmIGs2Fsd0KDdO5KqLcNqUTMwawaOMpSzj9CH
n2KAGrAnKpFRRKs33rg5yrn4F3gITADKVM74GQYNYIbr3YodJpcTClemzvEltzOs
n4mH176kvMZsngQ8NW7huZlHuw5hlIjE6LDe9ONuuUrZxg/siBtCjqqVh9Nb5/fK
mxoZCJ17kENsS2UEpTYy6mWQ0T7s6wM5CjZgUwC45oAGka4Ur5aVqYYAZNulfdou
lU/k3mFZi2aEkr6JDVvWCrLaEqe2V26wuj3uhG66v10VwqwQs3XElRKyJ6TXMdz6
3eItQTWlR9vonV80bKs8i1C+2QisqAUZpQfmh8dTD3L3DmzdezxyQAaSwCDh14iE
8SjBMMHH5VS+EfauezDis52ZcxlXwp3aREsXZdncVEyACy8wlVizHUwl6JZ/YtPT
76TRMy9O8k+131dQIqw9myQ7uQGZWZ74BIEKElnzR0Xy/RTdj3pMqkYB0nwcTQoQ
oIGzyQmTHnkSvxz0lqLLsGblQtbXAu49pWFPznr6vfLo/iyddcigit1268IV4Viw
oD3Kasiosv51IPPzeLRs7YkIPhV8ZOK1WhzCGFxWaeplzoahUWgH/JTyldFME1PN
f/Sw1obpe19BoWMEWcKcgI39ThermEn43uxO/iACAMrajYKXmpUf5KIZJwdEfqT4
L5OADz2ML3GuMTBYhwsjISJ/O6MeGbglBu6PfKP3OiyjXNOC3yEF6TvWYTgy52Td
3mO1t6mkoUhC9sZn3opJkmuYnDFZoEQvOEw7iqM3IswKXIuWmUszUzqOD+BPbWDX
NTl3iNmQLMGLDT+U5YL6qsyR2zL63l+iorVNPZh/VRNKJ6AFdafzENcb5+ihKaXl
PUf8oBsG9myMBGOmVdzW2yeHdadTfK+Rw6TKYmzcSEkS9ANNXf8cfxEzi5NxUtWq
eUzmY7NvYC1o10F1AwGkmgWHioWdALV4aqSvS8REAtw2B7NzC1bT8R1RhucuR7yI
y/H2lVovyLqRyUS2w/ve66OjDFLW1+jXFyRLDIRKf4FKQTvOYXPj2/vomLZCqY6k
zdIM/Jmng1fPc4X1QPn7QhlCALxnj1sBC4asbPAxFkiJRyWPoI6liIuSOBxh8ku0
AHZ67pzx2mx7jt+4bsRoXQc3C8KbnDHCAqX4Z0Rqk6HnLA0QGlMjB5o670YVQWWQ
D9ggy5GRtre5K9dj6hBtXFqGlFO0Avfl0/7N1PIzOZ7FTNxe5m5L82HAoBWME9Vr
5Kt+GnFpqRmtmgpapaigUSn6twwscBWwQPLHZ2dbYnXzPxfsZgU5epq1yX1X+EKC
YpFfde6JF5OBcQoCfjNsR4od1NMZBQWd7VpOxt0C0xy0HdCXdgCvIGzrFkgdKrtZ
GGYV1GbMHWZ0Qekq4w9yb9AjSEuDt99ArFffeXM7QEMYPn/y6FfQSBJoGcY0kBHm
k4YabYoceF493gxf8Ja6m9kGmJaaRVX75XOWLpM8J82hfEkHDgXpx0aCpaARFlay
59rQ8ZYQAhS283/7pJi/QioLHb9UBe0RkG9So6kDDmLIUGf21EKtIPKYXWk5fSvy
T9FfaeCOZ25prXA71WDLyXYdPjyOoIyKkR2GgNT282aYeank13qnacbax6GEhRp8
3CL6ytoFSpDYa0vpwZoVz+3wH9eP5Bhw1yI7xvt7n1NZG6lS9I6YZ1ias0qY1X7e
dHMyC4smCZ5hIdfbthBnHf+rhKcIuMjreyLM1GMaQ9yYGVqbHg218l34fs3EWjNx
17+EbRfnxPkMPaAuGCx75KyOEPE61BHj/5qbTtkC/MMA8DMz8/8vQciTyZ4S+WuL
58QU5lYlvtP6GxbjqFSqYxVcw9q8GmsTSAqvGZNhrCWiVg3q0tiRjfvyvK5htbkY
Kw2OtkxRnWj6Nn/8qiE5P9i3d+kfflXv05JmQ7r5puB9F7uXr0qHVBTLogOU29yN
3x+VRf/p3a7Ki9gDNlFJQReNVXyDNK0DjfV0RYKn+SxiCSvJaBwiTBuYY2NyblK1
Oeu1P1gPkklqSWcyUUZ2mJbfEdy8ku6dLNMWD7wev+1snA6HA+1qgW/fmywbx+xZ
/bTBMoTEulDGJOlUClQcN+midj0oJLfJ3snX6xAIabPFvk6j9au+LcZ9yE1cBclg
0rbXWKhIMXbNzA7UPt0WUUx8Yii1EwNS58/0t/w66735cchUw/ermZ49chb4F5Ll
qN+mGoEMR2Mq9NZovC0IJQLRaXufS09WXGwO2avwKyx14DdQGwhWRxzlYZYStWrH
yS9pNa90TAxgun0KUTaLXqViHmCR/6iNj8Rj0yhoxom0Oy3F1WrUDQIMv/B0PDSM
H/0SCHN9uawB1N3n8dr3pGEkSfFGmy76gyhEAYJDtOzmw9fILT2kqWpIBI0n/8LL
jWyr1FonOdFbIyY1XTykNO+5YRfDdEX7IdoInxpz/3V6pRn6+PEv9LH2cx9mEt0j
NRnBIti561lvriA4WwvCizqFddR4nduRe0xQp1ImzLnBA5YbCeTDf0pYbV3btplM
hZh54SabbiZc/oB0LOs+TCaoYWHWoCe4gBpq7/a0m5wHleiIRCBQYNs43pUiaWHw
R4tDYh3J1Hpa8zhyCm5LV6Si3uxzTp8lNsIdARYznfvQhURaWn7O5pR6IcSn64r+
fqVSdc9HwXGgzcvpoDkiQ6drOMUmcPpBEueem92ik98qXIMCr9J4Y8oPRAtqUmiw
65+Vmbyp7rh5WQ7Elp7BSU9TDN+L/84M9y53m++9cAgmNRaL4Ddyb+Veqr9cjxvk
/cSvkar8DXyJlQwyxevOo99FTWZyZwFovC6r+QrDQw5pKxvwc0UhYT41Y3KGSTYd
pLHjRic8yBX0SLq7K2rqPV8cwYb0BH/fOXs72hIOjujvc3bJ4/wdKDKQRrYKfXgj
FdKlRWiDRopyb1F3OoVnKLbztyx5sF2Gg4mD/8XvQ+wTMhPOU7NtUrep2pif9CZT
PaZfRIJU9BwB6eIqWHRah6BrCFCm6pxC0InA0jmG/hJV3XDzj6SKmEzN24V+lsSe
FZQMTQh3eU/SJltJpMvhCpCEVrLXyWZfDxyQKnAKjhHL7wHbM24lABzLforbqXrt
RC6qcXTYiQXM8+jFjRX3P2VRMMNyfq6lNIq0pJHhDGZ4y7T/pwlvQBax0+dwGh32
1mIEGkrGKzvy5FdSES6iiAl4E+ZL/d8KQvE+dpnXKzVor1xfrWmFBZ4E4r+CUGHx
vUutwSURLF55MvC2/PqFVvuWy6stTp59teq3rnn2Bv3L2TShEE+WRD3JpKFKKgbp
7dDNbZuAhVNBrltJGr4bkPsBNoa72liW6q1xMExeWVb0wozZIBboYFkmZXYFNjgf
9tJYHPUfVmLGBA9cRHqKCsgNv0AFU8nBlvIbcSdwkTcrtUe4EaOSIT1fU8YJFWMZ
UQr8KL5tFuO+zBQdyg7tJj7e2g03pBExv4hrJlrOCllkqlYJBI/8y000P1wny2q4
F03hTwZpaNp5v6ErkqWw9GepKIzVtbbQ5jA/QcaKa0Xz5xwT7pys5gO2QQVNmKtb
npnFkpnbcgazpapOgIeJM+OX1FgiKR9W9T/mpvOxw/MspO6s/NE2vfdQsLMBMLIB
MiTiLpy+86jMxQ1sjPsyWcCxvlc8Oi/KQOrY+EhXdg0ubiMEm3+Mqa4T9iwDC+/X
HQrK34gEUumCx/3YKRrQvBJ1Ahsfc4590MdlzzbwtwdVQIxIZFDziv0gtbLQYunf
jNV5bbjiMZNmftsT6xkBHLwXSIp1bbTCNiHmxmgtkqUlXp4VccD900TmSnRB/DKj
RAg3l/vWQKJIRgd5dL4m7k7yZ8ltzuce0asHagctbV+X6xYKqIoZxsGaw41rWWpm
Jel1KFO5KwJnC48z3aQysVVm1x0qFM8Q6rN21JY3L0ENmu57csXOOzAHlGm16toe
m/qh4L4d7meu2gOvN+TeUkh9s5XGRjlYrUW96zy7d1Ieo1gC4lJblzh1qHu1SWvD
FLoMaLqqbb4vdbSi7FLwHLCTyzzfSfvJzOKrYlcx59PSoCOQVMKtqYK0w0o66jMf
JwuHzki5fsqaHulU/JyCtzYapD7R+nvkjBCivi7Fjflf3MJzaZ9NH5KjFeBUdm8r
e8qQb3kk8kSnK8XvWTmfyrv6/ryJvniywmcfzo8e4BFyk9GqPcMEDqva23nbcZfz
bj0Ik8XY1kaY7f2as5+QQjhDN7GvrTx4aQ3Sa1v3MUDLhOPvVck1Ske9anDJYkEu
RgLq6ey5lKLHfB8750nkWj02WyvBjwwFR5URgZi5PIY8Y880JLFzPQWXV5Jc76wb
UTS1StSNH1zrPktQGyEzJQCeo51XbKozQffKXtJ6/3FhRUZTS15gICBWXsE1qIHu
NWG55kOAdtvFIxKf1ZmR0faXUGTQg8RKsvHgFoYR3Q87Gjzm5E45vfvKdtl98+Jx
xj1RXwdwAg0tmFTloM09yawVkuJfJlF439WO3UTZ2b3p308e0FKJpi4lCg4Dtx07
EkFX7VTiYmBud03PyMFcwAsBoqoxdT4WhmzIC8JqG7V62E3Z2c312XuN6kxvCycu
+QtWrBUathraNB9C1nG1aDJWOVNmOpmm6Yn9hFCs3MQgVVBsPCQpEFn01cn0wmD2
599cNvho2QpBF7yDIJFh6pi5P5YUzs/SPnkbjENRBb3R5pe2m5XTfv2ZVte1NW2h
/6WauOVqx5Ea7DTlF2NRQZwmLcpCcAcQNdExaTKzAPkZ/N/Gi8U/o3n/bEQNUaBg
YWkzAO4FJZgVLup9qRjQlLDVE22jeqKXibd1fdWIIRenQU8M1uDJbf8Y8TDFNdma
DXFiLs+oWx8kmvScfSpfzfZPScqlG29UeQpDjHAY1dEWfwbVNjdmvHARjn5LN0Wt
p9LUOkJ0+gxf9vdskZE/iBsfqRiw4/PCFxGks44vFisauNU2yHQv3SWpHnvZGjP8
eOZxn74EV6zxH4Tz+lSKXhzgzC1bVmTosKs9PZSADMad5kQwlOLbPPfHsMI5RFuM
U7XQd3wFwbdbei1uHbwr+cFI59PV5aXWrsGzWXUtgUma6VbMg/Wr5KFAAJtMnXll
vHP+UsWjcfPFoXYXG0YhbQJ0p9DnLJH9kz+iS/3GkQChlpJ6X1bnC8RXuYKsD4s+
TcsXYQKFsmO1Dt19EnZq4bscxRZEiP2wIZANCG8t85KVA/ZLVfhmeFD0BGswzRGQ
XOeNRgWYGpv4Hq0APTAYqN+HgjgHYvdqCEayqhFABpmykMEzl5QVhtmMr9REyFbi
+ClseG/FyOe7DwwMdkT6jnbXFg+XEXvdI9QsND5XU8ikOCwBTCfvTjPiGazsHu/S
/SpTeZyr8rfjmxr3PT4JgzikWbsPLtG7kTWnXn+RZQjQm9h16I/GeCJ+F2kDPtZD
WPZDMhTGUOCvdwTXwWXWgXZPZVBLGwZp/3JuXPyM/6tBvzCI2N5Yzle+VSn+Wcc1
p9YbUtkZPFppyPOeJdhC5Rxfpv4zDK/BhkAVsU9lR2g4qS3lIHC2P0SofzUf1GQa
AyFAiLuu+H1NC/7e/ARPdh+A1EfVJ0EtM2ggOWXHnFMs6Z0Hm8X9GmXhi/KUK/xk
1B2/lf72zrmpgi4eY87daZBFAcFfOdAufKxKn9/tzSwe52KitqsxxOKBFdvdDzVA
rlRzRM8EroTe8A3Tspxs42Az27x9cnfWG50M5DS4fCzb+kmAX6jL6b9Is7IZpVc0
Enrq/AEzYRd8AjlCS5HrGc7e1W+HiFoYKKle/gKfjxS9MPS01Q9aF9ldvfhAADls
NM7l6GbvK7UBrV+pHdvwvUe6RoGAu95St8LuMkYPRTU04U+vdFHlRpMkzUe8W20I
aTlYqj0nsxLyH6koyn9jX5HxRZqFreViRqf4e8Zd9xWleZmUM4XVQKnyt8a68RNG
Yv9yd2qczeHo8/ySJGuU62ZmKRHt24IH+vApu+p9Oz8nNb9YLtXv8Wh00Cja8ee1
xrFutwHMKHO/HRhbykc9BY4rgqjk06t2Qb1VulMCBB0kMEykkpgW7G5fJJGuqXBN
5DYICrPOXkbU6gnXTEepmsY2lxvfgp24pQ9aFw2ixTGuvF+/RBFy/LMSjEE7/qOk
y2FKRWBvhIZ5e0JR6MgC6cnf/EGmwNuaQQ0ybwpOUrZeF0dBg86Xc9F2+r3FdRI6
bn9WZ4cC2JewLWMLOElkVxEfReyD8AUHDlfqpC+p8pi2iuD6aPUFCCPAI5NRqmLR
mMHZRYsU/oIx7T0HIMm1xw0EyQLUCm3OtbcT/t7L3XMYk0S4fpqqjlqfMTMYhOWp
mS6ND+iNUeaeCAy+wMs8k7XCX0ilOMHCl2uzZCdK3cS+5BAc/igQUMs2xYO78PJ+
iIFOcTAPefZ2FNjaodv7fy4Z4zRoZALTaUP9NR7zid1CGzaSe96L0uYufjWeH5GB
i2y2jkNPzjxpZ83Ml+QcL7rFVWypFO3bF9EhdyGWZCvL1Ab/OxVNv1xmnJ1NXiyL
wUFwXvgG56/ZSyZ8jeWByomrtZpDCTJ98DcmoDO7wlL7mdOG+sfG/WCPBbzWuQ16
CWUhjWWmswr8lrMjvSH3Ua/gpT/WyzW60cCYJA039iexKR4mIeHnr3PG+mAnywTw
cylDys3JPXLCAf4YkWHLL53XYolEGY21nqOzlWbXB71MPlMob747wKKHWadLYhyy
MozzEot0eN0dbaQEbANQy2Va96Ov3GQDn8VFcXP8S/iiOixBDWYwsg32VYbAEFhH
uCOl+w6Xdch8o7KCuoiRS/JjF4nJUwrdZ8HYZ3FmBSqzGnSHsMgidBC8w9+huEZ3
OfAjnpHInPN0HZFAIA1hheiztDqCMe3Gjw1p/nbi+f4BbXvb5aH01vBnWzVTNScH
cRa4r8zzOhUbiQtJB+3OVQj9JC0fTphh+DP3LfLoIiSoFjECyZ3I/AzOs4/3COhM
D3G92o8f5HMxd14kOsOLylK6riohi/FeNg1qp2DjBbcPL+xmgbOkpkdO05qwy+8s
pHGZnwyQTwf+gRyjN7/AcdDvq+dlP51sMEHEUGNVQxzN73b1LVlZG1+Gr3qG3Cci
OFf+aoXcu4v0coAXX2eHfKxbO06/z2jM7KZsD8DztDQrh9Z++XovvsxGDVu1OdFS
nODjbaZCy9slzLkP6nEEloiUmCXBfKFh6YZUm1eWTYnA6md95rASqSkYg3Nke8Gb
RCxn43X3HWmeEH3NgnZWuknOp4xZuwoqMfoOBT43liz/jVzGef9IYE9y2NZom/Ax
PiuyrK+LHt/n+odcXR2cm8ZUmh3J5klm5sDa4seKgN6e38n6YB6WG6aSzol+3UXj
h7nizsPfVf5K9ifXu5eCt0yFiexcjsdHcU0onzcc9f2pwTSSWlbzMIutIDa5WzZj
/VXEDHM2KHobQNtv4mWJk2a/UIbeF2+7+XnExGBbZD3cVnVbNqU+JAztyoSw87Xu
SZ+rvYInMrOc//dwvZZGL/Fj3XOL8nMSyPHIc4wdeLaBC/m8KwkduowocjHFuKEu
dTVll0//zvBvs1vDhJ3TuHRIw1tsD9Rcqs8/vcf9WD8g1nuX7xQXPMnJ0JDA1Au8
LUvNJZzPHmECGhos121NWV/M/H5zYlKLmGrgblTI2b02vjnlYYz/XCBf9WhR5I07
9k1vHPSlGyF5aw8yiOQDcKxn/1/e7Gm2aE8yrC4LSay+Ts7UDuFHKxeW5ZnEhxBJ
Xbvz9D3i8le0uMlfWN6UFB4k2A/J3StgXsVKQlYhLrjZpu9SdllC4P6nYdhEjqIL
YR+JYmcHJIFGfnxo/tgcdb/3CtXm3CEZpGDo/aoe89wGffXBY39hivaVhGyYmy2f
1NbgjmyFMTpcGL+NZWUFPUDlaAteHet66T4UFdDp33SwGJ/gdGPaUAxr/RK6ak7S
SmkocfxdlcwtSLhFFYzxRtCbKjZaW6A/tLEnYH0PTC2OJP4FnOqFRK3xqpjb2gub
NRwFhAHLTStAC2/3Heyil+oPSALdN39w7KfuqJi8OLpXqpvu8tqVE0mf76kCBvK6
HtYOZV0zgmuSk92UbLkbfG/4bBjMITdRtSKww+XP7JWajYxFSen9c02JXmnvtiac
J7D6XG2AZGCpJ7eg/XSOEHfuomfvmpgdCsBEn6yolJt3MBU9JGC1BnmilY/9Qem+
B6aylpl1LrPy0umHYtNOWG4HdOW3yY6iM05VUJVFde/aL2cVjkBS/eqQnVFB7ogb
pl0NkHY35VTENyc1SVlI1k+b7nrhuu7vUcm4bneqxC4dkLla9ekHA9azhE0dpO5o
XyUL9QizqYpLR8XSe/0/zCAUlMqdCPR4Tf9kbJtZaBkm3HRwL/odfTMXsMuBMLPV
k28rUs6Saa2qCflKkyIIfNrwBjoe0nYzX/sEB4LgfR7dnBUdwj0n1A5YtEpEzNRI
yYVGgQYUXKz9/4hBf0CZ+Bg7Ez9cXoXTUsq1KplZhkWpzm8xYXD5v9b9UwVctwDO
UUHWbG0/Zqn6V+LAOg/GTf4N8GmxT1a6nrnI8wv3PQqRbRguSzMUz4MLCOAiZ9sU
9AbCCNzcOZHt1KiySh8xsnN35KWHIPa4ZcdsbMZVtHz4Ga/2XZEAF001aJAUStLA
n9bJ3BMOj1cexvhVvDhOdYF4LC8VIHMm2CEs9xz6xSRCEQs6odTpxBNgJvPsw3eE
ZwaNPHYVZ+8xOxV518APqgFPCTFVCDDTcypzU/zlNYRS0jcbKXjYBlmOlCAes5Za
j0uFyvWjEP8FqHYbRbRRlkHcjG4bN4BkvmTwn4sjMHnM4F0Z/8DT5LvhxB0WaEgU
H7b9hb3ZyFr+wbL7vReTbMkRR3wM5iCbWvVTPRpJmYZRITDNHOTEg/ISDRD5aNus
Us6yfu43m1sp8RK5PMfUhF70dOsVjnv3zlajYnGsnaL+VO0TVF1G0KcMkbNgSosh
T2ORfMaxaOuljoCaa1WJwKGC7G/hopCyz2Pv7yBp5bRPcOc+lyMg+MNQKPjOdjaH
tOu2QpzDq7kjWkPhPSt3zNBVLtcK7HiHkuODVAmN4w0DejJpy8daTZm82qRpgjyv
qBi8rKUDoV/e2Y7Yb+LabohBzv+Jm4teqKEBpWod8H6NHU140rImRwql9mHhNWAH
lsnDhN22s8YGQCQoRnwW5yNXj49MErUWyKsqMB9SJRUmJPMRod4GRpiQtl5sCqr5
aBxeeN/+UillS09xDaeYM0VYmG2ZJB4PvKRGbaN04Lfw8liFdcvWCrn3wwTSGMWT
64YPqUaBhr/PGIQlXU8nTU6xyFEr4jTMzxF1VniRc7chw9hoRt63B9L+jYCgBbmx
/EDlsuUEhHYo8SP+ay/YPquUvqMINdZvYkk0xWQKMSt0dGMzbZJB8ZifI/CEQUkC
CmHBjWnnHgTQMHdSBhpR00sRdUfdlqFQCJsRYWTrVLejZAMwjpU1gW3XAcGAM3Z/
k2O0Q961FP6HzHwOI9e8aE1aABx4Ez0k1gkhfX2khoA08miO/4eJWjHYXU7GVPp7
ak8Ebo6o9VwOOBXXYbjuMJVyNzYkDWpjZxV/ihnemI2UeepNR29hUs8clADWSH3W
bfQ4e5DfUhijgFTHNrTgk6VMtcO7mnnoeRpvt+A0hH3UldfmcqqdOEG3cKuejCUN
V7//x8ml00VF5zytEe5WreamyuShf2iH0TtfswXmPQtt3uj4gRgOFa+XlA0S17oB
vZZzfg5mN5u6ARJtyiix2tmzGjNM/aKl7+a3zCMUgn++2Tt8IsTQH+QpH8LnUnWR
y5aQBQaj++pVrHc+dP3eEfuU1isXztipb3bnkT48FlHPfKfqy+NYgw3IhIx4qVMr
Wzx2GGFTd8Hq6nssbSS/OYxvTU7lSx7wkU6S8OpSBEXHV2f6bzlm9mWbstO6pOvT
XNueablLTAcLW4bVHA8m8plOu/YWTjdUktY7Hj4dIVKtKjW2OHJ6SRh9QipZFTH7
6P4hDvTkAOXZB/+2W7YwGvyZVArxYPBwjcqjzaqcAREpkDLwFhWl5WxF4b2FNp60
1C0KebmjgNP9LH0sQWBl9Id6refYzlyebdVa2JCea6BN4ZYFfHE9OoylRULeYE3i
N9A6Dfnh/Nisb90XEW57Owbp7ZYLI5zBvTVfKzfvJOyHcN5Kse1guowtdIPnEyKW
yiUjEkCZ1rBW3mA9ESW8oL4gXZ+tFw3MA5A7KO8OwVSQO2IGurDT0UBthf7OfpIg
mwGm+bJGpEnwEnT+NJrl4PiBedNI0lfksPrM6cPo1TU4PFkalSz1444yL5ll3O9U
AKhGCOMwGiTh4En0AkX/PMwcaUXSrkxWOk4DyIHitdqJcxYFfhf5tVDnnueUuOXD
mP5Owf4QWFHogVBrpYHtsKELEycv33kNf9vhyOCsmAJEk0r8lNwSqSp+oFzI442n
GgSdQXJt+fk+pcYDiyLW2Dy6DHNNkPu2JGjPWA5cAjy58tFe+TQPDebJo2MqGPC2
K1H/uMIT+uhxsRONt0msdDJSoFlDeBHtKGXOOKIF5yVNZGzuWBfwYGH343snq6kH
Uj3/5tWZpyKVn8gbMBka8x3PYyB+KycutzNS/2OxamTEz5yrX9YqlwLdeRL9i2Hy
ic1oRwA/PBq2KeVgr9kmuiCTn2rAuroDuS1o590xkVsqbl30YtA7HeZD3EdIKZ3E
YdXmvUQhEOy6Nm2qlLnLjzC7sj5omcaUriBNuwZfSW6eZnah6u08gwFiyxkGUgQl
4HmpDWdqxY/NsuZGOBQLlVwLDwTFuANTe2BBko5vHpO6sb4QQh9NJLQ68oaIxWwT
kjxQwnauFtU2KrMDJ0/PZTQusTuIpa4OCsFk/hXcvbY6wbjKrOnwmwVM60xjdmgA
PeLaWlQVZ62+2dhvTiuyRVhbvZ93mzAqtFmtyqVPhkCddUC68we7GrXUbLS0jz4Q
6GvDzKLluIq4lKi5wIrX113WDWKbNWq+4nSXYkbegmsZHNRhls0mDcDIbX3UOpMR
1/Za13Fyijoau21XN2o4IFMFjybcvY1rbKIBB4IXQjB9S2MPWGiDz6xjthdOsoQH
CCx9w37RigchIWoq+el35p1x5Af371VxYG3ashEH0bhHfO8A83I0aLggs0rsyS/o
OOJpf5TEijllYSdFLHWjN9x/AjByXaEFViL54TYV8PnqKx7y9FhVVgxfktmCXeiV
1yZIazzIuHGbQqcyZqsITGo2QAWrrOvseGEU3ADPNBJFEEJ4ywzsKlTdWXDX69V3
3j/s0VQC2HHw33bhwA9gKr8hR70ZjgJb6nmeKrK68Cg2152R4cUZoFaSSVoQXbvT
4BY7ROUClM9eH7bvh/x7X5QrIEx7hz/G11dPoS0MvalPc4DoAKg5tTxN3SLfZ/7f
XUKOSzWYoCvihY1VbN07Km+5HV5gmE9zQ1CYRFAB3yw2Ryfek4SaibOUGUsnHEWN
bfDUTg5B9zmLBxlrzQMk/npdnvlfjaXV/XVV0EuVIOXjt9yyvSjSaqw2k+ZW0t+i
AC85Phv98RG5XHpp7NfN5mwJ5cYBt4G4ossry3Rzob78jlftrsqG9vtfgjv63zen
xcg7F2GdpbM6uMo2rgXhmvdJKIgljK6iRDYDMjaV9D+m1HRSwlQg7USosYAfirZI
+6c4RPiZGy+wlSl/ZVG+2VI18o8oK6DT2DeOASgLFaX+OkO+1E+Zgx/3OdtBrPax
vagtLn2dPtB3efQUkz5riq8S4h/f1xeqGJ8XckAMlpWNs6j/hnqHrQ78kTNT20IT
AfB/pmMVLUyVu5a6Fjz2R9rb13edVL77zOYvwW6Kr8p6MZaIoHfqktCbhX/HkO2h
qFC9XBIl20cPYqahCy2giHrV4zA8PFgb4+QOZKkLrYPgLhhuFIGpTqC7TS2PMAHe
2kpsujOAWqjmcNI+nm7PN55I8rlM4cxuNFVsF7PFDwKzePRucSJc0eT3Ep+KCHw/
hRZGlx1apOuvfdvBS9AzCQ8WwlQKqXsaANPzrKzAdZTCQqXjGWyFjWq+gaAka9ZG
ysmcDs1+oTTSxcMbPQE5cGXS5orYjGr7+s09DcPzecrWOVlux727CTnfHRuilxxk
GGF7lkFBZND2gfiPueYggq+TpNe06k1Vm2VGej2xWATnJOnZrOX222wpoT0Doq+J
qQ6yT/PFMcoPFSZvXdBcmCBaTSvtt72ct4CPfkxWICFF+gvE/GwynuPs2oXR//cu
32CcPgEHjmjZYXUyEknNprC+01Zy7ervtdNYnCXEDZKYE9mPb/y6lfYsLs20gA5x
wI8/3nnyjcrCe8rQnFM3PwAFov0QEmWibUeG9q00cleecwWjnAW15uQB67VreorB
tlPRX1jbMTRYo93vlo4WbEOoMwo5w/stXMc04/yQyNZCL6Lqdyf4vCRZTBCN6DVy
nkDXbQUPeF3TIylPHzK49UnvEx3cx9lnHcswgbi/D0pRCVbhiasTT30h7CAFlqvp
kb0+AnuFifN5TUmo2rlwuJvVUMrx+uozUn3lvb7kYAgpSLbxDzyWzq5/Kc3vdZaI
fFGbP+8skHF+HVW/u4NDCArEIuivY1YBTQVMFLG6OlOICdOr5o0fk5QLBlO47mDW
rc5DMlEbaRUSDGa3XAKl7moBTTloJtpRB9+AoexftC8lkBYPDbv8fpPvAhImvU6q
TZcBVMwts8Zjo4JqoxHaDsfqJ0uxxqWXILihUqIDnEZ4795k/6yNFm7thRwEQ2HJ
yYIvNeTo2K+1wj2/eNOFd93AIDYHrlaIDZOXF1eNkID2D4MARcU3EQcB3CbJIx1L
aJLjn4y7X9M30ZetoYok2QFZC83dEHePG27NdeEqG9Izg1jPOqzH0MDTv2NWXhz1
BMIiWacbuF74jYn6CD1t4ul8nXZDZIXIU/m0AWsAdP8uOWSD9NtmxxZErB4DeF4v
eSM8sGdIZ+aHNS5zOEe2Mzwk3j58JSHXcTPIfIdzfctujxHXZoeQShxQTIuHp9xA
0Lqo8cT5LMVCYRzX3i/1kRD7jPzexumGsRCb+ZifLmyKNwMCemB3MpAeLS/qoilt
0x02Kd8MHivfySTnAN5GlGQyqlJdP5wYJEL8w6j1pXwoS5cZzNmcPO0GX6GP3EZ0
f1ZIh+dv0H53TZ70fb0SusI4GZn/0SV+i4sslKlH1RD+5zR0fYwBmwKKIWpPbRk2
EXBP76LQH+MNhyQOzGoAdc8uWXRjTMUQTNqh011SvTPUCaJ/TY5B4DK1tF82EGRM
IAdhQ4n2jSYxi+v1mFQWX1q3VlI7krp0hIvAN/VjZOIEYvBdxhejyc/Di+sQYOGF
M42eClRavVPf+WPmO+ufNaBh5bn8eNdQudY5HP/nsToh2ETwrEZ4/dTRcbpAdi5Y
92M1MjNHImeZqhWwcT16kJQJr7NJq8ZXWvaPhZw1xRjoDKBl8Tx5/qj717YnPRXM
9JN7bO2DlMtaPdEJfo1m8Veo9edzoM11hieJdjVIKrY3j1Yje57jPzmP504ZVuSN
L1sGN4jQJgX26R5WEEkBz5m2sd5/bqHAgK1DQg67HGFwj38zrc3r4owI1Xhv69uN
cLOkKyjKgsfqrQkelSCv/UwIFeIv1csnj0ANYkXWChv25E3TiaVRbMoZ7IlHCa5/
jeX6G92f20gsO1fCBSAsvQ4CefLjADBADNKobscAKQ8U9NpYejp/Jm/x4H5YSWVz
OASzM6DIuKmv2PiiilaONhkVsjld40rbbaPaFT4mMXpe2qw0IUdgck1UNGJ7MCJv
2tTpRmrp2L8/l1TMg6hgcoLrU4CZ66vDi0xVMppWIBR5iUyMwkVLrhNJ+1/ZQf1C
/QT9mxcMKIedfwcODOHBbyXScNSdN0e1/BP9Uo5eijGjDRPFHPi/WqQfDF0OWF/4
WTFcN0RfEQtnhXb9w1h/ZdOXe+wFpQHK7kmrp09v/rINM8k2Sg7uYkttaTYx57h8
otOBJ3YAakF6WZHj35jiMHv9C/UFbvk9jqtpCXu5lPx1/vIPfxYuzFjGuXrefLuD
BTkU3FDNn7nfSf8PQbXgXWDmJXKvSo1I3m7G28HPM9u5csTvLhMk+xvEoqMVPg74
tyVQ7FfBTUpy6Dx81uWXgthmPvYCgQzkk11AlzxXjrtFtoHnZsNGyUrxeKv/Tm9S
1v1fDIBqw2OlLJ+embE2VgXimWU9njaNgkqhMzrqEO6dmcSeqm4itt9swHbZa+ap
lr99SyDui9+wSPHmpK4aWufAAp4kifO3Wz3O8GvJdhG4ufl1w+qZkYraEQNu/TYo
V4a9lurcqKqImshgmlEAJARihJStI/hsQ/ykbjCEYJEZfI+Vd9lw2CSYErUG+urk
9G/NGVL2TDwWXQN1A2ErbRWo50aG6gEa7d0CCayPmjoWYpTzda6vKQ/m9M5983qx
aBz1wvbP0fp6mJMFf0w0Gxf+8xanVALIsdOtu0jDF9mEyhoHvMcKJAzLhnZs7RB3
TYUrIZB638SJ6hHsrjva4hQBsErGrd7yE65Dl9uKfDXIEQFG+SlOvCBn9pBNZs/z
plMZAnN4c67sEyhDjLsK6gET4vNv4WYQHUfqbFBv2Dpo1tygzty3vRGGl2N/o6p8
XI7Wu0bZwRc+e3bEnkmHwO3VMkn/T7/hzAjjhy89lLX5e0nftOKZzE3Gv2Ha7spf
GnJzo9M+QifhFYwwEg1XaQVE4c6HB9X5BVdcsR5vuD25lW5SH2eW7IpERrztSgKD
VQgaYWSJXpLf6NlA7k4rZZNneUQF4RsB/wI6sa05+CwIYFaQ7Wj4cWoWd37ScRVY
BJHOQb2nqMJNcnSgaDxZh5KRluo+Om2bX1E+5gou270F1bYv1vGRrxlVty/S3Jfy
m6L1oot6gkMN6JqwI7+Rx6I39leACu28L+Ed+YKfFcRbunLw0LR1gbZIRAfWIyG8
ivwjx3t3L58BQsfDCOL6wE8GtufOKVt3wwTk7Nt6/bC3EiU9roh4421fqzy459kG
Y06LrysJkxSFDvlQ9zm4tR/NYNEybaj+yyJYaPNjrt2yevHRuDSxI0Op444lrQq8
xeiLpsi2soMpDGZRph1Wz9Ox4ZDQ8GwbF0tC4MxXH9Icxffar2UBCAygw7tjpXYq
atCmWP3dgaUCUU06VZ70RL/aaHIncHJzslvWcosMcY5yOfMjsb6/altkeSVmYGLe
FdQQg9YwfnHBOwnF9hHwmcEtsxj6QvZrzWwM1wENj6Aqnr/fcNx0KMaXzarGGZzM
xpBQZ1znDkREq+OUpscHix1DM/oAjTKz2jnx9vKLyA9v1tlnLEFZZGaePyNdbzMu
FbF/TWbnc6sb9XqLkrZzWKtSRSzph4/d9U9EgkW74Vn8I9LqDBrYXVLrEdIBhli8
NOfFR8W9mKpCY+avKdqM0WaY1WhWZ+pzgth3nbLK+sM+BDmuz23fQK6SFXAIwZUG
V+Lc/pV7Oi3gu0ByTMbyH1nU9+xYTO4Ceit9nu6cmVzuxwWF9R5VChDr0RD5Dx8F
4GNmUS3pVFpt+TQiqpagB1E2VEHliOrCQ3pGHeAU/YaW8nYXS7SRFfRUSayzbjWl
D+e/m/tZCsrJCT9Wg024dgevpHASC4uWYjfAvlTiy0IpEx1zjaFt6HaLO615Gszz
l92dte0MG3sdk2Ja+g45T3GFPXzP8u9wzva7WmY3DBg/KZRgLwQQEQ5xtbynDv0s
HHXVLHNzNkGY/6rFPKBzB5sIkENRZZpNHF/yawQMd4nkwGu8op5UbNPKWcJVP1wB
9hEMdGL4fgDdzcS24eG6Y4NKPX/3i2KE8p/d2rUycUSQElfC+b/AVHPnvylR1VP/
EFe4hoFwvjkteipjAmgckBIUjVFzMshQ/7lX7spIb8XEEyitr+hCHq1Cc6UWben6
Avc778n3OdN1yFMPtkXXCTCthC0wEExfDTci4iIuvLZJglVlmzpuuLsdhrbxCpT9
71DNHPcHRYDiMLQMnAXDP8QVa1Ru/MeuxEogT2EGuvykUYnHuLh344Db77xFhaUh
qxU5/q/KkUiowoYyyFO+CKVteZ0miYS8dSYac4PPiRHCzLub9A+5z8hxk4n1CJDx
9gNXQ3N6ym9Q82fWjCBt1O5AkuWp7fZ3hSAfoBQP7AuQJT5i4JA4cQ+2sRSNT2oN
YYaKzOTJW6cv1Td8CR9ldunuR9FJNOQvnt2ooblilHAFBcpGxNqzB3UUwoFcBuCG
mPIVad7RHYaI+FU/IVrMQsTWynQwVM8iNywMMgT+0Hu82uhgT+tIBq03glN5GDHX
wCqMn/HBQHjRT98ZWlrNSherkYESgQLxLw6HmSiWYqILrZC0e2dU8ra3SpUfnxS8
1lzWESf9I4FkLWxKYJW9TpJEygyuSeAocwjrzEjMXg0jdVJC7weePsneVFvGnzIR
IhEtDC+xwCzPSKk3P30iEJIQ0lLoCbm53LLGO/LcyabPHlUPE5Bqg3ubP2JrXhY0
m3PylMjuIB/hLUudgr9z58N5YZM8mH2JrpgnmLSsbNdEqygjd+Ondbk6TH6M+IJs
rjCEr7irQ175Zphx/2rrZPVmjVb/sIB965C8Swn/q2BJCl3iqmJqSNYjGc4V7MmO
mQVI+ijQ1WQ80sJdVC+JdPo3mQGGPjalLwzACReuKtU4IlaEEaaYCDCTDmobnb+B
agwbJbhOd8Um745v1EMLyjo5DrtrwIrYYVOB5RYiyS2J89FjEzLVd42IGb3bw9//
EI3NfTz6fpMjf0Mz55+hdTmgaHXhZya+DaMnmugLQiNd8JBuMn6hmV5xSS5MMJ5o
1EfHF5bEb90RmMZG0p8nsqv+XiYt3d0uqN3Iw3r+CqtGCQ38ywHRAoU9nf47ecbF
IOsMt9sntXbtOFG9XP2xGZmQ6hWN2gEyPX2G9WRx64VI4xygJceWkOVvpw4TEiwP
aNPnMCkkQDwGYMPWekTOfUxx4VrHZZvKQmCqbXzHQBVCYkkVMb6n9OoVHhrEWIrY
oGaT1j7JKam49OS3lwzWeGFytc8ds1nc1M4MmQ+KkPzaNz/rcmM1kyr7rAhlB3mp
8WjaMrjM/RJyF22kTZBnmzz8DLuRdHCcCcykgUhOj8h5lAnZvZ+ImY1iJaT9oXrj
OhV642rPi9IEYxPJQY6uatEmbF/oqF1BY+gb009KdkHKZrPKS31jfvqNuVojtXat
4xRae2cS1oBD7+CheW6wKf/UuSoAYJ7vBrQAXffF3IVYlgmLx2cE2G9kHIVxF4/7
wyi2P08Nh7A9Wa0BWMGBBVaNq3lDic176I+IbZc6G4Z3uPDJpEBPSbrNSfvctnxA
7gJ8fDZa0ioOC/VWsA3YJNkYOpFGs3P1FGiF9X+524alxgx8M1hFqSw4Qf7gd89A
EdCzVF4zHluX1SYbeg2YCT9EpcE4VGpNzhrH64sm8BqasLeOsmEYRUxSWVHQgRS8
RDrxFYngu8BrJfxLYQOwLDDtpIKervJQK5myCiX3YnUPnnQJ83nNhol0YB+skl77
90+Jpgd/cdxjT9upEbpPOzfVHdyzjmnNdwkT5ydtanDXj9Xl3zs9lNVGJbkXRBHh
NtqWQHH8YC08YJGFulnsTc/49R9I95KBWTucPRodT49zpn1h3SQ3iGXXeoQ7BigN
ZYKq1cGcQnRRZ+WldLjFfW+LRHnZlMXnAOQrJO+j8q+Q+zQoKIOEARsV3vRQzoQN
5lXbFzc4Wl2cep9I97DV2JoRT2/7Z0od2bUj44ktnyiBxlfLUYfcNJ7SZKItdLrk
D4JGyj1h87AZEiOKcr18roHMBq5NM28OeQBDD7zTROe60aV5FLOfevLx8VK44JQw
MZcEurpIAHbFLoQct/ZDg9aGypWyYHjxWpzugwyE+cs9i/D23F43nboHTPwMP3u8
B8dfxm+JTZbnDwwmgUubEzXl/mQ3Bc1YJOXlFih9tLjKXHl0YjajXZq3ByPycvtk
nvmfkB+apuksbcv/G1EgN0k1fN2bDp3npDmj3VXZyaq+7klEqnuKUrGwHxfJPry9
ctXOMQ6vw39B1y1R+ImEjUEkOiv9na31R4zWyHkkjydoOVzx3JIkfH+gRNbexkyw
H8WXapnLyLee22Z/MRfpqbnm5akyC3mMSv1Af/kK6cWHl0h6eBBzDHxn4tXVjpNo
bnEmv5MnetLB22mT2/7COvif7rBGb7SBZSSBvo+zvKHcxe0b/bS/Z7gT3ZmTJY59
kSTb+PXE/gvH0pD0x6dh1775uX0qie/zDlUkZyT+LZYwPj8Du9MKwrI6HuxpNZjI
FRGwnxfj62p03DjqEXkECNSuEySwTeHnhps5nBLIq8dCzVqxIM5Zk6bErqK4lxtN
u4laM8udIGi7J/FvEAJQ5fDfGijlbyG6cuHDgpmtaR1r+ThXdf83zkI6k5RC4GNM
J045I9/oOutjf4lNr2J+ljkKwLGRtyXmhY1CzdBC00p9PB6clhKJxPVHkfnvozTD
7z7irTz4bnFWbmQ9kQFmIVUr+7FRzAZPgBTpIBs3xeiLzVGdYoS0fpenQ8hucJIe
bwRFbtMmSF/g3bnxFpmft1CEG/PXkWb6MV3kIU9LIOVwE9h/VspicBLtPoQFluFi
+e/yfrqLO46OIHDU4k8eimuti+GaIBPpEvIsh/Wj+EDT5Kaci3sngvDGJapFDTSN
AvSaUdgdUHf+lGegax07xjwjMo0PPwV6EC755j8TEdjmH+PubrHf/wEOTYS30TiS
emZiNiINoSfTLKmplHTlcYLNgeKrWQcTKznR01lpgvk31oIagYpi4rzQGfeIwmpC
ujUDlfzgl4Shs+7RrC2+hleU+LJpP9Y77IEQKpbXUHqCgy5j+2d3FLxt894deC5W
b1Dgzp4Ik/KJq0BXkwPXsPNVuDNDXA6PX7BZsb9E6/hDka2MabO/t5117oyNLhAp
gAFrgKvLTK6nlL298Oj/JIRdCM0FH/ot6b+Cp0nYpeiO+eCpHEWHYyLFaKRkzYhe
Id+lJfj+4vWlPdnkQeXi6R2rBE5+5Dkf3/wDKxTSy9K9uFyE0zSNnw7V0HksXxaj
kjkf4hLZxNWUtWwZEJ7uNOkRUe0AtsZpGUJDJK6u1gYp2i4P2QG7c4YHFCBt6cza
N/mq3yzmNszzm1Zf7nqShZLyJ+r5N/VyURvfiKgfLXWmr0rDDWlDiVeu7as6oD3o
rvPuiZODDbVog6UAGyC2NXojmNYKDXzIXPR2KJO7Av9ODG9d+tC1HgIm0STzK54J
WAs3e8B2hC7KNnXIlD0a2N9FhPNDOC2G25qa5gad8wLu0Y33LNbROlbnQukImV1v
hZ2N12pCd3jBPPBfs+mp35x5bmCEgWRHEI8m196HLYDHPMCpVh9eOxNCnDEk63T5
/EFDz0DbJOyMpdh0u2fVSTLi3rOD1yAEIY1b0+uwTdBc/xghR7RcuJ/6piU1bddp
NAt48I89KgC2NLQwIJq0/iSJdih+mAFG4pm5kEfZgwXeXJxJJqUbOxksCeS+As6R
qBfB1qmDlYJPjV5b/mxoF2jrxMemyYv26VvVUt3LEqLpRtklKRxeT47cKV9p6pJV
oBYxhzu8RAMa60mFIVtmBTCAybimRu964/3STPKaNRCjvSae+EtFDdVXR0ywKUEx
iLkg7+JWbnGmUSbaAKO26GF5yyEIyzkS4fhhii98BmW91bnDmngheDENRsnjn2Am
m7MGZqxPAuAGMoaKhjTSA1bW5bUbuO/UD0XQaLfk8vQriUMlkuC4bIkVWIOznBcG
OFfSUU9TyDKUmv5OUaA6JdAiGSx61Y7XdSbqyR0VWoHBNolNWS0YI/WLSWkfslbh
YD6iW/0hlJLIGj5uY5yCDmaNmRKd/PKJZdoOrgFz8l81msYI+otNn7Al/3CXQIio
lCEH8/whHCHGxvISy+Ph8w/j1sCK+v3+gIhnEdQiHEO66zNGH20IT6tNB6EJmjci
cY4B4T8epL5ampqDEqY/I+3YaqrWzHB5C0zp6/AEy5QusBB26dxJbmbzfTJlomA1
L8LtIxox6ym2PuilpataBMqpnflzsAGOyApBYPDRHu150J7LrpAXpb4+TdxAXCMp
LaQ8XC4elSa9vyHrMUjfs4kd0+Az9eeA9olQejZq+HCtsDV6/hckqbmKvHSsFr0N
6vUohZQj52asmxcNsR1CAhPjJTUSSKACJ6uEcfvf+z7gMxS36aXfj3m4/0uKe4zJ
2aFNiS31ZHNam+36iuTfVFOGkRveFUg1zMIp7dlA8TGtogbNVF6IJDJvhncaKAHu
eLAxVoOcGfR5a1g0fS9bwwdlLqQSvQ3k1NswrLFBgziW/RyCgir3s8zFznz27IyK
gy7xXnTpsr5LJSFtCg/lY706R7wnITW2+g2NegkGC9p8F2zpd0jVnwmrvwgLmtAE
5RlxBROQQKxQuwdrYXbUTy9cD/Q8ZoO0vOhIDOSFkw5t9v0rLokcrzXGy9pIHmp7
6frroRo0llZYJPIyObXL3OpRkHoHSKx7gkhXQSIzVxpYmwY8IwgKFPyopvVft2ml
iglehZmtHQDpUxCPbd9TYaVqnLFj4FzN9mH42Wa8hNDu2iL3kSGzlJ6cEXJFsftT
/sNw1uALnRJ2kJV7sy5KaVZPN6GUnZe78Rgeljdy6JtRHw2FrXXT9nn0NXlpR3+l
OY0ZkL1+5NhkXLDOmIwMvB2WSaxyA4CB5ZELh+oWEY1RzspGn759gA4CtiZGeJfe
SvRXIrSrumY0QIgYHQZ+4Lz8Xo9n2ZeWnwq59XrmSXNHUphY0f8T1C53BKyvv4q2
OuoVsJpoM4e417SvW3/yI/MxQ8f48u8cjAlY/ywd5b/+b4FJKRhC2F5CLe/YlEC3
nPCWhb9b6bgYvwQcXmr04phVyZUW0kYp3S4DklTKr+QHzoadofNGPGNoz6Tt3kBw
vrPFvSu/hnC12hozbMf5eYNOD7iXp9vbWcMTVxSH8uDN0dnsIsVeTyHB3HWKjGmG
6NEMaXtckItt48q7Cka9Zh+P3AGDtHFxHEAVIxQllplk9VU1EqERR75CRNm8yyrR
x6UzsGPK9XUsL9F/irYpgboRxNW3i2RIJLewMciUkxlXiUuh2xHkR2rvFi/NE+ou
uNMJ7LI/53Gktf7sbuQ0qHwXjn+0tjfeyzjXsOTmdDjWTgFyxFNsWuPgZWEVJXYh
Saj8ZefsRRz50CjiIPL2EBHbRAPq4PCDtAxJ4XH/i9au6D9nsVJilllFZGcu8g9C
u7QFg3auUGRFrQOPSISvNAyGr/Z/CtFU8GCqDrEdwV+cjUxCuNSvPZU0wVyGtGOQ
TCogahSreFmKMvz+wkckI0D+LMjxv0mdG7bUunZWfyPilXqtoV/Y8Ow2PkTfB97a
wD3WphPK6v6F956j/FdCAhYSRW96p0hnBzc8FpyOqi94zj/MiYUbhnYdf6sdvdgJ
49IeNyC/B2wBjmhqOSO7zWaJqJhSJK+UuFMmrOuLOAOhhIs/TLrWnFsgQ8Nl39HL
vhEfCYFSLiMHDLmbwFZeTS+muX3UmbKZi7+r+BKjzc6kPYSBkzlYmBbb/AjPP55D
gYsOLgIvzheZlJtrIC1iR7zfCYbeygL2slhgMDif77IrRuY739oab7soHLzDPz5f
YmZhbi6axYgS04JMPr/w9wbgK08FiGlpFBq72My/VQMfilTIm5GDiz8aoPV87Y9O
ki2D8/zQfWvrVMP6jJO8SKZ1TgdL0pqzSudPCtPDwQnGFrkRkN8xpnb5IcBtDF7j
MhebV0UL3pVI/nLyyM7UBFgV69pbN7EQHmWD8+LpBlo7gBKb6m1DigFyb1D4odS4
k0y2iHwGe+v9KbAv/IMP2DI1uDAI9GScXRCEEvtJCooSd5J/NqiLx3MaRymY2qbx
ov3GE07wls62SnzbnWwKTfGPKm2E5+qBnUAbFv45bxmciKnOz9EmZnamO7q3Wa8Z
j1V7bvJzcUNGdAT3mjUp/uADNd9hpqpkKJf+dP2bdIw0p9UCQ5rCgS0LqiOEkzB2
He0EQDFHGnNSF/2cSTPBEdPzOcObDAXfzyuavm9rNbW0uJ7ASN6d8YLgijnhdw9R
e1q1naWDckGYm3gEfuFpIVrz2761c8qknp+jPPgLfrJcc6sT7efwdHcfvH0DAc9B
7a60cHe3nmZ/XNYaYtqEc9QOXYKAY91LIE+GQQ9q5zRMAvIJ0i5qDgqFvZ5EnlRX
DZfcrXUKt/xcHJiUKyeZ8LTtUoGr18TTB70Hilfy5nYqq4YwJKJFVNGK2URGw3jX
QLQRfmnO2t1EkEyD2NmBt98D7UyNM0V0imIRRqdxMncNmjBB9SqyVjyi0+8HYtWt
SBC8cS/T1GRgXZnrOG3zybUOBeGlhw96carPRE5r4y80QWVvrFNU+IVynDjpTWG3
gtpb5TS+o6i6BOmEVakCaVBjzSsCO1LuViLTYrUqk1l+KGrbz0BkucKfq1soueQw
yQG7P+zdexEqpoGnem0mz95N+L3TitHUmGlzNzTGX3aQp1t1FDPTS/qcMm86C7Ce
bTtjcTYdkY9WHwRY2VYAtvsPqoxSnWEssWFcOuTmhoyb3siCz9fWz6O/AqWKz09d
bAILvLgx2tjc4DCLqJr1MHI7X+ut4JKo4A2ImbO2oTxCBX/8H2lVyuWvjmrduM33
uyH4BHuZK8yYzE0RVaLAh5hGSba4wYv1k7hoTpx0iS2V9j6w+jgZmNMvTf61s4+H
KX6cK7QTG2NkT3K0vu0uK7zObyVzlbvRaYYNmg8BIYGW4AHrEnPZTAcBxwoqbI8U
PFcOV4SyzqOEpUIwV/OwJ5YV11q0zrmKJht1cukbx+QdY9a5StfGWor+LPr+wJJP
29JdysNuYgQ1UAnZQq/dni3SkO6i/gIognyHYIc9rQe4MUC5USYCu/z6T5CNn8Ef
g57b1BApXFezdrnj57urVSHl6UIsB0uvSfeVAG8BQj2YdQXUS0BztJYLlJYFqsOQ
UoGDCnEOARnU/yzMWNP8ghtkW5CtYo8lKFC8qWSqZXNyCz1NsNvj6bCHyDRoUH3d
t0Wec94Elc+JXYztLL1l378m2USIBA4BVuyuaX3E8HbqgP3zIHZsaCWNSqphV4x1
soQGr3Wb55PIJWdvESb3BUlmXMVNsG1UgeROYjTh23sC1kcydDGCsiCJTr/N1+TT
iTxaOFCnP+JG4BhsTUnpqjKHsGvGqW9DBeu4rdv1bVcY3tOnVXDFwVTD7/UK2USi
SImWWHeEt2NvTWtSbxl3CY9mqittRGB7gTYh01DWGKUer9dOqkV+xeKYpcK0fl9M
kUz8wey54FPWhK2+sxiMIsiCAbNdlWohEnZbf3BYSpGW+jkJib2hCVD0dQnbQtfZ
GynYEmTkrNzvH7anlA9KX/e8kvqH7e1WpC4gO9D6DQS9J1XBzXCTVsT2FcXd4/3l
zTReG856ySMlQeOHVILuH38ZGXYpZW2gCypdBxZMi0YEs6jhe0ZNXJtZafFP8tnJ
/26F56FHbhSx0a5kXIsWA31gTQeOsTPqWCBglY+4YRDXtp0DgN+m8KG92W3UayJV
ZHt4/gbwyjvDb+10eH5Znz2dfOd5RvYPARbFiCxMy7Bi8yoLrJrZdxvpiX/Bi66o
8a/yYcfz2LVJFba1+Cv6qEYsDgc0PG1IRZsMt40LuIAmf0423wuSGEQ4thY6qCtr
1AgFusO8D5EvZPH1+LQE4WXSWXp3QHAOBMHzu6tD1/1oz7m13svWrjMczNLAlB9O
4rAj3bRYvyiArup79L2soSaH6SvR4U0SCQ5v4wjcz+Ak/BMTmXFGkYkN12yMxlsU
GDJjmajP7pEv3T52hHKBPvRCVYv7u7deexFKzCPUMwSfUC2kr8fyaBkHx0XoweRm
cLOqU+5G+b8qm6rG70GiJt2M8dK9pjZqBfV3qi1KPNcbsxzqt4aq9GMkh5WJhJMo
oD/IRtlR6m881+uMd4zJFYzlvG3Z/F1x2/eneWaRDqW1S6ArgmtHEwoEmhA6rO22
4HzLYhPiZdp4Vl2ISP8gtJH+VjPME/ZXhip+uhBkaQ35OsnzGnfCOX/wkfJ7jUYi
JnjsnmstPphMOoUut2/X9v6CBWgoS/w44NivDqplrXnhg2b0yVUThgZ7i6CdZHfl
E+F0G1acbhJT0LDc+YkDrD/Auyb42HK5GG3eV4KkgpX54n8I92ezOy7gbpshg5Fs
OBWyfg/PlG+DmqChi1DcokkNzWL/+Z1m6Nr+TY71A6MgNs7MWZ2YvZnfaQau9Kbg
eD/+5ukvJht/IhX5Af+Emj97PCg41WhPvdop8t50urgVScEwX/exny6GH4HafzZV
aDuSGfUTm+qtgIg6Otfhk+zJRuPEpqGzEESgnmvsHeP5Q3G280SKPYte3AEoYJee
A5YwArqTcpl4BBF+vdGoQKlIhVqUsJDF+nRtfZN0++YaXKCN/2zwJSHh8cluDIco
o/QOZz878gPjLMr6ZompEXWuzRzZqFLAd+rApqN+qGXq4EzAz/fkhwaLnPdXhrwV
7NCKki0m2VuGB1AdUOG+hyB3sCZiLrAutJH3rbxOxqidCYy3bZQuS+jzObH27irt
/tJRHnRjOsjmLJa1v6mquBnE4+J7dOy/N9Om8RjK35a22CFDtFDqIGnnqX5/vgUP
8/zXh6mmr0T//Tbdlk6/PIDnW6AvQlQU8dxS38pqQd41zCa4HDJtlgFPb1wGhR13
al9z22LkbJBfbl7gTYaTB6A1HEUn/cYPeoqo1qRHk028YqiindVbjqnYdPsr8Y85
svw9PHhaH1Prrm5o0/QvoyNbVQa2g0/GQNRqVEk9lr6KHljIldYIoKlAXiNeavcc
nREoEpwP3369+W0OSu6oZZNXiDLuKPvArXm4Aum+ZjHBhL+6cLqnA0ta749x8Fiy
qpb2Mzm1NQ5axlbXVGb5notLaTYLKObfmEGfxFoHliUjd7Tf+BASKcVEJ79ouUv9
32G2vnF8/SSUYJvD2D4Ob2v412wHD+KcjkeGSTtEH3CBt3EKvPqXy76kWRRkyD44
8gIms98mKW5L/o516wq47jC2H8mrQu5iWAdnPQj7Bl2gYhlHZfEb2pWa5IM5lf8q
W4FUlAYllpGYNS8rdwHlas17En/quslAYFLTwek43TTzgvPMG9B3WxIG18ByZ15/
e6yB3m/ZPXEovJwCqa2BO/0uPjCoN+ecHAnzYCQdAzmZiMDQqoyRAKpzXnh+SXqr
GF3wn6Stp+S014MKu9FqJz6UQ2RZa+CV4+vLuvS2qanDzbogRN6BGy0yf39OX5bA
69VGyNiEunq3n4Dd3ps4U3U6FNTii5ZFQhtR+kPjBIsxQGTK1wRq83h++3F6RzTi
R37sVJqYaN86mB+ANmAu/5yKpWPT/XpUBRY1N6mGsKhhMyADbKpqSbCAOEBC0ZLF
4bXfZsvQkyyWv6LuVLTe2p2YLasghZVukfCt7KYnXLSTRORC20afgoDuCnfwneZA
qyBOlwOK9pOHxfoDV7WPaG4OYe34/Po7dBGeM2n6YSyciaiDqNzYZ9aj2XAfHKxp
aQJjOx+aQy+yRsMAuiUL9vd5CP2f8PVVqNADhV69ZX1TtcVBnQ75Ds7tszt6usWJ
z5Rh5RxYYBV4zGVOJVCdDd+pPSlSj8vHmEO3cdpj0MNAuJgXeRXIyZbN9MnUPBiq
`protect END_PROTECTED
