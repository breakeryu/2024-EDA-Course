`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7IQyo7VZkRPCwIufhAgrVzDF2KdJugIIcAyNKvpVmPOK/u0xVA2JBUyD00T+J0F
FDRjaa7uvkEcZ7SS4VjKi71X+bg1RtsNinZDfLuNhHadVBXxx9hseWlxLPMClkIZ
WCXH14O59xwIm3HQTOXqUmct1LGEy0J4shXeB5JAZaibtkiILXkFJ7VG1fQ+nDqj
W9kP1lW7IAyBhfZDlzSFZhBS1DaTztSIPUHJ/Qj0PffQgJqFzx8c4MiB+fPjlqr2
ILYoXT8bdP1MO7x5maxfQaEtrq6WmAVWoqgmkVQ+6QnPysq/HVlYv8spifBF1dAG
wmKXKFUCJcY3tE67wKDVQdrFXMLc40g9X5XRLngc9AjIuAPfLQhm9uPxNhnpdsCG
zptM59d32KSdccE0vBTaynrZiFDu6Rk0w8zPkJK+tWbGJI6YtM5ErAv54IFylLvZ
peDx5+GxcAqWB35U7SQGX6j5ZxDVN7aw/P/1J5kowYTA806qa1PV07kETm6gcqDt
ge2ZmlLbw+1l1HCKYdpJOP3PWfGJN71OFK1zIfcSXKKwf0CsevP0cot3Gm1l8ZUh
ViEnOK3nAjvJdsoBN0RgzYnt5nqWSElRcNxx6i/5B80nQxDQ0ffg6tJU3ed8wfaI
8XickLGn4odmsaY1K3Mp8EAupHB5DHI5wYsgVCD9/SumV3Ux2KAHGp6rCtrkci8+
tPLp1vsnRu3aG9Qn41A6Suv9mhqoLwafyN2Kjxi8GZFsNRJN3h/ddfFpzbPI0I0O
RYB+Jp71DG7Y5I67FRu2fCM6U2RbiPr5Q/aGLR000i5VeHDGWxWgkAPQ76qRMqRQ
+oFjwW2+ZDrqPUGTvwHCl4jegncjF/jNVxBC4oXnI/vBFgXV8Ss/hC2Gy/6OnIJw
YlTSFz0TBThQKSSiMjzcVXN1k7vpDarlV2FR8znxImECr+MOL/ictQbtPBHL/fYV
kiGckUCKrmxyQvTu95ee7s4uIdu9pHBjEDX81nUbt7tRT2Q0TbQ/XB597AATbWQP
0OY2/1RonjbM1IY6S5FrCC3OPw6HdJK/vvf+24BF1kjX5g3dBmszXGRROZ6Jfl0l
Oqh1+Jzagaul40c7DfIOASQvnWQULyjGIcSa9aIkdD3jyVwWVDnMkm85a6q/RKnx
J1TGyH9J4uanXNuwXapJGznSRWrzEbvdp85KplxCJ00DqxxRmTtgGrurXa7Fj6S3
QWoEiwbGzRu2fz5kEqx9YZYZC+CcB74YYElAtwh/xg33q0zcceWp8S4ShMxEGpL1
HiidgEQV/Gx9aFrw4k3hyoEVnpOTqUaGfAlnie4uYESEjewyQXwid58CWPsUCCyX
Uv92icsbC8Sn15XFBJjurXv2jz/+C8mD4DbT5LKQb+MqtWR+yC/nFIDRIOHveIdP
z7ZkmiEiC6h3mlCMFxTgXEK3mdY8m1jmXI6yyHVJ3tD/zC2RXEIoV9Q7HewAtqt1
UTfPxGz7z99tTbd/N8GH8zigIFB1/0WRIuiZU72gMiPdjeog/EhagUgnM635B8r+
FfzHJ9zUkFHWNTZaqqeVp2uPFUZ/c+5IPNEhovkaw2RSwV3J+YtXTwpOM6ei8BOi
DtIrE1VPW8KjXTEdfJKlBKGx15JBWjAzA0wqK0xhlNbAmGz4/YX4rdmctoAvzQvc
3i7DwfKkixBoaO4Qfq6gJBkP4PhO3U9oGQasNIHIv3OWhtVQN0SkXzoEfqL1bq22
KnX8Fn7tiI7aqP0KuBntUqgH0nVvHnZFSpj1QMKCSRamodhVvsRMy/UJ4xb8NEmJ
gGUSD2sdhEcszyrEUY5BEjsdA08TsEBj3wu9+Kn+oILeVQCu+Jj0pGL4poJtuSIZ
HJT/UVAfNf3hli6Wpg1XtOCv6Fwy8szBXTlmDv/Bc9apDzfnrupjSsK57rDj1X/n
1aZyPblMVLY4AP1EDKijQ+hbnop1eejEUuUlPVshBDT5zne1qGd/GYEPNfTW52wu
DFDsn89RG1quF6goUxi/n+SKSEwtOt7wLHKVkdtHivrR65rGfvbshOimKpFstqEh
yZXNqZqWc7r9dUdbAyMc6cPdSTu+C89bvIaMP/YdcZdQbAoIbbI0Z0SlGNTL3rs7
lk+jmxbKHDOZtn5+b5M+gzwrX2MO90VsAPHHm9hwhjNH74G8V7WH0+ldw7UEBVxp
TMajjPGdrTeEVimZCRyscStU5eq7WDprb19K51V/sFDwDkqKlEX7kmMdMIcXGXhT
lPzqyKYzS8W8HKALyrZ/LSy6uGDmPXz2ThjQaIK8LD4AK/Mk0YDVxDHjNSev90m+
O6YQnZryNeRuRLk7zq6OVpc0cQm3wByKwrmEY/m2bcKYU6vpa2xafZscNcQfeXbH
Ojo91nOkwW/aJWDuybFlCdxoJjbUfZ+Iw8nZHB33jtR263znf8IPofdVDx76LQZ1
lPbbVq5LSmQmgmZBVpPukyyU3XmrL1q+w3Vrkj95Zz/PIn0NPBKHwnKFU6ghTQTS
GOg+Aq45vloaBGu+M6npn2aaiFmlzL6PF67EJQg5o5D+slsVfLtC+dXFuuSDWRLn
EV1wRtlMPamaua7UIxZmPsA3kYfTlEvVfOt4n73vg3RYihjmODhs8zyk9w1hYgV8
ekaHjEt7YjRxbeqFOIEyKCwPVGIu1VhqDC7B5DnktiVcatnijfEkM1yeNb3Cdthg
n0TioQ8OMRteF4AL8odds8jsV2Y7pPXK6N/XaF7yrR5UgfSJ/6DgvACZqzpwXkhY
dLf/Mh3i11MblO3KeSZ1A8Zud1T1AkfZh8aHHgUKln5K00Ze/c7CVLpBdBZ5PE/D
YcDeuc6AEBq6p4adfC6IFBh6FTiNIeDatEdC4Eg+2vyLURDMD22cZ+SfIYMBbrFx
PNhLkPtdctshtLvJjuHaOrMATeyS5sL6zCfTffIINBNXS+vh/dabwscEfQ4GVEhe
qMXKhHVXi4WO0q9vJYnv5F++1DLKfWe2wCSq0bx6vEwLuZktN6mL8jyh4z+IZa86
7ytVRMhce1sfSbdTcnh6oH7ONZZxmIQ7CvT0AFQW9Fjtkbe4egw7DvRw1iA3chbG
MkXLDVbiBKTzF1vdnkx0bU7WaLnYbNwhksG9F/fzbRnZCElIC/Nn7t5orikOIYbs
Mnew5y5sj4xCRkWUQVt4GaxhfDB0wXsNFgoXJp9HbWlZpR4J181fKO5XVlhN7GUx
6bp3oCRYWgWGCVQVrZ0j2e6RD2DmTaDKrJRjHLTtTyHWeJf92JfARpX526RpIuOx
dj254K2wmx29uESMNwfxobkAlJV9omFWyy/JPM8wejzu+AaYaiuTeAwOaKikcIx2
LazVmnSrqoPr7FNOpS4xZ4sOTjYgBtww+O/oPGnOzUhKdAtZVHfkZ0ZVnb82S6VJ
ey76PXV/lXNLUnBZ/BDI3S5OlZmB1rwQzzoi1UIX2vUE2OQ0NTM1wZecWtFcIcAR
LM3tidtjOO7+Nh7Upa+7biGNCXx5EDFCnyrZqLM9J5aI3sKFb5dCvoLQMiZJUz3n
P6ceZUKA25ERHgyeKkNmy3OE3zMPvq/exI0/elbE7vEieF7QUQDmvJIgRt6HMIJJ
DsnllqPlmE/NcxGUl1zbUERpx3/5FOvqs74FW8KZAwyLpzbFK3wuDA5BwePAkdLt
tdIVPynXW3+kUDMPOv8Y3GkwbaLAmJ1s6J52GQXmzm31AfoU4AWmr+mWDGm0V1gA
n0Kab6IkrtGMxnc1940kpELilblNFPtzOTYqm4r0gn9hWeQOS7jH+gSE/UrTmhH0
xeqx+CfrOQij8MOZ/d/2239zP0PLEwL8OVdpPowjrJS5t2bCX0h/QdEZa1E92A91
wHjh7TlUpQ//+IJlgGtsdIBmkqxYIRQdpUBHbJIcxL7BpiklQ8ft6wx+LYl02CqX
8fIc9bKbbYHaQg1zJwYU5ELB/X2LyaRo19r3ymfZ3BfnMkgGHG7zaeizgCL0ixe4
VQADCSeuwsty8uc7h6L58+EU9D/f6SwUPiVL+Uu0LOfmIXeSJ6ptMmAoFd/C7ewY
Ac5/sVw6rn4Mi6s7t13EgaaHxcG2GshROCVj3wzaeIYqxWb7MsmdJSAsU6bO7uOL
4U4u5eITvW7bWsCL5AkAtkm6Jxg2Y0T+AHpKdenVk41VKrCKvRLogr+FRDp1JlB1
AU6QdVA1/7d1mwGPd1b527QUGGHQSfj1tZ8SXC1yxai0TjOGIZ4tx7u4PKFU1N2V
VKxPzS5En1uEYe5AsAgEmkxdIZ2Q7yHyWB9Qnt8NrC3u3b24THprFDUgDBcqX65m
kZdM2p6iCfVSJheXiUR8g7XFzXfpDJE3kCPfFKx9oa4jA6iYLaVMue3194Ejkb3u
2tkq/VLo7yFC+L+x+Qajd5Y/Wkw6iqKOaEotF/TopHSCsAWr/grM8IYidZJh8A4V
/ulKCPc6kV6M/3HIFKF1uexnP6BHjg8M0ZSdAH5nflShfnHKJ28/r7IJHgRPcT4T
ErOSJoJ49K4upS3DOxq98Vc8hpQBsB6nfhYIgy2nVTK6Vqj5L5+Gyiu06F13zkva
iS0jMtujJHel9ZcXfstmyFDXad85THV4jlqUtGZNCTrT1NXGC+bLBTUx2VP94yn2
ydThkSrHCdv5f9+F1RugrMPowME6Pvwp3pt+mn3co4fdKjn9ZrMrwhMJ1Tnesjw4
t1G5uE5R4yKS9TxwniNjBoo47NS2LxXBNMir6gPJ6zUX1JJBDuxmC7TW3CRDIv0L
NQXnBDSqBe5O3ObQj2kpv9UA6nr45NpIHc6PI5cWXIv6CbVpwhGTMp6n0dUQelp8
SkAJyQ/qbZUON+2+aBlchCBlpOSFRW9QHcLzrd9DXulNfKMj/MOGoG2ugBJqWvFv
+ZZ9VLLMQgusc4Jlj5AQErfJayXq6fx7Rjpkncb6zXW7cG+rwMJBVl5svqbKrH4m
71VTovzZJZB206zJKh9JPrev2qyyi8cyr/auAbkjMZ+1nkHR8fc3sRamTsw7xAuR
43dJhh2bf4NY1156lq5GzzfXUKzRcT346P6HxDRhZ6lJWDnlGGRG2IISKBHHf+tp
a3GAiEQ1FCcPjdKEB+DLznDPQq0cSVrOVnI6urmhC3e5vOPzZNL8fWcJIqMqQeER
JwAxHWZoOLNDFWlZZzfPxUpCAUxdPhFYqrNRzuFdLlptzgObk7MAvoWxM5+5NiUA
ZSXL+DOP/cIRbOTdvFpi21f0gAlbCS0BmkcO5TY2Pv/F2ZVg72CXbpXhA38gMIm9
yRApaLramXFcRXdHNjw/aA==
`protect END_PROTECTED
