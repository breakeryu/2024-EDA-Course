`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkGNqVH6QlCzgX5s5m9YTa0/qUGcekrNalmIKNH/IuuzpfTAUWVXfJpd+KJ1CeOh
RfVTbGNof8ytfruVTpV8SL/xZHuDeER7laGjA7y4l2kQfJPq++lLOrhXRjebCkdP
X7yqdC1QyrOcthykEl7fa9rxl32cBKXCY0XhXVMjQki5bJ4KdvgoQU8QshWnBAfT
8TfkCl43Rbrooj7b54tmpos6v9TvezrrVkVdoYLdBzHNV/bKwiKk/gdnwscSCHRF
iainHlz4MdIXnYUwlfVRDlDZQ4JlqPft4XIegQzz5o+HaiXGp3NKuNLby9t2sKoc
xhe73TymXt1rtpwM2y/HrSvlJT4qU6JSoz6B9bGGvNoxmSIsKqcIBSnO8LHjOl9I
XqvRjk/z5Ph2bARvZy2uzgf16CPlUhSyywaMZ0r5K0dPlO29wxdvxpY7WAjWoQoj
DpF6JoYImFcV6NjPx3m1EcKU1S8Vqi+1q1E3Q9lO4ytYDDszF/TyDfz9svGMqV41
pW88mrrEm+YZbMOuv05OXYkmX9B4RanAOzIP0dw4q4RXYFliNyETuexn45I3nGqq
t973IyMxPPFZRjlJMDZqPj/JvRH8Klul6AuRu960E9r7ACYeA790br8AllKC2MPD
5T7arfm9MlqxfbPsqJj/IK+YXSQ1LAyuQpR33IafkmJyStjer//laXKKApHI82ws
V5/lA0u3umKDpUGRV2SnKhweuflbqfIIyHhLlTeHLEZ9Y3zzVsxjQj/OhrmG3S7G
rpg6gln0ajMWKZOjaKEbQhGO28vCja+dKcAiEar6IoBLlcT/Ol1nYlzaHDIZkb5d
8V/GwLxLe4F5i1yTOBLrRPYFMowmdvRaYXeD18FOqBLK+7oGsLoAGJOBX2aiJkyo
UDefbgtKs2O7yBGaOPnf0rWzCWsX19e2MJmNEKDP4tT6/yGSyqQQjPu0M6DwRfzA
F9tAQVv8ijJtJxfz8z6TdH2gxVWK6sALpXsEAOMud1KHADMc8IANKoOmjtmA3Zsq
bjtFDK1+dQEww8u8f91+/vVEp6Id1L69UjwvJINU5EPP7rg9plroCVS48ABOWaWL
k1h10Vz5jtAgRInakbvcGkxE1yx8ocB5jczQuiP+i+Tn/ReJNTRJecv3fs0ibUBK
w7v7qTFEHtHXn+2tqnOYMzIlilP7D8GvIU4DcUU/oZ2nEuJW9rLVHaFhUfTN9+0K
sST4zg6+z3tm42CwGEKHfkL9hxEFhwj3UBh6qFSQCyOKoTsJfFWhzZnuAtOkUqdC
Ptu8FgP7yshQSblIfcIsU6ia99qEvjerBokkE3SjmUA3oA73txJq1CDv+VacfUPn
k0qN/tTMoCYV+Tox3R2iSUzYIP9yRmEBSsl7fg3uMz0VgSlnVZ4Oubsqd6+G15lA
nh3zzCRUq4fwmPbZMr7xXSlSEAZMGjh1Tks5dben5accObwBSGpedr/hltbaKJ56
SeKxKBBZzjc1F4xLtA0ze+45KttueohY+0J2ERco6bGxRGWJ4c0kUecKqS2eZaHK
WrYBzQBKMjpPOAzkXd31KSlasW9KRN0rdEt373u8hbaHFUfN/3L9z3SVsOtVnRdB
C17mBvZk1Vb9jdaUvEzZL5pZYv/EfYm35GjhPR/QcQIkPpgdtDqebwjSKmhUKmgu
dTBfLgxgP1h0i1ATh8i+LvFafaAnto2lH7oqC9ApoS19I+r0qUYuDmIsDu9hiwfX
75SZqB3LaaP/PKwlYl3bdXmLpSQ7upKMZdUz1fq5oYBFutzQysXA4Wjaa2w2DuK5
ilkeYBhtj6bVFAcciWrd4U0Y8qFV0IiZpXH5VwdUaByFAeiEz2nnZwn50NnO2FDe
CBpzYo0Ew8wQoubpGNYpj0cpEzTeJ0942afWVq+e3OuD5PLLN2Xvdkk2bdVhGBp0
tdgeMwVihDzDvB6mgK6cPuHh6cw1kYccpZddDmxrl+gtaLNmxyWksUxKHwDZb5dR
U4X4nMHngzCxj7jnwVBpJClva8PNBST+9Ve+bS49ezkM3BEM9gxUkp18XwUOaBtD
IHOx0b/r2TUjQCV9HwLELP+clqwt15vxQpbh4FJ+kKTvy9Z5AkyCWlN+8DLJU8I7
ktJax7hR7OA4+3g0r2s0XIfRcCoy2/h3XcC+cv7G3Up9Wk5CQ85tPWi7DzSkEMnb
s3zY0LyiSvqoxgpqC6n1QEmw6Ww2zwI9ijdWS/7nrYYzWsTqidyI+i22/E+cqvqJ
Qs3CtgBHgytT5ZNFyE1l5iNAdf7S+1XbsBMve8sCZVyveHVwrW2tPVxGJecFdC4s
p6Aur6+wnPR869phsMZraYya7QaFd6G2GmYSPmfKTbxlWBy19JdW7MSzD/8/I3vS
O5aCaQTmwTnqIF00dOUoPc5ASAoW1b8AHuCLYVizpGhuuQr3aJGP+muJc3S9TUjr
uj8twykwhp3UHjdMIYIQpNeqV/mpQzLWHq4s667eVbU6v1RfJACe043nW32MT1RC
gkOENA2A3rs3wUSRXT6PEHk/m3YOenCsabdoXgcjRl/01+kLatiOK0dc/XS9H8My
iIBivRrzuzLVv68SAI8U4yOQr71bG1jS79xu3ekBH+fhReTMWx28n7SP0MX8SiK7
rM/hJfk//Cak6veoxFWhXUv0X3slXJNzmRFlqH2ZMjFJ8pqGZ0qWvDHsait+cJmQ
qsW7BpF4gJMn3pNO/sfw7bAj+8JfD8fy1SLLaDRkrBNcKDCKR4SGuJQDXYWJuM3F
qB2w1Nvxp3mZUlcNfmaMQRQfv84ZV2X905WimTvP0uV7EQlPAcI4YjCUjXGZ+6UR
9k4LNdwP8b0v0R49/vVkS6Fg7x5vhRofS1WVazyc/uxPamIbrAKRd8/h9X8WSIWr
LLYC15LHAwl/3E2xXGV9+f3yx2q5f9NXENckfanaOvRNW+ZVvpnvQ6u8cuoE9wmy
CKz22OLgvcI+HdE1ZvJG2wMbY/gCKxPj7VonBo3ftJqyJEQLoMi1Nk8rny6LUPUu
ZEGEma89GbE4h0iHrwINzJ9NZzXh4/2VA4McbaxXf06tK5JOWMLMC+yt66/VHBAA
0wSEeEdb19iGLngeDGC6T6dtv0u13ZUWCvYlXisyae+1jEQAHcdYXvJNVtBwjJoj
jDKpsUGfRNol2Jk/Qbc84zYtUKVnuSlALiHh9m71k/aD0Z76qfsvMJY/R7r6p6KB
LXZVuY6RV4w+bF/jLFYGIUjKrTHUO1bIScvGynwQ1Jrqoe9EhC78orJK8mEC3z7a
qKAbyhnjZCd7igamGN+AehDX8TOOkWMldqcwkKXd3yoWixowFlV+ufJC/jh7A0oc
pTXWxObSr5/cYjtMHkIWELRIZEd5nUkitS7174hRyiSqFosWItGEqZJuAzAPhdKa
SKsSVEGM9/svvwwKGdsMfmU5MeRUGlL/1ZepxgcAYaQ9sgr/ZRHgBOe9AcZy/5EB
vuse97LBONgfaDrdPBFV4oDHwcmNjlh4Vqm0uc/YQJDU08HU2Dc+dcuyk2bl/6oh
KbAMW4W7T+Zke6YlquAi8+4XOiDgSR3U2io3ndarhDzxY9AejjJ2l+I2SDyH1dW/
fr+Y5gBDzErAR9wG0AA7+FpbfNj67AC5I+MGcQLKfQ/vdNzHA53AZ/FOoQXcumIz
FCrsf9wO1jncSVCjcaMOGZbohjc5bZpd8Lokx57Ftzwz2spLOODlvP3AHxpLe6zl
spBXfErUlZ96IXNGiQH42L9C1zC/9Ym9vgTy7B2L8UX/8xdaPs1WqN2VDJR1mA+h
fSU5VKixrI58uAa2SEEdYG5S58HR4+QLp0Zs2rayU9EeYTSTYzCqkdDEbOyGz5dq
sOW8ep8AATTMxAWJl+d9yteYz3kijCX7DakrgAddPOKepUTIf8SnPy28rhFmsd0t
oKPjCFp0HA5fmQmHsCCbOTYJUpPYb2pb2IsZow4wIKbyqAO0XYEMJ60XT+s2N4+V
vVUWYDXlZzjVE7P7CxJ2o5K28q7X4lyMInoAbcZxU4JoSyThx7TV9yQQ+SzbWDjT
3WXnme1o0BqEL2Wa7nHizmqbJJhXDPsNiLbInv1yHoSP4VlTzrIdBH0FwcqEXZjO
lue51GIiyI4p4DGZ8Zio/ISVvy4fwF5nWh/Xyjtq8dREpdtojWR9kAOrnDgvxtsN
eMpanh4iHEAS1X9k0PqDgS6v/v1atHLvDJAJF4AMGwTc3tUarGfJFOdGgDPiVKsH
kNkTPlnZvcA+wc0YkTMLDxLFNlyp/z6gUiNC3x3S3KHVMt7aJbYqPbuJDcD/hLOx
SQIn1EBQ6whIdAMeAVMHZlFWt/uea4nCfodyDxGAyeis3OxRotsr9LhDKfGs7hGX
FohvfL7uQeJwSywc/rDq+z1jmCJo7PAM+GElrh2P7pPcMzDrDnb/2oF5p1bEQxt0
SgG2L63W9D2nje1hKNktGco8IX91RZOaypCLsr5RA6sTbyYJJziPoDH01JQ3aTUV
r0bK2i6pkmmcqA9DVFObwNtqa88mQAEhdaRSCcfAVsEq4APNkcivtVKwu2AYNxsc
OXs65+0OFPvQF3t+qmJ6VXv5K6qxP7ccL2lBxeJ2ILBgDDYkUBolsQaTq4MXdmey
UvkmZY2be7qbOfOxR9ScVXs91DIfbjEQU9wktEruZs1zZvwIWLVYL4eru9vhtJG4
4gr/Jl0bzyrX7WwNH+J7cePVtZsrOrbYXSffDWszD3r4j/Kc8zy2EQUyaJbyWl0Q
PcstsMtGXP1FfwTXaazG0nG64TNCJZtiIWPjXQJzRyKWnzeCfI+wanZkEEIr9XRM
3lM19krm4LQ00aFXFi3HIAmcnDDTyb1ofT+XsCTiELQgOZlXfu3fk+OkvCMHdbKa
a5Fb2B0AqY6Ku6kctlocec4Fw7eK6zGO/qVER5CKeeagWfCU/8jeLiwDbgYWRInm
f+c9n+RcWx2hmK9OruHHa54jf+e4k07xQE3bC3sa+e8aTlTpoUqfT069EXz7Ot5a
omZvuZ9ZgK2520ilIpe9y/1dPvlR7FfWAttKj3vlrDbuutOa1LSVFYgojCRPFkks
fiR8Sylab2yWPgHgS3l+5OEPefi33Zw9LmRS3e+CtzfawkLnOmkoHL+Sx16gHQ/3
4ENl3oA5TkGBn6tOFzri6NYNLZNRI5Qw8kCkO6zmz/49YnJvNoRuTj8EMjVqShIa
xO0X8deLdd28U6C7pqMDjW2qZJg09pJjeH5KyCre3NDwoVpwpMijosHFmjCedYDt
TDhBPUrtyFqu8gmZZH2X7Kee/3kQCD0a1B+WjIl+4HQKVCUQzEH+xLxyyZISOjpb
rPdvyQbh4ipQF1k9O+dxF7sJs7WiwqrEE7mhW9eYyLhqnky4HaOuCxup8Y9asOEk
eBv3GI/tdPHtUcwBpIy0zdc7cn3OxkzfxwkGSdw9LWlOGd+iXJebWd7kBOq9xPAx
LrpDn4q2mgdYfqXBYkVc400B8dZfPeI+9GLaU16DxqLPD57PwiSLc4dM8e+c3XIf
hT/DFGUxv+Oadjw2pPAhdRh/6+vnwbB3c5zJhhwekhtmCqHBs7Hhy9GTDM27fE5f
yafM8W+3hGUPYqwp3WLHHiW4BM1lTmpx0USXG4JfZ5mLub7AHzEyWXvOlqitbpr0
4OQ4iLyugNQVcZwE8G9BQkRWfdW/Kts284s7cuJQDfOIMxTMRSPR5eraGO9ctfAe
QzuwlrR0EnSjD56NMh5y5lL77jZlq/47Z1Z1tWndInndD39XoKQutdHMWjYVrxtz
GAfSEvTscGi/91zaTvzhwmN4bVdqakCiuf4Br2mCiNf7hiGceysgnLdyExoiB5dS
phHzZ1bZIQhOpv/lVqsTqb+dS7zZEjA1sHEb1IUUswwHBpe22uofv+cmBHR434YF
xpdbk61hOAXGNjHQiLLkpUkIl8j8evRvM68e+vf3lOaAhLAfHZtA6qRHts1pxs39
PPDRDo3PFhS169esWwJmvGPZWAUVg0aMLIX/8C/O3ZF5hHvAbDtIP3TqoCSMI804
bPRUV89de9/w91RVyARZJiafGypUl1sFKSAbHleJVUUnXGjqOjeySRcJYk3Iylg3
kHTugZZupMlzIVrhOQyX3wNVsxbDqO8z9I9wrUWSrS4uAzZIzDuXK4oJQEcfoA+L
f8qdGZXuMPTj4kbnHpxETZ+ciXgkP+9MCEupXB4N4VxsuuYNi5CSV4RbzMSE9hNH
J6s7D2xWI3GKlQswToCb5B++A2mKQFFCWDO/AyfYuoITeMGuFaIuKm0bKl+FGQOz
3bITmdi+bpA8EgoFGuEcdmorc5/uyKUkDjumRKv+IPbVFyEF2QRJDeX/wlcWd/B3
/uVw32Ytod/lZD1eU0fM/HT4d2+ZMrYw8wm5d/xegAjp1aI2R5DEzeQwL9ZvS5CZ
0WDdm5vL4Yrvltj931oQ7BF+a8fjqoK6A0syGTcDWUZYXp9oJ9uXPT0L0Q9mC8aG
PcZQgFTdhQ6D3RQ0l7Haa075U38SnWyNJWPD5NbSf94qin4yJiXxBMhT3otdjNNN
VQfmnvgzW422q3Vro+OJDbf9ZACO1YXJHob5nV4xkZj96xP/PwTLgguV8nSaNBVD
ysJT5pR2jIZSqeCRqI+QzTg9Gb1QYFB+qg746jp6BE64gRiugk/A6SUOMkECTcyu
58/OXl0Vo53is+Lp8ly7mWYHHkn/ONC1vkdX0ZzyCf5Jt0FOc5vXe7qmfTjU1NfK
8YioqjvXMgAiax/Vty6ER03Nnzho84yMYmEatVb3lx0H1S0bxt99O8w3nesEXboZ
Y3EYpiXdfk8P25lJfz9eTv0th/5OVdWGDZvq7AnpoG8A9bcNrtjdx1TFnIVNeDQc
1c74fTBsFCcA0i1ReSQncU7+JEZr8cK/W1KGzUYvveJcqxrgCyCaunAJxavAdaDV
afOBqDQjGT5lIUF2B7/x+whzvpeU4vZJGNpbxsqHRcCxdMyXt4HFzmJyR8L72kau
GnvyUE2+4nj6Qk1K3MRF6Nx6wmVdDF815SAdeUDEMn8obsyToL9zncbnwz9wkuY8
8HCspdNcYqz/82v4ZiInW/UNEx5Lyuzk3+z6JEP9t5t9ka7cKJA2NkUXN32iUcqt
j455iOKuQ8tG5dI+70SNjR3rF5xDlwFaeOdxrTWx57RBm07ekmSzJIO6bbyqY910
31GsdTnxWOH4BxKMaw/WBpBzjedK72zyD4Xdi4lXh8oYe2s0lqnGZRI0m3DrmdTz
0Cg4gdrwbi9c02EGzaJzDpkplG1Ic1go+LT0H1o/vRGgx7P6RcM73LVv2/sChdzt
YuFDy1cLn5/tBs1HtFs9wg==
`protect END_PROTECTED
