`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yNTCciBrKGQm3ed6I8tQjRWXepGu+s3v/C4DuAsG6kq3Gon2kHzLf2+jXY62o/UC
LP/zlYimi5U1yCGvgNAF6SedEqHMCJMIgvOJeldnBY3vRXMtm3IzWqq2abo/ICyF
qird5M2Ob8qBkpsRfUYgcniAjTh2psGbSR6gbZE152PBLC6Gri5OwgKZsClPlQlM
9BcfmK98z6N8/LWX7FYVydbw1ZbrK93UoG2W1UcibC6H6fHV//GFwVOiTnzsIKgS
kRy6T+rx1yfaRZ/jsM6QjtCqlhjFpp/W955vnvqX0SbvBB6afZ7KlwOgZOua26Gf
ibKwq731S10h4wOb7plup7VLNP9nDvwKDmUVzn7LCC5OIiOgNS+suKLWpx9VEuFJ
e0clE7CTuObDYtPJEFl8ZfDAgIU4Vb2ULJ1HWzQ9AzEywMxnR1VCUvY737Eia8i6
300PecjVgtX/Iqh161NfE+Afsio3OvNSYIx8xe4iBHQ7qreTRcv5GHZsZfzdyaH8
1uu+k5Dtj8jFAo/A79lKSDcODMmKly79lvRqJwIxTh2u20Dvhhvtrq5MnHS9P7rd
cHbnK1dkApj/tfDhkEvLFP408P2X2EG/S9FKFb/blPjZkMSODCB6NYieUb03ydtl
BFT2jMMSn8oJcB7oK6zdbZGV74BXF5A719hexpwpsNMLzYlzNSAKqRRNcKZDrkVy
ELv5WxfJ7kaqbTFPhhFjYJLJu8onq4iLB1MmGlNryiVT38nyhRx2jyhEqv4nJPxn
Ypeo0rUoqK06FrGcU5DQ2WixoXISIgNjN6xUr5vACrbEcgH+wI6MIj4r1Ja5jp0K
fswrMxsI3wvw9soZwOEs3NJvhK2vRT3UXlqI2P/nCHkpHJH0eDE9VnAoYRe2S/5I
FpfJ5QwUbHXdn2JGEhjToWsTKKquW20/okjEJ4UOUVU/X9cafdQ74et1SvEiVA3r
qmdw875We7DBjfe7ugmb9UZaerh8qJkQO66XfLQo0usDkqoQjWPU21p5Rc+tIoH0
cZdOqC08h6zBYaMxGwx3HFbD3LhRqnEvgYqKbuzGLKnGSa7QPx1m+oFjpDi8BqL6
cI/taNJnZpDt76AZyUbvQILthhu0jGEqRwBvbRIl4gbHt/HwEKFzV7MFKG/PLGEc
/MxxRui93tuWFXuo3p1HjZCkS3/6i2ieMm7gJEkDWe5QrdzosTFOcwbSR6ZGEqar
XDZb/NlOp6By/8qSKN755u5PWd0bn+UYlLMLR3exsTo7Em3L2NrlhaZRyuJfjZzz
5Rd/JIVYkm8Nwl6uWY3TH1970/CJbafPEiaXKr7e3YvLrPJJaN0zNSv8zXXg+cTt
ZTKgtrkAfWmCh4ptYpChecLLmDXbvhP0eUXvfL2Zs69bsRQkFjEqZfI75Lg6QO+d
+pRrSmj8P/yFP3PH7Oo7dW2YjdbeJWS5lpR3ttHMhZyN2WJ9wgsvcIZX0bChLhPu
A1yL7Etvpz2y657Ro/nUnmjkuEXNs8SqMVg9qITbhkSU34fFWGuNI2uy8iu487IO
9SRT4cuBD/UsTVJDg1s//txqtYQRGw5fvuImVUy16lFL2VNjl++1ARwUQbTouS0f
zqpru4wSqzAfDv6zvG5uny5vAMIDkaK3uL9HtSvRkTkXz+eCBuXnBHTurjPBDpwa
W6ivoZt9vnK2+NxFT34vP+RLorExxTNalFhhvNymbVKI31UZ/NzaPt6MPK/BeOMX
Oy6bHbLngQuX8IAJanzTjaqwAP/y+5AJ40agKhwcjnuXBdl83PqcNvV+lfUvSQHB
1kkSOkmVhTCmZnqIw7Fjva4jjgbLOq41s7YUQjVVM9q44zHtAPvNYGWAGBY5azg6
uzZepx/wKKFEX7HOPMVz5VC9pP9MFtm50bPTEFqD0raU98gvJT46pj5aETHTzVOS
KSwymhYOT9ohy1Qb6UqXlYjlOlMForUf0o6p8itcWrod3IdLLOxXZEI3DHwHgEHR
qeVDY9RhBfV3lX6Qf6OnPdw0aE0ZioSLPJgby+EpHjy+RwB4QC3uvRe3oyRCeR2L
/pNil6lTUmutDKOL8hUBLt+rvmB5iKjJC75n8PTPxkOxW8jXh9dSTn6UWo6yXbJj
i6RhMz+LBJHQbdIbp9QIOA10EOS9RL3IBB7TPUar6JOCLxbTIa0k02xFakKKmoJw
UM1j7RioX4XEomR1DhqOADR2hfctqhjhXjph4d5yoqSB4xlClGrP/GyVI9w/Qx9j
ux9Cpp454vsrZZYJbYM6Lt5957kLXKQi8pWT6N2IhH5qQ5hM1vXzGf6R4mUiYPbh
HrUsBKbmw0+4ouVVHd9C5fojSQRWgc/gWOFirCiT6Ytx+3hrOA/ZTSsxRGJ/4TFi
4BqfklJnbwBl7K6itfNnE+UJ7wbAkONtMq/q/hFtm3hg9IduE8qlRCrSbg+oBdB8
B9Jy0AaipNJwFfzXaW5/ENcyOLd82tCUrOT+EHfn6ozegKFP0IEuTzKF8PYsyeEX
+CayB6ZYBRdoAOKqoGimYc5jly5dPW2GmlEL6m8lmbPvhX087arqpXfmJua1CpEs
iOlysq5VWm9wpU/IAA0rAyWbsioOVSOZZYMJWXz+6mMucuYmcJXO91EdE3+tgBmF
nwXuQ8yYQlRvHaZCLv/yVkgv0SoFzl107BaHYumidbk3u8pEp4s/UEfwqV55jTjV
jPq3PZt/hn3q9WIi4ckXDib++ruj3NXiJ/KGCysfjxikss/Om6Qq2CEdRV0JBbJq
FfwuD10NYLOU3XECj9930+7HZD0M3V2MhKv67fSFq40BOacUji4K/0+NGieK6COl
TkzWKPm43ZRvpnWzJlzuUcxlU4RhvDEShTJbpkl7JDcfPYim+BYw/pfm6RO8SUr8
OkaN7o4nspEvo3mVrENFCoTQjiQ/MuHFUGGdYF4D8uE=
`protect END_PROTECTED
