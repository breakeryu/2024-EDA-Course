`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OrYggdYRFo9LVa/2E11+BkNcIJ68XvKSZifkuD+im/maahdSOxdsnbI2/uANjT6
ZS4ATIhQ0SJ/ucCQNRF7gBe9bZu/rrWpPU+GqRW/3aUryyaZN7EBbZWpw+cDxTq6
tzsckcdpP6KyGh5foWLOETq6WYLBU6Hv7SianfvupUWVwWD5n+O1/rCDNdqIIv42
zwCsygbbDfiFK8PO+wHoUgeDpyJ+E3t349DG094A67lINstwmf6RM/khra3xqq/A
RMrutzBVOCdZdwjOj+pMaGuEV5Hpd0KSrvWclMB0lnuWjHilUNGfXenLB5GhEDFz
MVMd8IceuNVka/MdWmmyU5RblRskxKqAfxv6bgWCOHP8MJiTKHDO673H/6oyHmvY
I0qOgnY9URquaSP5M6UzaptmPYWq5i/y1D9BpmydnqLsb08/8L5B4TD7f5b10Xuk
mBrA7BjmenocryU1LDUM7MuKfOj08EcAZBK0hBZ7KK1i3KN4RUWa1DkHG/dwr0/+
fckwpEdjZJh+CFZdnj3kgnxEvUmyxUL6aJGM0BQa0u8w1TMDACuw26he1PFP9ymQ
LpTcNZvUR/xHr2KDQ9QIzxydEANqYTfm5F/TxaDEpCCOyD0ffPz2PZZ9iXLmilSY
X5+tYXN4XBBW41Kdj4F9XUVNu/I3fmtWwEwyz2uG/wO11ZuaqMVaAOdt7H5s1grB
Cy23sJM/wbD6lmVxJNA8mh9V874E877gXwjl1/eaBm9KqO2jPzrIfJE/e7Bluq5Y
xA0Dh+JOeu6qtootFrwMtANimaXfzcY16aj9iQwhrnl0xH7Kk9i4SMY18mXsyqHa
Ukws9mAhKfa6neGbQ0eO7G3bEW7kfHbzq4qrcH1PJx1VMkCeWKnrSlxJNs57Uq47
iTI9hD+IunHDeCAP3Kzd/+pEpLQv/UkSFSDOEzYOzNLX4FdpR0QXqFYryHfF3UwQ
/5GTCZCx0EuayrO+MWcRWhq31uywBfiGen53rrb8cT6v64yX0H13amMTJMWA2Qzv
wEe0QSsZT1DvZwLY5qLkbVFiAV0Q8qAeeXrrZ8Eu7ysIxdtHgO9am7iqeMm/BWr0
RAiELvrrugg5dnugKki0iLYubAOHgqoeTOHq7yiBQ9Kia5xK93JgWA3vPt+cXggX
YTAo39mVb+OlRaur/ZjT18+HVGvLTHvbhkMfXL6T+WFgBh7Dn9ZOetwOWk5uoJQU
UAhX+qChtvCmUHSgvAbjH9svEg2JSOUU1pH2bL9AaWOzxhu5tL5ibQXAy+B5YOMw
5t4+KeVqEucwjPUYydTLc+jCuErJYfp+z2hrbJl6YXxnX8FwbhbnrcnK8WaC1zR7
w6ysHwCgPjqBQtoL5qd3sPevxVjKa0WfMjb8WK06YOrYQ90x7aTomhH2RLgTOkMq
V2qVEtnZv6hGqEEOX2AIbXLQCpvenvpjT8RcFZvTbnh3j5s/c1WYPiE7VM7CkFGz
FSBu+WGvfJBh9NO083+3L98cIsEmam4WtZwkODLL8lFSZNegBO3DRCnZ78XvVpgH
MMOjpHUqC1btyqxIS8zKg3s6bbOA/xmgEbyDGmokQQpivvCwYp7LClGpYocvqijf
392b0aKn3L16CG1hbfegkfdNF6IO4YIlq8kJziD5Wt0FO7dShwrDyJZK31gvTUEk
Pm6S32aOFDq2gQyR9T3hrztijIHMx1Uq+czr+rD1rVdwtpXdfJDY1OtWuk5/JaD7
7n/KgmlN2rq8RrVxAmEtmbeGOgafwkUIcKTukNIRYe392bS/+PTWKoQZjm0VV8/P
4BTigTNhtpe6VpvrRy+R8r8f4Iq4UAMd9D3wQNyTDIT5iR7K5sm4K64A+Q3gvL6Y
b7zhqfeUwlgR8a2tyXemRIQ86yvtuKbsr5QoxyZzb6wxu0sVFARGh1Umr9hXc9Qw
njRyc3KhoWw5Che1U21zSHFAv1bxB1N1VeljpbNXY6jEEejr6vNcJJzX4M8if7Nh
1rzuWC87BKu1oNRQmNvhzscdqTgDSKkDfNX2k2goHcfKysrgyf0nki9xJgYFa/Dh
WKkPA74jgEK1sDPoaFZBq2Q/QNzxG4qr40PdAY6kCluuqqYcV7Y0GZh7uH+eB0mL
tufA2czoCC8s5lJrtK/lZSMhLYUnmnNfPphJEwNYKQPxkOL7gkm/v54uSu5V8udv
UCASu4mXGZ6Qi15dExc/DZy9pDPpCXkmCz0jnelfL092c9vfOHsN5LcuNK/rkwfw
RCFlu6ozH+mB0wqafT+NZEm5t7bD2xszj8w/Xi/VVpEBRZuFjMjjhsk0qMoItk9u
CERKg/U1wSPZwdkrCFIZMTx3WEauEFhkgUN/x/5DSHtEQ+lTOoSuWGF5HjMGbmpA
dqt6JTsk1K4MJOoIxmfW5g==
`protect END_PROTECTED
