`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9BKYzbsCSngLjQsE2dIJ8HbM0j+MPjea3PkVqOQHxiWyg6SKz/1a9riJL2TQyJo
5bjK80MLPYBhoOTSYnEYr8tAYY8knZlzqlDoFxhb/g1wMWoE9D909R62K99y9X3L
rUdWVUvlPMMRqMD2iUNbduIu2och0SsyDo7nOEqeExqioO6jOhZDCtD2uh2vpK7P
7byD0WQUUEtL2SU2qomNa/8rELYh/R+iWoD9OQ+/8FL2UtdEG3Iayk21P/f+ycOF
1xGjk0Pok3h7nJeE2JNYkxRqGdzTuAJwak+gc1oEN0MaknWx8n7M/LGarYWtFGvG
ZcP2D2R+akAUYBjs2I1tBoILQ5+KNZw84qCWY15C2b4DjYGOnmSioNdbj+JMSUmQ
UyQajuljFAJIANISIOe6pbI1rrqsmx0Im4FlWTZbIPr/nkcY0yKzBArzS9zCt4Xe
6Ea3ooNslQ0Xd8ZqytecunqBdq9q2mAEcuEl8cpY/Xegpv7Qa118y6XRsOmIxVx2
cHnp5whUBBi37uOMnMOosnNELUczYNIDtmEbHv7ZpoHPstznlp/0K8samTfRC+k3
7Iz07QaANHmHv7HRLprMKsKD6NIiap6LM0J0uV0BSIM7M7QOMZRBmncMwgkSV+xP
Y3nBqcME3ZHBzylwKZGptOZwhucaxC6kN20ToL/Ljb5z/+WMUYC7SeQXvXKbkvd5
FSER4sYcp3Q5x8It85tPpbIhTWlXnk1e5dpXV+DRb3ifxJz8JIOCAKbkg3WtWx6G
rLdY7+D/bUtRqsm0kT+ZvJxvQtO+WFZ4qO5miYqWDM1VFQYL/yG+mfRA47JtL0pd
oWlONfiYyWh6pGw5XzAfvCBDwuBlTktc2HYg7znsU7+PxrZv8FM1qcnwrCqb7SFn
T6waWxixwtLVk5QL4s4R3xweTNoJCFijOPHNh7TgSoxFWCuIt2STzqCNLhfFxKmq
ylI/qTMA11MbUAocPB7xS0z5aLuJkhYu51TcfkEJ666+dskWOCIQtQ9jNT21RHO/
ZwRLrwtTi0m6XJBhbTER8znHALMHqMyoFrGAmI3ogCaSe4M4NqHvbTxEJXW2xy/m
pXNj0QHMUvs2kaRfb3YpraGYmiaLu6dxq3A9T//9irTeg0QtiPvbflp7S9ib8Mey
G80UV7yjl9VTBQB08TFP2jqYR/WKfBm9RPg9+Y8uFcUx+p23+Tuvhno87Zsmgfvs
k5l5w2TwcPVyCuiyCzoHcvaxVBV5M17vWW/ZL6oFcg1VXsf6moYzBhrmXIUuuq7x
OGr/kQLg4EuJy99s2WU1ZZVCACjLblysyJJJ+xz5//MiAg3gclTaNiUoZDNPVgOE
sQm+hNr0isbJzX+1i4+xl/u1BwNgY7byF9Be/bjnHMYnAB34RevIF9kfPhF17INW
iqyM1GfYDY8WyPtsH8yNmaGvBZ1K8J4q4T6fmps9Lnajmf1/V89fNElLwzBJOPDL
0AscxXbIIQmBLE5i6iko5i3NtOp39MD5EXfEVk+vJTCqZQFfjEktPeRQMEoYlbKQ
YSQsfsbkDNG48qtkm2b5UYbdA1x4ZM4Abg+QNisBiBDRtSVfm0g3NjAd3xxfy/nB
vuNe8Q7J07CF1XVGAsa5iVhGLIFFkXfdNmp9lBQcVhu3dMq5lem2s6PF6bRVdXRC
351RiylJs5okGUrcqfcK93gIBrBcWANgpVJi05cHcleTjLW0gCkhah6Q6sXjTR6g
dYyPgaKNvBTCzvbelwUmM/MW3bmh1ir+kShOcI7iriu6pkUzcUgBheD38saAPGpp
0II+kKEJOgPmlziyNt9+1uX9Mt8M3w0opsQQN2D5q67Pmq+9/dnfJZaysX4GUsDO
1VBZ3RTBQB8kZ8n9LpYNASQoRfpJJzNTG9GVdezYsBnqKX6NrzxpIFwLPjUV++de
0MkCaP07Df1bhKbsJvdWWB6S3g824+o8akFMoofNXBgkqaBfHzbFe3of/+PEUf8/
o23GCbvTMNR2K4tYnZcvBkt6669eBMZrC83P8ou6pdHUZx/S3S3ALLGmpNhlSAuR
t1B0hkhQS/Teg5UIGPrBDGc8dfAqcTQE+a7avfAMkf7RHjp8EqY+5AdGazhUlFCB
Ek5Ru167gyRbkK1TBduuGHA82hhMEMWvlJqSyPZzeneWoVubrjASA/w1AEzEBZQb
wJV0885ClwE//5hcOOZjXe/FmtMEnjwoXBOBBiMyWExrVeL+d8loCuZeVUbUmngO
ZoF0FAR36F8LuXPZuDoTHmPyQp3srvIAzmdfVGIa5SmzExQ7D4DdVHwjqNMMfBWB
MXMYVuGPbEdrAEtGFr/6lWgVSTxmAS1i5AsPHW+nhyDg3aCJtSp1fWxCzFVbkafr
HA4xCStEp8slfATIX/wq/Zrz9szrKDoB/SCRzLe5vKF9lJnnnkUOmwxxW6zjM4V3
tbZMF3J0Y6MOzNhCvUEffo9gMEmWvVfBtZ3qgeG3g9wMHn9HP62ZkTsPtnLdDyHn
GXzX89vXaxbaWOwEj9fatoWvaBXvULsosgonuB3DtfWc3j+PsMkTFR2urG46Dj0w
ScwfGPYnBoeT3MbON7Zz4KarxbOns4py9QfZBCxm9gEYrJGcTe11OsPsH9kcwJAW
Dv0bP+br/1lviU1++ToSWc1GlR0tdZeh6LOm37BF5I1hHqrAbSuiTi6RTrAu94I0
PSsyEnaON+pfqc/2s/HT5HyCpujhEwmkg/oXZr7x1DPiyjij4ULJjvT/rGtJ+R14
/ZMdi0GY1eXDEyPNs7xNCOb9DlVPpSsF2nRqmgocfX8tR5HSzkzUNQIeQdZOxF9y
qE+B3GIploEMteimZKsFpHl2RGGE0J75wkHl3yahxpCQJncSF0pZg0FIazmFMS9L
JNnZB1qmMMuLgqy/+Q7mGgiMav+9Fw/UE7yRV/X1rgtT72bLTKErQAkz7kN8SaQY
Gy3F8rM7OJn1kxeq2b93KKkn0UTC7NkxDjF39OVD7cklUwEK/u99QpYPKKM8EJnJ
Xgq5hYlAf+kcw8N56km9OivxIPtDVmrN87sxqZSjyp9RFtRBzge042Yj004NySRz
WN8vCtyUCdYoXhBCdSj51e1mgp7fgz1N0/ps+9pu0dnURxYgySzsdILuK2r5Jy3p
glIrQzNWRXX0UldEqE9saNC3R/LVJd0DFjWpGol/1cYlTwzSP2PwdrhvnH9Jd9Yl
IbIiQtwfZ3mnnnYeCl37q+LkX7Umob7KLKZmlQkUnVhZCXvSWGro10vBH0OhwQiv
z8GS0xugbvDIty+M/kXQqbnb0fzV3efECwaqaJ7ZQVv5NvdtS6hgPDQNWGsC277M
wOUJPTAs7hfqvOIenL5KVQmbjJvZZIncdYgzGimLv88bJ/QY7vT+QbQ5aYs8qzWH
teXqbrd+Fk3ZcOP6vgjFNrCB18LdgGLx6s0p4iuf8fkUZlnMAkjsWLWKzCA/lpOG
m9hSnGRH2tSOUf/BeWQcmwa/Sm/NGyPnNGefl07W8jM7jDXn98zIpMxrkEJMeHzc
ciYWZO4UZLZTh7kzC28qwPD9Mq8JSzmmwIrxRd+krW5fqbTMivayYf+b1Cr6NL6b
O5ZU+uv9il61LgcQijRt1FOd2+DclUjvIXO3XDK6ZdyIJ+YuxRWHhn9Ie8Og+7Zl
tsR/Pu8lZLrCpv1l2zmMVy07YSJudZOZ3hpmxxSzSyHcfj4a00H4XTb+7Qresy4g
rY0HCL5F0zHQ/poHIQ+EgNJHKqpZGdKgCENpQj635V3mB2pETtFVgwvCmK6KxGIi
+K0xPgmU0T18yFrPOZysbkh6+y0xHu74LTNFhgUa/SCSbcMhFwip3qi8vkJnO27o
fNvCTocsty7nzJz3om1ykvIiHyW2cRyv0mu+NMvMiFWVI15SAr1flThGdkh/tHUu
NpazuPp6GVF2H81JqVBZd9El9M97AiTW+3wDCeEVvThTCHuH/VROcGcWUvr3dxPc
u9gB58s/RUezkZtmCstYOJHvYgpu+5lEJRXFURkJlz7bHG/PRdxbo/9NnjMnCmPS
oZIfqK4FUaHoWsE2z3DL+htM3YeqW4t63dcwKsckmftgv8xZNy3hqptWG5aToGeI
Kk4H5YYH7KBoe5W3Ld9sZ93VrSvCaZ3QV0QNE43JiglML7RG5FJHXsEMUqbFz/QB
o5zLYGlDFU3BwMSrzqp/evUkZk4N/03OvgNfAfhAoR5Af7y1OncXNL/f/IWfLBu7
+hwj2UJXMuidrXhFiWmtOkCiA+LG3A8M0GqwvHEO93zUSEstdGrj8RkMSo0bTCaM
lEc/mcPuILTWwfdMEn886FjdCJ6GBQFW+E/z8vlLeLiRwL+41JCRczCU991yvpuF
L+si1xzwEh1dm6EMji7d6vhKV8Uhld3J9WupY53DBNlaNO8eOj4Eby8vz/RWSMQu
3HL984j4LM1vJgAC+Ii3FWDLnQrqvnhXkL0nzdyGyOB/0gfkkrKEwan8OwiH3wu8
ewB5hVYk1vlBXSqBXdX8YeSXgdakdMQE+rwtiTAy2+plpvasaZ2JPjs+eMvYgNz6
FY5f6P5UL9xWIoFMelv3PdWZfpObc0h6Ijt8ECVUEljq3889J52PGQj3jRenW3TF
azrMyKyKRYNTx6wldeIeYQamBS6H4hU2yEhpgIr6DL/gaVXqSqE+HzPrtIlFc9MQ
618GLe46KNQawrg3yz688Cf/DfzPdasWal6mnOlqGJOHUkWpu85xWXJVZjm4lwyt
XuCGDRsMTTURpMyn/gN+rysi8QiPz2Wd6Nesvf9PlRjFizMWf2iG+boNqAO6Ikir
XaMgDPPsVKHk0Ivismz406+ttIN4uIWDEQ7A0jAWKnmYXw9qbtAQG58ckk7Q1qVk
mpyQaanO+Au9jWdtmWmUHoVvL+5062FIS4AaMqWdfwo7tT9XRxiIs4cSj8JfJBXR
8lJ+VrO7I2ltwN7S66a7Td4QQwmuY+pgOBh3Ao2tUspxTCyge45cMddoN/TJG2FA
edZMFMtLlPeHFkiByjId0QcJD0wRpf8CoXknVy9y7kqzjhSbvpSBSjdI3JajC5Ok
3hCsT6Y7+OuC2K4m2oJy3IgQ7MsMLo7zgLOtaktljYdeGWVyjGTTkAYOWo5PW55c
oLLpOdLD3VFD8CtJEzRX56ILIygmVeWal1Wd8ggwOyP+6J05mAclCFEzJsKU1c6Y
688nnV+YAo0WB7RwPo8UXIvGiYzRsSsSO8CkMKyK5ZNdqsQ2Q3S/Jmyq47/SdfrH
0HZEAvAQ8LXTLHb+CpsVQnQE1gc0gryB9Fmnd6kqJq+mOLFK1hsR7zgLtKyONfIr
UpqEXjqLKxE8abtGqurz5ne92DtZc0gfR5+plfAhyXE1E+jbPldxTsF2lgUwdXnz
ZchSz91FTK8UZG2mYz6GGgEkzQ+vxMno3bMWCdtX6FYM9W3UcNrWYeprG5Zn14Z6
/1EoJZZRpmkBv0egI7TLhuFINnNzwySpq3fIcS5lOKOgTekKXqxgKy8c9atklImK
nZlbXVuiRxyyhdKhjwTOZ1rOOaUTM0LSFJKnf2sqjWBlYN82NXJClawr8VF6Hfq2
eM0wiwsCMci+qXYrKMY/QDchOReWlu9U3yNDD0gTWfRapAYz8i0Kb9LKPZotvboz
3RYUuxQ2IQ8jXZuPXGrtcU8tszKQtImFb7yV/qSv4xPSyyWzKtTkLYcNbOtEFwU/
QfxWPx2/87weAm4brVGSeGzkvKtp8GqCWNocYQGgXRjz8hRhaRfx5tlucU77BCC8
DBLGzPfwUfHesUXEmFrNGpX0q/KTeP0zOQr5xJT6xsalG+BXnX7vKTzY59gxD70k
Mq03PcgnVq6N/nBpAYmhMaQLDUDv3RcDomWwXJSGr2gltFnlGe16gK3DRCVDtTLV
lR0a9W/0qN4keVM/B2E501zAQfEiLeTvaf1H8yV4luPcPDYETxEYIOD1AyM46lS9
XS9rhdOKP+4vRUOcju8YRuT6jWwxBtNphVqx8m1pF6f5E/8PSRib+DPsvLWHePbI
G69K/sTlfUimyDxOxsOJnfYi7ANqlWZjMFOSyqOK4aOpnT9dxbwjFrV18nJqxnvu
bZphyQpyWevtmHBGFaOs+kOtKPa291aj/sacYKXg8+fYH2u/xUs+z8pp4KNuo81D
Mvvu97J39pFMf7n2+6Udl6DeJdgpJrWy1sW6l91Uk7lkVVLKjGE3OWyy2bvMFoZQ
NxtLqwYCwj4qPbg9GMrIBgVlbBZ+iDIkSvJ7rG8ErZvgKoIF6LcqXlCDR7ndRGWt
D7cX0eO77Soi0ggaHlcQ0jWo+Wtz8btRxNVtctsBuHu3fXq+oKjxcUZivVlHB3V3
cPQ58Ik4Iy3TcxWqbps1HST+j9iicwUI2oGXkxLVhHNbBWlSjKhbaucAKdPbQqa5
oG8YfuI/bHe7uNkjoqDa2Hjlpc2teNun4x90UV3gVuEcXIqFrEJfyPqwO82tZ1Mz
f4JrtAO41bQGX4iYDLvhla93oaiNHG7KOETyk3q4k8pLeU7VuzV8vRoB5lKDdaQq
asSVD327QMbYhD3gugS1XwnPHNExPKrZ87Ql2DvGcLHMi7j8xD4+PaXpeXYgSia2
+S6VJxGGXenxEfeyDEvDRyckOqbTBjYx0FxmyE3RzijbYn1s61gLKg3yAcPu/d56
CMx+G3GZ4hrgIZ6F3VwWy82/CnPPUjAivYc+JWiH7zsSmBOohfmemAmVGC/fruIP
tCRmngyMjp9nxLmqGU55hYFGV3YwrPG8LS4enlsnRaCibkNaulEKjkXw2Nddw3uA
+fuB/oUDAOms1aIF9FhWsBL2zGgEvbb3e/8I7nIhY57n8Vp9MulSg8AO3U7Np9UV
`protect END_PROTECTED
