`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4IwYDntR/1KBMXwDYnB+JvyDxHYkBU8cnve/2rkVORuridecM8PaVrNJO8rWXsh5
FHVSMgU+1CYjHiSCMkOizvVOpii02SZ49y9SPxugJftM6d1J7CJYLXibUCI18lhS
SkHvDqBeIRobn2f7difhIIrzePfwb5IlA2KuB/RM4dKQlN8mgpLWf0Nx4Cfe5j8d
8zr51PrYOme6vbqV/rLEBGRp15p9pEhjeYOhf6EANBwPit8ESME1J2dtcfJBYhPX
ikzeKCoS0V3wtGJnSDCtPVU6FQKbrOzVGctx5gfOMQY1uf1sSHHXo9a+MS4qMQIQ
qA3cRsfxHbaMyRK8i19GTzCZYJ1r/cvUc0RQcfv08Qgq8kEoH+63Lu8uCsemH0w2
G+MUJwF6nq7coODlFCvp4lfYrH9+av1sXXyWX3eB4CTrWPo5AllhXlc0/9veJRr9
d1yEnHhJ1T3DvxWfqjztowrv2Y8CUGknqwkf22ojhvMZ+vkm5wFLSch22W7Lpt8v
xvF0kDA5fzWo4WvSYC7N5Xk6/JylTWXenMtiSQ5HmQRXoxJwfd3Jq2vNO9Nbype6
VsOjs5sFJ4JSWXW0OYLChNSVxduqxKeShldTvr29rMT7OQbL3HO3nIhspg84jesR
eEDs3iI00yk1l8Zh6EvbA6z6rwpVyJYQpswcCB79Pz0KZ/0NCWKv5Lc7lp94NKtF
TVbGVmixJU1JUBHF1BtH7pC5ftaY1e52aOfwfjWjpCzXA6dQmUSmvJOCqn6DGKzj
EQODB2g4qGLzjSUQWX3YgA0y/ykvxi0cyIkRQ5u44YJ35av4l/sxzf0vmoeLKhG0
qJWu0Z2nZR+fO0+uHkHKiFbNsYxDD8Fpwjdhrk8IskNwow3g8JRC/m0lcgjLlHM3
eiM/jhTvYI2xkitqLxQT1Sd3Uz28NTbcGiZ1nL/Z5wyzyfNVzY2pfjxmLOqCiNr1
sm9ghdKJn3ACh4tXjJmIzUpR9kqTe5hWAhh59StWswIji6NpmPHUPOa8HHJp0hb+
F2DQzx3M3+xsdDvbkZ5imPVbG1IbFaUSnxwucvHZwwS7nUK24aICpehzfHJPextt
XsscMwMeAu9VCicsCMXB0OrI+Z0NlZguauuFkqcEhBMngraZh8RegM1e1WATWtme
Ix/QPCNb8ulGPI6fb1T2v4jYG42qsVqQSp+kSLvuNJvZske8l4g8nI2uIXnhMJw5
XHcmDQJ1coOj9LLigYt++WisYN7pK2rTvuI9AT0m87c7I0lvS+FTFXsg4lbJ3PVR
cR4ZlzPkr7otl54Y4jB0fOdPHyYo9T2pvNPqeDwI3UJCEGRvApDOgQvre83AGRDv
QMba9yvHFs28BQQ+Q+avzbV2FNSv+JmEp38Z+6ogUbWe5IP0fh6RkdLbLMzTNtLP
dpbFORkNJ1JpPqN6XU0bcyOfglZCVKY00H/pLCxqWmXscfVfL/giIxLJXjdRS9Lv
QWNMPkqS3f1Mi/CYa/WeDw3cpzrZ7m4GgycIMkB3kjaEmbR88QeMgrrNb4RIFHig
0IVpAYr3gZg/Y79MULkEnDeFEXT+CFgU7Sqd1nFCnNpJhuDa1iZ0eWJWTsWNTfiu
SkoTe/lkg1XfsfjHtG5Sa2fFylOp7YZBqFRYDYUfpLIteXbtoZwrAAMayrvwbJMy
uH/XcCrlzlw0VIWjOVtip05XQeo1mpxZ+G5YHZqCi5OBt1T4qQRoxx8MQyjhTHQL
qNaydFpRV+2W7Zwj1ku3sRZzfAzlGv0HUkss/I45t/rygEZ7Pb5IL820Y9lHSsKR
`protect END_PROTECTED
