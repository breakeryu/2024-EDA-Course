`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7V0Vu5j2N6QKSmmprZ19uKVF4L8KCp9nX2X+vnSlmpC0H7H0SNGsDxxBA92RHx2L
F15B3Mt2tGtSXS/FwIDwN7eCNOpQYi3jXC8zO4WAARiv5TbjzwYwQQxwi8ALFjBw
m1e+FdG4mDoptZh/mRSObSdNq0CEJdt/xH/KoFsIJc7pGxXj75BC3QdoKWzZ8cz4
zjFqL5vDzhia2EgevazRcfhT5mm2HVJYDef4Nyrvqc5PBnJYKd2jMnyuwdZcA6Z0
PRb2n2Guf16Eo9eX1MBcRtPwHCW4+I8VKhQutgD+He1BUpCFPTOt7r0Ml89nUDhC
/w12+snt6htJxDM/7c+dJkz976tIKDkSV1Im+rTLg14/l/g2tV3HDizaNO42CYAS
p4n0+Y+PmKGE0gIl9eseCO3sN6OLayq2CcoWupwqpB/l4A3LRDXzOqeL+AN+M1kV
InG4FO9L/MOZHEiNV+NXLn2rHksUlRWRwkjIQyPpRKFRABM0Be9jHcekh5VnSH6v
FA5FlyTcLB0DrIDx2O+8/H406myV553YZciN8/9TeAy0zNZuUa+M8Ii+PLcBoLh8
92fckli0OIuyQcbToeVFzk/ywFqTNRxvhb+LzGDjrr82Je+BrpgYJ4CCKBc8Pk8N
diIDEZYb8uOFTTMukxK/KW7USAG2rreRHTmrabUu3OFSxLLgRUMonE9wRavJ4K0c
sdn9itKus35Ph/MNcc09fho1UVU642xheYRDKKQ+FzvndGg7EzC+PYMsbbffaszv
ujsPC0w9nDieS71EJQ16Z2L51PCOfBy136xHSeeJfnIVWiV6zWGHJVsgWJLww9Gk
10DaIgLHvINyT7ekiiUg7P2W7PwGz7dWsQ5H5132aD1AuR4AO7zVcTdxjtAO5bf2
0WE+WrRpi4rjSzop2u5hmpefhupCgGjFZhnhihbmW5Dcx46D2iLIwXBlVy4h9Vr5
ExobspJjXtDP2EMKSMv5F9HbEs7Njod4vBh/J7QePEOwhpDdt9sy9p2w9UHBrWqo
SwtpWcLsRIC6uiVd/06KRd3RFKT7KdiUBqW5r58LFEKtJZIPBAOXfRL7p0/OyVLQ
ZWevWfFOJ9iiIrW1nYzxq1lSVM4lrb99nEcJ2OqFeJTvie5rEblo84sky7BiSKIQ
oCb68XRwiyngW3DQViIeT7aRAOvtz+n42gGz9UCeqZXa0htXkITfdIMz+EP2cV0o
zLstBAcT1K0p+MWOfcmwtJ9ZqFiJlwTguo3hdED0v6WiYCM+hd8UE2/eLxT1FFv1
+xQKCjghGVWNOttDwmS2adVB3GWl2eRAuPw6ScCGuBKdkb+9jhCZ6bqyLv89RMGq
ipFCG2Dx/Gp57bMwAgYUD3DdF+7j8PmtMjaY2sN4sNmsB8A9eb1yfJazB+5gP4FZ
qQgxVGdD9Xpoo7knxhY7HE+97vw1MOK12s+rSqvVIOfTWctPxH7DAHG8B42y0aH1
dQM8LOynjKWCm87o5b2FoIpJLr02VRtAw5WKcQ0G+oU1gwm7mrCScZcdqijPbSss
1eE0r+UbXTlqvuiINGeK2SjJt2nxdn38vaztE8D72IPGyATziHDovvodtiLwNdYK
nVKqP4sSsdZklALNbRWM79JWZqIvBDY5I1r1xDoKO1uhL8Fe3A3LbT6BSqxFWi2c
+PFslAAsSEn4OfPmsjf4o6YR201VZfJRfnCoYPmSYK9zNe/DPRZUGognoy+om+ea
ZOuBMnUqVaOAxezo7PyIobooNFlLX9bvlDrnD2XXFxPrYyKvNb3DM3GG3g+wcpg9
N6aCBvjNMB5mLBh24uDxbP6rHl/ojW4Ji7S/pB8DVIAR+9riTpdXIrO4vbB+gV0+
oTVsgHJrZTvvVNfdW7F0uO6j8srJhKfHK8KdPI+xnienK9p1cQYaddF/VNzwMboD
HEHRFsce97g/NU4WOS2wh64/bRI1fFYZKYP2mC1T3eHiQacs1H0ZTLcdIIGwhsjC
8hhnzyIBaJnPG+nTZxX+Ugn/HGmIqYlGognFET0u+cKl1TxLR5a6Rnt3TA41/54P
G/VbW03rlM5mJW+cnsYbqN6i+2OJirP6IgF5M1rY/41px1E7mG1AxrBTVNIlWoyF
QBNmxcYT2VqcxiwM7CJnbXPYmpTwV40rU/FqoK+R1eC4bWN4W6J57yavpolDqVd0
tkEukJzntbS8q9s9V+nhKtLfZyNY0eAq8r8qxAzEGJgbYYVhEsCS0JHeBMN3I2jv
EEP5Z5SeUWbBkn2OOPxLL9Sp/FqL9IeBgvLgviqgU2NpHkSGWvNprFvyOaFuMlHJ
FAzSqUNRBkZCMsKIAOHcijQMmK0gwEZckBfwsc4uvnyO/vxu/fwnGKdgol822wNh
+VkHphHrv5qUcrIbbxsNec6uiqPir3D2GFQAWElK74ab558jmKBNRm3V8Gk+Li88
J3WgmHP/EiOGlNqFr5oYjXcqnw3Bccp+laLEfSNNROiCM3v4c4o2hFlhvkfJYeEh
BNEyXx0kR9aE5Nfn6vD0yX7tqwWwU8jBsjnHoRda8ZBUIrbqaU28iJ/LZqgE6mDl
frnlfw7ouecq5r/MOrDLxWo/hMW2VgE4clRhtCzIk/BU/0ZhDoWIwfMjHxLDUTf1
1rqvIc5fcowKe43Mhitg7vNPsYPlPdVuSRtB9IrYUs3rYGUywkVb9ZhRjUTTeDVK
PD6So8RGpsoYZSJpGWEJOxk0KWgCipWPXna1gGJEB1EVr7HyonGyPBEarqpnoBiJ
80KQHieQkYwQkzJ/BF+fZ178H2lWz9mjQQb+fa+tKJq+YkfhEja9g3DJfUlDgmOl
jyU0EfOpPEnRzdatPXgU7/PTNfU85pa8l/oJQPYhqj0zfSnF8l0akV1U3Zh9Efjt
N65FQ7QzxA1eYxsZYGhWzk4us9N354koWK4BkuLFuQUSoLwweHAypniEwNLEsHk2
/jME8B8hju00hRISurRvwhnPQydW8o7UfWg4aVztZUKaosE8/j94MPVsgN4zYMd4
n9sbFed10Htvj2996ROzzkHICE+ooPpO2p+ffaRJ+ddq0I1AyesS4y5FxI0pmc1+
M1x3goPYULAkua7PVkvCa6/1ZjPxUOgpz0I4osZTcSSt6PH9vz/xaaN30d+EdBjX
8OZnmAMPECmL0u8NelpqL1olGB8zHnxs/RCjnZQSoPkoWMUE8EOPZ3VTvd/oMIn/
C+Q9jzEWWIk3/ydq8q7781/AAtD7aHZ0gHnpUFDwfhFP9gsGv70pZhJbPtGzBvwY
A0WVrNjp/a3I14asrvLtOhFkHcDKHkZEBb1YD63/kOhpVRGGBHR9WbOKON6pcWk0
udzL/hRMkh5Ai6BZECp6yQC40LK3bPfTJTmA3vGtjZUKwMN56xBP0jWOPvMwmS06
5j0n1LXic8D989BzTTV8bkWceUxO2Ov6QcmFp92F0cvAuEP/tYZaA25cXiXySLiM
Ptt+Bq2a+Jk6e2vdmcfGkwE3kkMjzT7zTcYxi/WTcKt4dFOgbGpdZKitxLsUHHlk
Uti+H0KDVuy/D9D05CsWhoyQB5ot691jm1fRN12CV2ZXt/s1vGDQYZeYyLdQCDki
R+pm3agsNuCMS5FAPRvYvJ7skwQXrkpXkL2PBLZigwKMXOyZC43e11M8LsZyrbeh
80xkUJTNgdABH2tHL5+cU0pMbyR2HCWpGn4pHxBzbVs/d5bJvaD7NQAeX5sQc/Ea
zW5i4HH+zKRvN+vFx/r+hxzffHTR/Cbm8NUNb4A2xq8VUL5yOxuYIEdTqibfpZl4
Zpt4ACUr95xihCx5aO9yRS14jQXHPnQZeLmK7ccC3SF7cIM4765yXd0xGJpCrEBy
nV5vXF8QrR3v5V5gL0YImOzUCXwZDsmtfFh206wv7zBB5H6Hyqnu/U8cq+d6WrY/
eO3LFeTsfw/LzK9BG1rKQHYlbNCkeeIkSPV+CHcTR5rvXahvsHtuSVTz/zoZsbg2
0wPUgTq+LbH062oIQhbe8WR5pNilRvK79LilYzYG0C6ZGSSb2iXpvCXj52riOmHv
TxAh7xOsndMP3ZmAOmE51Wim3it7hzfnHQhLtw+10ZlklJa+60T0bIERXubFeilM
iCeqse2QcwAg5zOzxUyQWD2dlmxx24Z3x8Q5KxODzsVZL2AkBzwkp08HN2hvRYqz
UIkRJ7J93+So41zninyiWhCpsFuF0un3D99e6et9nssGJNqjjrZFU6juvX1I82q3
rJhGcQ8QfYeMGRqf0D3qpXLFlHUUBLdh/Kmt/8FY/DCHkVgbOxBZHrk7Ly5uoBUJ
JvO5pyZNdrtC0fFZRbB+kj8zKhkWNmZ+rdfH/WlGX9Bq96X0vFwZC8kM+MRVdHSE
1kiqByGSQpwMHoOEI2teLDPuHNtDh8lNdgLGXgHMzyMMprngwQrzg+d6U6CZJKsn
HsX/dfYZn/iieoSIqsxeR8BiURh5BQPz3Jtg+wBzOp1espbRDCnAbV8oUzfU9KOC
zABbLThq48GP4PWI7n1em3eI7lMZwHlX/2uk5r3dnX0tJxd9e3b9K9jMN9bcSAXe
Ub0dR/amMfTxvri5urOywyJWh4M7lpsxOVklM3eKgXWXjvaVlJr58vJ7/FC3Nckf
/UuiNi281BmgE9dCNntgr1p7DDuWKQexJ97wvsHdkS/kWdq1W877fSqgN8z092Oq
S5LIc1c9Xt3hjAKJUSVJfAL0S3LRh0KH6k6se+poAqYiP7QDmN0XqJMAbnmvzr2x
t8HRDtJsvuF4oumCCJLetvpztW1u8GkTEd82FjLyc4NF6esziIYZIbkji4DiTJ24
PIpFT3ubHXVi5W5x7fWpnAMUMAN6mpFW7Xz8QYIt4HnuLwAxxSU7XTZa6xX9Aud0
HNDTXlyiyTiO1wr6wDfts36hi33VaTeSEWeP4qf+xwVX/gQSuf0udO/0uaMeYOGZ
H1gG6810rh0uUNQ7/mxzIOvFEFxcOFAQIl09doh6VTSI8nVlLDjwiKVbDZbB18IQ
g0rCaO0s8eLesp0zPY0qWYiHPySg+1D1wy1F+0sotS4+N3y1te/Aid9VNn278Q+p
bXGfgpZjS+MgmgqQaEoN5ko3SZQrFsKp2Kj9IZaXdtm+Pd9Be8tAbr6hTuJGRdNd
Q0perTKqAsoA5+8gQn9pvf60zLBhlvKWXSnbP3TzrF7C1FF3uJ5EaIn6gBmKfMX9
69/ZBq2evXLSJr47if/c9cSPoO5vDZttOQFARvtgyIXGeBPhzzNicMEyHxTC/P63
IqzPB199M12xcJ8U0qLXD6MXb0NvFHbm/2u3hFmXwc+N6TTubvNRKrHgQ0OE8ap3
tsfdgiGI+EGFYnfEEkGeCfFye2cvkrCg5sHg0g/BfwLnVz0zSjj+edAO0FpOwyDk
2BJOgSwcJB9+YMxB2qE6iraImqa9oVzklcVLVLc1GIx4W4fXlZx9zyp4oAF031Cx
FNQLo5AVdnGQH3JK3jxx97IYGv+7u3H/uImuxCOWSbbdRT0ogPvyxGem+gj4ehZq
eP9/BkK/q6macxC75WRD0p7ufU2IYkVpuw6oxcAVxJfipD/bOJ6p8tC4cP1f4DSQ
y+SJFKH9xK1xusNfmiK9hGiABNdHqapAhzN1mGcKPEt8TxCKyRSeVG+/zEaxS5Q1
3Gy11txd1GQ/Re4NuigLkTJyj4Nh1Vox6ck/4+eIigQLLEIXY7HsKVBSLHt5qTeX
Eq4DLTmxyb2MubBqoU5R8Z5P/MTiECb6Y9yV+bH8LPjlQQp7RzVWbtF7f5wo1Iuq
nhvjusZAy40JljYpXeSGL9EIkyWHsm/yGaK3KBVM3ctpgONI2FPgf97pnYExdESn
AjEsdbffDcroIa1jwT2Pvudfh+zADQTkBly/ypnVtdprsvO2yqmUtKT49mNfKPVM
Ru0u9siRUOMt6wxsvtinnPJcqJy0YBO+tdL7KW0g6DolfFPPSDodvLB2uK90mtke
CWXMa9g9+fLpea8El5Hm99UWufV/NQdOpp7fqCcrNxCyA4gCBVHLcJ/kevoQU5mI
3pkrk/XRYlwcU58Dn/1I0womBl2Xq4+yRw/s/Wd01b3Rze446hI4xOVaFo+KQNgn
+34yoan7AnF4zuXW39b2UG3q+Kh1JzR370lecb7VHYfKX6mXFUDx1LQtbL9P/KfA
324M25DRKS2dAbM4bk423HUH6Y3LugrWMSfeBTUH8DVVhgknUaRzDgIHYquZ9LJ5
BkIMBCKHsJeD7/BXcVcvMaHAp7mY6ExU/HDF34K6pWfly9XNoTKkHOCfNpvgrfCf
U/qLtcsv7yuyvQEhsXgHqS5Y8U7zy9PfkLkUDvASB0YBBO577e6rxAa803O23jW7
BNcqa+lK+2qmEiNfiPJdIkdORMYS5QWG9teR3PLYIYSlO8vT5sCFnDz18+gctxBV
IjBUNV5C8AkqA8gCJUjyF2KyjDSZxEjxzAphAgwm5rXZqDDVM9FZKPMyHPABKxyX
LAePQCtY6FAd8Rrs6fiy8vzPfQlBrOV0nVIEpbKAGeNAYZXc0/0yQDxy4opimUz6
o8ZLOpR4XmYzRED1Bs0oTNOznzX/3k/UJ8WWKtRpNotNBY0JdxoCvqk5NGBplMPo
DXcUcdh5UadhHNN8aa0h5cUU9bWTC0idsdLlFck23yHKQXmcXZhTcpaLyNDdTjCt
A7s9YfuS0ZxOZpysTrhoHdLunyF0H/1aV3Djzp/0hxHG8QDkHUwFQjVg/kYMfHi6
Y4556RB9sQ10TYfO9/eCWcDkDeBGqBWGgmuByQqwn8o6uwo/rp3UyGgRXkbAYtzh
IsgJC9YwLF0QZGDukW27sBoJWR64ZCStRcDa01kCOgPzqLd/eLPDohQW4fuy14r0
npNbiuDGJAoHgXNNyYiFjz4vZuPsk+ZloEHwD/iPbeOFIbPayQw9vNW2lYEfScDA
JiZ4jq79VpqIMl+/lf6s0nxekrtxnzkl9cqmXz+jP0ry+Fh/D0IxGU+5G+MvMVxc
zrjrvscP+BkowVbcRwyuob6krZXL6CjurnPC4XnmFI5OTu/RPxfmrHLnJRHsMFi8
MH37hzncS0Rs2jVDaB/+BkOzifrYbpvdICorYODmzdGHLNyXVg2IY8O7MmpiCsYq
0EvlT310ZrtCgU0aPf7DyshmkakGl4odOcvkb8lIol2ltTyySxOAcdyKohvGeQaz
xVh9jTIzH5Xz+khpRjk2Ryf1lOUEqZCmNDdbB6e+PiWNnxIY/W+dzeqIxkwwAdTL
KyfWTtetM0tfA1tp4XvkuvqaHZmFzGACCvo3C6nt3FUPtbl/59FoNd1vk2U9ol6/
Q3ciMbJ1ElUtiOOhDR4AbP9BdBhrZHgskozf5A4yIhHyYZmCGf1McyLF66FBi278
CY8fCb7pTJadTJI+GX38zfLafjEdMSsqBbHxB5/6JjwGVfv+VravS156TV4nhgd/
PI7spd/Gh6hcuJ5gt/UvWlNog4bECT5I1Uj3vcnyxnrp+VW9sY6o+NLlKgxLcp1F
xKiyXsU82GF4jRXQjJbTV24fZIvacEw110wKfP+WrXzA8Hj+LdPkrbPmkH64Z8fb
mLxvIIdMAe70pffpOECWfatg+7QjVO6camAuUK/hMUavRfcNcq/x/sJvXb0t1xMK
WPUNm/hWoPa5kYyOjXjegsdEmv9Gt1enCwsjkGyxuZIDaWjLPJFLhtff3p0t3AXk
SVmkiXmhjAmvFSenxG5FDFmdppNI9fg1aa0pNw84cFjsRlgGsKd4k+Id0XTfkGNa
+VObm5JIq4WnMgGylrpsbK8TnjPFZu7ApjqOP0gU57dAEcgVtIu0+2TK1C7vnt8Y
wUOwM6lQ3KtHG+Aj06woHjKLl0ubf+RwVEBh23SUqbj2skkSBJx65BaI4pOSKIas
h1PtK1rBPeG5LUnKsXtpAjQwr4ZnjBYzaHrb++lUj8ftHpl+CFTX7xJYd8A6MpnM
cT4/Y9dPyZ/iLJUTsJJjXOg/DsrreFAW8/4uABGjnYiLwr2qJdNtuy99sSUwaHtA
o2IOW9dQqXaN1nE3+Y0kfkrArZGYzV0VHLWRk5Yo5d/5CwwkxuARvs9gR/JsTYaN
13BjwasRcPnz4d/mtLTWuOdV/Ne81IFvijNN/ABD2vEKRuDpCAMx/63yzuGbViZi
/h7IZ5PR0mZxLvy1cqahui/zHND7WpDxwDERohw8CtXRd1CNyjlY9gsQ3+1ywVPM
2WsTIjkFb8U7S4DWlkknn1BfYzd8emRX2mShcbUfBNjS95nV76GGVJ7XYKsn5cNP
LmDiOHeh7iu/Z2i3yARw6oHyX1MDYRsqGmSrRpUY6rZUy79UE+mM9zhx006VsANu
zexapBIeR6fAvc3f1JFzzeS49JhFLsmUSMxld5wsQ1k/UgoyFSItJzPcGmKMuUp6
CxFqfNVr77cszXNyQI3QK+icYisbJcylufds9LCpQTnGdvRPJs5DB+XMpQkUErZH
dYi7rrzaAeDhnYzlmTH4lPAaD9cwGUe812AOQCe84PKLu6LW/bwwRXpjKZulUayw
NDHrhUE51cgY74Sil4EXzTYYTCK6ZRF5CXGkkhn58zsIWj3Jo4+8e9QA0VkmbKmo
cIUKTuL4OkcwhGCsyTof297CNHURcUJXFiUaOFJxfpf7E25Sg4MEBVv/NpkpplN0
7lBqISwxZeFmfnvWQFpthPlRACFYnth0H74aq0kZvSFHxuP0Qoq6H3twIudsVp5B
2MU7LAEWckT5To9i1KC0/Hb58RxMSdQvrqv/2/5NVVEjMbOPTXQntlH8KrcyBX+i
wxTK/yLbTpCN6xQzLwNX2lVkZdir6pBsrLBQ/5PIJibzH4GDu/ki/c+uhHMVKQxS
ZD/WWZV3dJFbsyNpmA5lPiT87zchy7X1GVdn1CELVNZM1xUpp0A6cuvucARr0iLS
HGGzsPsF4s2ymxCnjuONb/orpU14CmYWFp8wQmGgQvzxcqvSvKmpVD+Bf9U8fH9d
JMRM3NU4nmcHohiAkwpCghc8lMaKglfVs/p5G1zU3z1/GhE6JU+FC5V2imUrqm4e
D+maJfVN/XkhMBGUGevpPY7wMVXjxST2OZFjSUKd54bhXvfFlKhjRdpRpFV9Umhj
0mxUuj0Eo8l3pY2HJRZSliZxIppUojAPMERoGYVSORj+tziIkNrS+W0HAayTcPWi
KRpP215IZddsP19vur//V8H6bKM/5GBf7gNUpdgkY8YfkwKvz3YRShgRl+bct9tn
T75RyHyfAqby/kZyp62TJOQy5MviBuKEB+lyNBBL2PUPitJnA8RDMy2jhHMue5WF
y3iu3D0FY/4CEdWJpHJqvBqX58upvAeb/7PJLbo52paep30Wx8HhcOXvaydAbCOQ
eGKFx/nX0TpgSBz3RyT4/TufPTXl8mT4KsAB1vwp27TWMyx7K+brK1aBzS+AvXng
oDgb6/B4MiiBYLKCImI3li7HINBQ5F9+1xwiDZWo+25A+amf6TyGIlO6GM3vcDjJ
QDlbJlLcVFBhN0cwyYK43lNzZgdE2vRexwFbC/+8EXt7dLGXjiViVZErXG058bXI
JJ07WGCRY6zFB/nzYiUG6yccBbyskD/6ggDqjJZ3gIRhrdiTkfq0eJ0Rwn56/5bz
au3lDsg9o0jIaVAdzW3wUHzAbtcBrzeBFYjKyuX6TNxFf5AhdgtvPTgv9qQAtBDR
sZWTsiiYk5Ulfy3RpiDiwihJ4R/Pe6T6Nb/VtXSet7cxBRFBEr7SWAaI1ip1reFl
6xhrjQlvm9X2zzr4LMYWISjeqpxOsMSUs3p9/+ZCLrX2bhQv83uGwjeyGuLytclP
GdiBQ16SOE9lA3Vl5nEOn1pvGq/9bXD67Eoz00w0yQfaBVSfH3URGzr17HusNLXB
Dx/2z8nadrL675F7CC5/AeD++Nle5ZMmwRAtxqNiMB+PBLVOfhByhwmIM1yZ7E/7
tFUNH51LpjZO6tgcuMaaWCuFP/X9S3282tWrKZpHN3bonm7rR9jE06EvD6UTaBdS
lqlb4Vdx3RJXOrzNlT9FRZD3XSp1SGSq/Pr7JHG90idIoOMENUFCUWeFtssqZDak
IQOhvJFKT84kCEKWku6YbqRuL9rrAfGdGCWkFoWiPuWF5gTlRXtb6YPjsvQCdNDN
c4JjUtbIRLm+SexPsdXK5CnGluapCJr75JC19eO0LZGLkYlx8TreFSE83ZRyE5gP
Soer17o4LBVCHmb0fOne9TxiQZj/sFFTOe51KZLIXf5bU3ibTIdbvXGNy8GMJG7Z
h6P64cfz2pAZbWSEHv2vsRvIY4jaqB4tCXtkwPXyHVgMw5JkTRlXFC5aNRZuQlBF
wVjB3w7BPHzFVZve3BwjoBaZLlAvaiau4djRh4bAGVH8+uL6YSR8j8Gowc9HRwRZ
e9sOgtPBQZKhRPcPkJbBYgYluAkCmmELk4UiB8pZO8W8Pulo/T0UmWwGNw261gYA
P35j97I3CqtpHTVV3isigwChDrI0aDwaae05cDepE+0kMYM6/M0JSgVBRVuxkyMw
xWjm7I3DNUX2fQCOn/R2Z4It9cv4iHmsYfFDSygLYkHCBn0kwHETtYQtZ+7w2IK1
bHZxYyoUUy8cqhzBOdgy7/DymBs7YQ6OWS8I7xbv6i1i87aaHQdHgjZBlkzXYMGp
kpOwVlry6voxbMGMDccfVhGyAdzgnkc3x0TpZhMRoEdoqJkTygZXmnNeSbkWnVHT
X2LQ736DoFv1B5eqyQNaZtnWimadinGYBQPpyPsGTnDjBk5XNKBfNXA42fa99/+h
39c2NmuRYOH+4l5L6xlZ0uZARIJYcPfomCOF5iyh+q2zRNOLES4AxkJbMnEmHw9b
KOdPZx965OP9xERdRlbxoqVMwp4PmAL+1VMsxQBEiRpI+TLKmBif7/M9LQLTjegH
KnaKZztLJky+rX/enuT9YG9horw+WFfAjohrXBDevbgj1AUfNPSEjsT268bEGb2m
ZBrdcrJOoyLO/tkYtF8WcuyloB/BR/5YdYpwLFmqibmnI9wkjrQmRlZgiGL0m03j
4zXwYZwmCNKnqOlGECBzm3+vXigMHc2SGjGmDLiQUk+Zi8VrytmFtsweoL6oRhz7
KooALVinTBvN3QYYgdwQt8fM/hUzXfCE37YHG6v1FZPJRxXH/QAEStSt+Dr6nESL
skhQCs1T7OCzh8KOQg+BIic8W5D3cAReaVUiz52laku8iCbnLaofb7B6g9Z1MXAn
E6O2B0gtyyjGZTVBNEhMv5jc0q/IGBp0/AFz0SQh0njuqrVJgcUV4h8rbgsQRFk0
c+Dhrso6SEneN3ZhhDUcgc414zNU3hcfrz9le67j5qj6fNhbVsfqO7fUz9syDzII
083CBfTdsYrNLdfFXS3MSQh9R/nkEJI5GPZAFQt7w9c655zB3IN1PAc6Qr/2vN+l
awpLzvjw5PUkoHSta5A+HCw9xQ74RVS0Eq2gfC0QFj3ayhWrvQUBjwDUGn0dYVAp
R/WefrYC4WU3UZcV6TazqbshDi6PMUwnK/aXc7M791dbSsdmpa08GBv/AGZHULIQ
wiGYG+zDHByiR9oLOiizetrCDEz682ZTtxV2LUkrlPMwgsQPZLSeHFsHNezJ+DH4
yw12v6KnGdDXWgK2MpjXBQ8ArG3s3Bim9bX/WMIoCt+kkINp8qEzrWNtStz+f/x0
wVIHl0Hx6eJ4o09mLGdaKhQ8Wcmv8jWDFlycZWqAFPCcjNlZMBZj+ecP86A1rVoK
nNvQqVwEhI3TAODMJP0AQUpgWGJ0Vs6b/CsuCoCfs6VPyzTr4P0KVb7PI1e6WTiD
6fnH6BgZUddTxx5/xxzKZs3CUTeMmM4N+2h72Oovs/dnPZYfzDlFuEOvRcxW3fHp
hcfGXK3IZBN/DRyk4dEC269EFs4ROyKeRz3IIl05+Qc9lA5fEaRmGd+9wCO55PL7
35He2cZLInS75ILWFvgw0ChOlqgdx9DrCBg4lTxwcbA8kBgRPCH7K5SWbr3A/5BH
Tr4GDipOf3qeqa6PeWYgHwd0LdikZWcF1gAQKAI2DVEzcBV0AqSoxNSsAEIm1OVL
2qk/nZfjXge8rpx3tzJiyLe5aIBZSX5nDnlYTknkEUYJVcFHZQqwHwKEvUmrSTDs
AhoI5jjY1uuHXXOprI4bWCsR1KnHg7yONsyKOrE3I9hNqj5A4BIgtFvgrwDez3Xy
/d1kQ0inJsygvcyuqzevTDmoPGDLmMb8uHQLe1d0E8Qygk32p/fytr06VAPS136T
NJkzv6UiE4PkHkAW7EXe36VHcpAXkktIgrxv4817iiGnHtKzHAPpSi2vp6f51iqU
M+luN49kFWSkqK2nG0282wYNbw4yb6jsuz2KplGsIDWXkaE1T5SVDEkmnOysxZvx
GvK4kg6Y93rrnFT/rQVlLN/AVaLBcM7tG+lAsQ1Bhh8zWxLgQz0/xSbOHuI98vJf
a5GkJyNEpbMaxyYITD4ZD/zLMcNv+bzxegZHdIQIP8xFF71XpJ6s/tDM4VSoYXmG
fP62nhpofQy55rwlaRJJG7cIAklFtutHU9euU3Oja/SbL4fWJwNZhJtBB4t79jq5
5PXzKACSHY0KTRzOYgJQsY3KK8KoJJP3hMJkp+fAjwSgVuHq6XTAqWheEiBvGKdQ
roqgLb7D5DviiMDcNw1W1a4ro++x/cRHnGfeLSRypT0hWeiEZFNoDYyfYsqqfM++
XJCv0SkqveqTbCUS17IQ5A==
`protect END_PROTECTED
