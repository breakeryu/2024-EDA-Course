`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eKchkhAgPF05gZLExabn/Q6t847E9JAed9ZfY95PQgsmtnrIQBCc8VmFIkkwL/2K
0WQvad35r+XpvnRIAX0PGVHErzmF+ZHRJDsffbMscgckNpO4/XaX9+Tn1KVIwiEa
h91F+MQU44+vQS2TrV5agvIh1H2ILrfUlvH+NxEoqlmtzCWzA3FJRydNscntSaaG
K31ooxRjL4e56FwT8STUT1Bu7nzV+EK89o0docPFSAAydTTnJRZO8n8YgCPU/soJ
Np+BjXiz9iC+qHwvVJIYmEBRJU3VsG7ny6NcS496ieEyli+WCCyrLsboC6OWrWiw
sTxODAO7GwiaaMtpIJMlWeoWluSldVh9GHsfs6nZcCwtLiE+/J9Vw9j/mUK/6jdb
3RcjdQmaOxY6JdvhoUh1qpCo2nMTxomSKM48TrYQ6MM38Zw95zLDPUpNb4NZaxAW
YisTgRNLTlJmzGBiHEgzdmsisP5nIn8tVIDa1+mowHmpmBfcRj9QbyvPNa7taAQq
SvtCXAEwXt6O/n7Yk6nJGlV/tS4JU3Y6UKY7rtjozbpa2crtmmKE8ijNsCzIZHvC
40wNTO0uHX3kjy6/P2BemY742RVjUYeBGPB6XbDeNl01Bib5tT6upH/VJEHdq2mV
0bM18yF2rkefS7uiaWgPGl0NnX5780TtO+0Usku4VzdNyUNEm1a/0DXEZyMrfGxZ
WW/YuNBvfmYYZYU1B4DsjyuIxfro9C+lGjK4B5NJS6K1iBDhmtHgLyyg7H1TO+Hq
pmw6lWVHTvS5Q2fl4SInK1qjtkOVbhR4tvssHUrManbHxcBp+nbppjOAVPBQH1DJ
IjXt7H+B7rxvCfnk3zXopWTw7TlbY4zNhCrjkjfNqEXymGUwXKON/nplhOF6mRow
Rrrlr4ytbTowKB+W9ASiUR31z193XKMHpLBEbA46uEZbMkzXYtM99KC6u/cRwm/4
czTRRYJfzhw0iMgSErKxko0TpMg2FaxyvdHv72gVULjaS3AqLwcBCC5sOwc9xmuL
VRpwJTl6prAV9KLDfLxukRDtjzkwg01lPn+3TAP49BHhjhS+uJt5nFm3qWBDq2r9
Q0NF5ABF54nPJf4ofOkLyvc94o+ca+4BnWq3HBniJqI4AK7H41Vq6oeJkNb80YX/
SmnW2scL4wgDHZ8SMPSso0mTdzkyzlLZ3CepfJCvPcCBQrxKIRhQ+PsX3WgsMJra
3AGbwBy4jFjYb9FKmvi9NUZf8ptB6aSjqKfXNtGOFOjMyRz+RQH0fsqo0bST0n4I
IJN0tg/9zGaRXS9ffS9ZDBewXKp3qT9r90lOriuDajVOvBcBaJd3b/71VKbgg1tx
jyCd8IgZKUi+GB9gbGhCyrzCzhxsC9ZEwtwFMdCO+soztf13x1ioJkXbONone2ML
JaN83vvav9Yp/0odb3aBjDVIcYAv84jrlGC2JJsKdOFIow5Cbbgwn9f6d/uLgK2A
Zz7P0O5uYElhSZgu2RM/g3/KpvuA3SdwJUwQcBx1pId+TuPCjA1eWzrrzQ1OePXs
poSwu+8rf4qSBknr4ONOSQnT9RmjaQnAEeNYyB1tk5bUPCAyaALOPDp7+7q1Q2IA
Pcw0rDpniNPbysAUTSSuR9/gWqMHGRSWS1rWX335hhukHRVRlSYtl78JfHC/OzRT
tJs/GMrnKUezSvgv6nC99n/DVs+7DKfCpFyaHqHALP0L0xKs28GunnfCxF3YpZx2
AaEp+CWcXkEY8x5hQGxgvFGt4uyAvUUY36ijl6Yx0jLLITER8xWjIZcijUtSNT0k
/+8H2MMy+D0C0OP8QOXJHMf5UKEFU0sCedwcz+SeRycyUb2mYVc9lferI0p6xaeT
EOaYOcbmXWHN7CopZas47+Xk9gR5XHH2dIG5K1TCjIPZ9UoNRFtI47zq4QdHgCJ1
hGtl3cheIjl/Kl5rk8IL1VM2hEkmcV+Ed4PSfBK8WboZHS5UxP4hq2W5DhmPshdx
9HSJ6gyzBiNcC5P6R6Q0eiQJO9D7sDwg+4+QP13NAmPcb4+DzYKpXANY+KePt824
gCy7IkbQEMvthM33Mo1qkmPw5mVQvNl13U1+zqwFvRS7DcquB0eMWIhC53iWo25s
SZxB6WQH91O+yQ+CBu4uNBE3O3eadJFszfVc8BhptpNBwdK8bQOyuqbgr/xxERRq
N7fBA4ZJMQ/McuLHmbXm0y+t2IDs+VhmTLqas2Jp/zEHNjQmdE7bTgX9A/HkQdN+
/WbCFX0AQvuXfnIk68d8Ua/PURzlixvJNUCmWedowdDocq7bCmCH+p3QLF+fP5gZ
AA1/oBwquloHRv8RcyRvX6vRrG3c/igZXL61FGkf37zIuLBc7gVbyJBSAPQZw4TJ
`protect END_PROTECTED
