`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zh98+r+CbktB3eK/4UGmHGFasr+eYvCnSAHaYI4fWCRJ/csJ6pGdPVYmwqV3TIK4
lS/HJlmgU5SrjgB3dqMPxqvlqay/MuEkUm4F4Gz7HlYWk9Hgq/mwQoU/pPRx0n4l
4WmiQNSmg2mUknfkeRlWZA1ZM3TSap+AlG4Ik3iMlVoFKjGYmNyHly1q1Ete2T+h
i5J0O73HHJUyD57pa+1/sKUHNxy7FpSfZE1lBd9B9vXh5odVEF/0LikSaTZst1jX
jU9bl3WOc+R/FWiDqhonkkJzs7P3OYkwjwmFqO/oKJVNToqmnDQsFBjkbfhvXaHi
oONCKJn9ZWQN3jbElOSD9VhrGRvu7I/rIGykE8fhE9AZNsIYA00ZN0+pbQi7Odmn
4xbNd7eLd30IqliJdpCX14huzCg6fWvVqOf775Hboy5QEm+/5CAl8o849EdYhM4j
`protect END_PROTECTED
