`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1HnkV+2qB8LwgQBD3fGyqiKhY/1oreRH5b8sd6vkV9pJgOGp8/QnWenqwWX0xE7y
X2RhMTKX8QiGIGPTZHzy3Yb6OQzHYrdweCS6CKjjLNlJMcAWh0ITr5kOunYUA5hb
ovBroAt9TFXBuyifLEO1EW6bFCm736hizoeqmIv1jL3Ff0fxs+9m7x9+Eu/4u88s
tkcSMzV6bbwdlty2gg9DM3trkW86RDNY1+nEIjGW/KsBo3ms1jDaqwNu0CcgaN/D
IZGcr0KgyWGJTTR/jGeN6w/t+/4i+cNqpCIIe6NLEN69mCpRbun3mD11KMInDE1o
ake5aLO5o4Jv0/ma7kZlSxXOk+thL3YIyxWYQrTOPumToGNrLHwur+ZljrUenKcn
D/f9kTuIK48rodg6HnQu50dia/ppWUmv/cc7MVA8HJhVNwdExWPI60/C1bJpgz05
uVt5yfPMCl3cKwPl7ZOfmlLNiY0mspJoOhESvo9OmHD63ay+nXj/KGC7vnePUNM8
wWLCazOEzEzfZdyVZuoUGSD3/bVgCl6DKBNnfiYIsdx3s/6/mxvcTpqfKQ7joUVL
esVc3yEE165wRMuPqjyDukHZKOR8LmUIqLiExzVXh8WUpsAouWrhqMFHSMZiB/6+
+e7V42t/9DqGvvFv5mJAbMEAGOWKqXBJGzhJaX+rJwRSar6lwmI661QVGjiARpgU
HRYlcCmfVOUHhHufasvaHn+qxFYRiHRWYFDvCGLzIpALDBtZFIxlkUO/MIolBXgS
NulUe/yRGiDYL43NQ/6r+MJ7UZ/2nQ3v4FQ4MMRdJDdGuBJOETl9XRFIlDvQtr2T
AoY9JqMd+DNbazRpsY6xzUJhrrNY4cXumxFnG/pdeYSgXXLwW702Cs3JLO9hAwLi
QuUML9Z0xtQ4mC4WXdrmigV0/aBkRRi8yvwxvmJ3fL+1Ud0SR7stle1A7ATEIsgw
Ods7z3j6V7RtuvtbQcNS6UFx9EtXhajCnEgPphCBiw7lESUzy8VpsAT0fTqZxhav
oivPlMB5qgIUH9KPBRbUlLk2B1MS/m+Z1BdkggUlpedhKQTZejAFHYPR8DIdeK8F
99mI8+HanopCDpRF9TxUnwgOdhtC2ql5N0MWWNiVlsFNPIEl2SwoLkqoXTDE4LOx
TIh1MI2pA6dZ2ksHeJLq/3jj/HKpqoyIDAyX5aHsRqTwYTAaxwxuy0Uipa869IOb
nJ6QrS0j+lVlq42EVihytfi8LCgD9Pf1xqFSIzDJ5uSRKxapjKQdo1A+DzLZ/srp
3P/ueHGgyP0gkqKwNNNAYMpDdlfkYQJTgqpmJ4QWo6NwjPH/xsQ/JQVUWqfytMWL
+tY7SPfbkunMR6haiYcj1Zfx90ZMu/8D9NEAaEVyw4SrbwFVWgfNYVEczqWD5qRk
TPE7JbDuE84r98ggDbOGOwZ/suBMjuFBlMXe4sg1cMdU+4kJsdTTCNGxLRpyTj23
uKYzzPtMYYLXFUygI0RsM+cU2TkiSNEjxOkyv4bbVofkYbfZ/hwV/32RWuMQA6x5
LV+fxj3sG3njj9wXr9FKZ3TRJgHhkdTT/sxDBjTQrwYO0GRSPWdDi2CXHQkXOuT8
VmG4m1q2fMObeeM0dMrBoery53Y6xZwEbWTqRASOW8aKdUr9SlwCnNGoIj4a+eAx
1yFFkhxaCtyo81x4VvOSRrEEpjDbyDOp3C56uL14g8f0LZbSjdXIjSdx8Z19LhI5
MLLqk+UhHsejQsz4VZsofZN7TOh00VREGNxZKd/nrAO/STVuOpeWvDZx0Isc5thy
DxVFyQeuTkljxFgBp9y3lEfTDHMm1v65yduNtNX69vNHvxMBCAVriLcSSCkI7QDT
brwXFmULTkk8HSkJtr1FQ2EADCE3SeaAHz76ce154oZFza/tlne6sBJ9NbtTZQI3
iQYz2HoCABwi9jM3c+XA+rHQWdbx8mTGoHqUyqLzb7dlEqodr7YcFYHQxoy0IcSc
r2qvVjRcpYdP/8z1MT/0RPdDCLezpTWVKguhZgSPY7kNA86GLmvG7zN4s/WGLZSo
J8tP/t2QR1ecUVdO1l7yqxXto/kNdK054POrkLSRq131OaINwm5zWn7HU4jJbpGI
7qwPDcQv/yT2MmENXH/K6nVYcAIaV3bzbgozUD/9YOhjiZR2QeaozED5Mfsf9+tq
aU7tN0GIy36xheeDU744WugCQ27ugTEeIY5MQKgea/kK3RfMAFFS4jT1ADJKDeJo
VqsKZWpLQ8oaNHCYz5kd/j3Q02QgSsoEXA67d0LIElDETzDSJ87FokZukDY8T87N
r1JMvKBgdFVRTFtJiEcbd8N01S+MmjBJv39zKzqLTOa6kEyO8wT1knABI31un0yI
B5hbKpT5y3aunPrGE1nmzbtqyQSh5o7dauma2m1PVoay7ryCI/wvgGnmPqPJ1LDs
K+Pr1uR+iZVmYvd8+qip4u6QjpGygsV9IGxn9AQLHP+sELlARy06IJKBX/0+0lxM
KvYYW95YjsRa09emDZ5tq5gQsV49zV2sL3J3lbLvGKP4Ty9SzegBSEYm+hUgtU1E
+2ubNOoTWU3HLnDbmR9YtFsVpS81e6yB24XcuFJp5eztsSNWyjf9MP2JG86bPxDC
rySbySfc7ZsuwvC2KDldF6M7oY4ta1fjWMiz1WGVvYr41jlPTj1gqNZfBg3lwxRR
nYmD8XNIHjaaHTgwXbGsMfT8q7UMF7tuYHdH2eor/YrfnkdAgY2J2iiyJJ5EVUEF
yN0BnwpSHZWGZOsDQji/ZBtS/fqLYPsO0+lZ3BjwrtW8H6RY6SlMcgtEgd2bO40z
5pOqg/1rzf8P6diJ90O7OphZhan14AibCF46+oV5eU01FGGeePDGQUMrQUYMejg6
+8hEaN1igXsTVcVFyDt2ePm/nFO551GawyDvik1OFnunZmjo/2v/IoANeCs50zaI
fEgzgRYjBrDx6KGaiqSOlyfL5uLIIckqmyVBOzFU2zviZ/md5ReJWrpF7JuvX2tn
35SxFxbmzuYPc+hYEY5z0Vy5seRoF2b7mlRoztQODS4ZbmhtggfqW/PA2sBn1Mpu
O63G+bL207GeuJnMJOoZpYbMJCWAPA3suq0WK/pksBCed8mcc902nfbt2DEYw4fy
Ii0vBoRDzQCQjxWs10VR+vEUsxW+HcjIyaVFPgTgx/Er24w9y+s/J/U7pqkUuED0
8uVHLCt/kYp1neKDlf0qTIqsSSkBdjzJnE+VeU16Ig3eoreEKmKgT/wVQSm/DjXr
EmY8+uAgYTreEB9cAnwBBcnq9ZvhrcmJpchCrPWZsILHJ46Q08JE9cMZeFhXRuyL
WzHj09u/AipBhUe5d+GakXn8FPpdQcf1e9cPaXBdIXGvnK4z3RLp8ccE2pWoVIRX
7A6ozCm3O4ROnK5WcPsBXXOdJrakhE3H0tSaxB/ABBzYIwWfzRXfVAsk3OpqS5Ss
PCWzyTcJNWVckAH1e3RDUvGdEmp7H6WpZVnZjs2cHUpGU6iFcXQmyPp2J4XY92Wm
cYAQw3VkgL+H/MUtZhXKMnlilJ7DJPZ0TnD538rXHH1wHPpnFjMPpx769LjSL2mv
XTQYeVl0J37d4QH483JtQjX6LkBxS0Rhy0QanspzJ7DmLm9cJxAExpM8thOPpbOI
5FdDkI4vmJvOIZr+ZxXIar1KAqzFClN6W15nN3fQ1tL3/D3rPfkzBtm/q8JEdPAE
aJT5+eEu7SC8/BLdgYY+dL7KLl1kR8JFCnhf06lbeWXlYyK9QZjaMfk/MEaQ1hVV
c1U2Z3rCifm4xme4DqPCPNTvL+5tQNF/oNKyDk846WFw+A8vogmW3akb0h8Xs6/t
UlKLfJrtH9sZ29TZYcKhSCdfbkXboyLi+HzRDFjJzTShoXqDv77OQWUL7RpeC4DB
N5i1ghiS1e+6/Hw7Nvel44pyAmilnlPHodM4LN2ISMJeriNX2u1Zx0CD0D81GFuv
OCAU97+XTOrLn97zU3/zXV8R5aFb5KF/7NPKpiKxPGv5+TyO0q8fkwv6Ual3dbtV
hIbkFCkZD1SZ8aM8NvX+sk7/yt78CMma5zE08HsMvVYmwE+akoebnk316YABUv2L
2VshUkFx9TVOj4KUXL3qrT2q82mCbGpL9zjg+xgHztR+qXttP2ulqz41qOUjjc1A
M5CcXX4lySWTMXWOkxUQA9eU6VTve0df/3IEW98JjQ/c3+boU4XZardohU1wHQkC
EfVB9Q++sqiNAHmyqZGT+FV0GKFXgZL5LZy+0W6UycPsWshuK9uCS2xjiaCxiV/5
OBOE2rdeY77p0itvZGW3+9bShlX29leQnHTffJSB5fjj1RnzAffP1Yt1aAZRzvK/
H3BMHSZUH0Q2JfOPSfoB1ezots18/nFp1jROfViDwmcD4qxB59JTD78jZeN+6g3y
YGpn4fGU1ckj3xMmXeHZWlIkfIKYScFGZDvkvvOABD0aMom0K4AQykkYwdvNfci6
Gzj+kakawYi+pSNKz22m0ga+uALS42UN6+22EvRhEpkfoYkATPwWv2pXhvURAPnF
01saJHACpA82oAqaVJTtcP5V50ZsybWnH6WlMBLgwp6+Qxe5rZdWmT2+c5+xp1Km
`protect END_PROTECTED
