`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fbwDTdz1kboX0+Iz6jfvYctzrqqIlBEcw7MPfQ+ueRJQN1Q2ghX59+wVwbMtkzfH
na3JtDsReJp5MyowpX6lmOrJCuNUxRbxJLO7Mms/OTC4BG64R+e8Oixh3s2GswUE
m5bGCDoLzdBljczY33N6vkS6miwd9hcXcDqUSvfGNf67VMGci7TseS6GKm0MSkY6
/2wLUFaTdSmqJqwERlRXU6RWjJBwtbbu9x0xE48ExC0WD9GtfV/6HcqE+zXj0DIy
kpSuA/jbxWIIfXP2rJA38qleFQZZxPFlc25mnk7ttPmUvrAnZgGHH8XbA7w2l5Lf
uMy5YDuXg//q7Kd2V2kTrnS3467ICFci0ywSyOPgwOHrh03zZiqONSDHoEVJpcS1
ZaLrHcQljaqqsn3uNV6/iQ==
`protect END_PROTECTED
