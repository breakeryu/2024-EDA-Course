`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PdmC6t/aeEdzmFPEgsIg27P17R2GM8FECj2ugGnH2OAtlUlJiq+0jSsvt9U3igW4
CIksXU+Z+3K6vbpp2661rRZVSvQs5douW5uszB8PXN7Azc1lSf+U19qan2MY0wrv
kZXFauoBc8sUq7NSO99+9fU3vFwcnVX/Joh2TztC6eHa+JA5C9zGVljtZlhKch45
Dr3J06frPAup6ZPDbG9WPnPQl4CrHtA57XC0CQ0UjIBJFJk2bwFKH+pC8MkghM5Q
o2Rp7WqEauvEfDB5HJTdhAy8k0rTANnolMNGW4cpEOuejia4leakoptAiApt1QhW
IvoOg+Q8b0yAfLXvLkXzc8pb7MR4UyyB/0fXNoTJQ2HqFP3SvO1XVtKBmcFPiv1g
Pzgk2s8O3s6SfuZys7vq9HhoshGYJI8MG9SWbyJ7khWCT52QMtAWXxQMVKRRcDc+
/yacLX091P6R64z/xKjhsdChX2LHp5r1sGXhiLXR/JXaPGijdshp5uoxc7YxTC25
jETCmEIwSzjrAwoQrFodjxoGwUqJzbGUjcb+5kEsnWhatAloRD79hEHTScouCR8q
QwP3f3hOjR1QfzGnjK+UpadWY6daBuGbsAKOswadPIaW4jtyjhtN7hOupsIAE6QL
3af/sJPm3wt8GYFHLQPTIiAkPWEnQcog8azquC/j0YHEYVZFv010dBk+XqzvFMW4
yBS6hvJqdROTUpiD28a+hJKsV6l/nfNUSnN6bjqpF58raT3rPwbydxYyGsW53cku
ehzF45Gf5KOQcR8QmgcxQYjEs6dUCFyd1K+Sie6WM/8oE+IpkR0iPT5kiBAoMfeP
4ELM6VT1RCreYYbGUNe4d0zhVzuiSo+99m+MyKHmGB9synJPUO529Zne7Fo7m7mY
9fu8wEiDp74PaG6DSt54HNIAyychRYp6JCtMxdTj17JJ/H9Ii/8Sx6UF6Du+onYV
flKLGYJ8SWNPMnhjuhV3V6aQjt+6GEkk5flGjm8L/da+jvjUi5JOlC6C5TsBd2Uv
IGo69OizeBJcx+F4vPVMKTveMfJaAuvSvc3/dh5KKJTiDOMgDsguYX4SMrMqzo+C
UnSfbKG1DyzyxnHtwQJ9u2tXqkfdth8r6aq9vzVhs6wH5VfiN9wzILKEjDYVospW
N2O0Rdn5XW7KsAB1zlVZUQoQ6tUXUW/uctmCjTlieF4s/1+CydRlWssnWp3OFMzB
ZZ36a/ru/VytoiRzA+xsC/FyqVcG3LIpIPF0k6EjxF3vKLa1LtctwdXtHxSSqMcw
wCB+AUwIJeTlBLI/FWzoFKcx6THKQT20C0yBRfQbulZUtmezE1BgCqoHmkgsmDZw
JqK8li6JzSEsjTjCeW8xmEo7Njq9tTev5I+QVMdGoCmh9tUbUmaRH0EE153YqKPJ
4W825Sxg2zJJ4H2hmV7/b/Ri9YHhg5mPVcxtytTu88wnGyuIbaJuVj2zZKZscnCr
nqLkM9N+9OCePklrR9HvdTv3dAhWYu5YVA7lyj9fQJJ4j40cl/uiZrTJmkqet4BR
pHhldkuSa5EE0xXHe5D9wego29cPVKD060+Km/CgnX5aDQ9GodKAxf0WgXMcPaxZ
0Fy9x03+JIIXmRvfa0sz4qBswjVqv7h3yM3TKorEvg5nxuzBoZY96ZlRZjmu3RAs
5Er7WV4TSLwS8lH8Uorw18MuoKDGc0XgToPOciivMrl7wiqPVSOSNmzwWeALYqWj
0gYarjnWm894xi9FpS7S/Yw4Q5AviJA37pEchEYtC2N6S5wy+zuAeKOCHQh+7xpk
dFIo0nxAFJbKHIQbxxsDfamfMJfeE/GZw9EWNO4d3Fha48l/7FTfsQc9nJYfHys3
IbrfKLvH8cDMVoAr65J5rCWOmvoe0v3ZBJpQcwOe4b4Tf9KXJntvv2ZWG74IOYKM
SbDBBLNnjpjSRoLQqBWnD8tnqEwpE/VtYMtW89Lqn5RsKu/5KGNVkh8kM3fg3y7c
Uh/FMuLF9kHeQsuFN6OlVp5J5Y7tbjEc3VQsQNcezprPLAIeCYRLaByfTpclsOeT
sef6UWzou56E0tkbvW7Q5yxp3vOdHtuNqWubatredRPB3Pf1ZWiF2NogdMicaRVK
Es8GlPJ1n0PetH2B7MLUlTqxuxtZyfwPAM93in1vME5ry1TdpjaW8xNbMljDqKGK
D18VUXzYJVjn6ZYoOKI4PYVKx0UmH3reBATY/hux1ZaIfC1nR3xhel+sZCQIhow0
pJhYJl0kKXe8jHikMUnkPsojKldHnSfN7p7E/l00yKq3byDvy21nbzjeQDbg166n
ubP17JEZqJIoeHiyd1af4MHf2QdOC51dDa6gPqR+TMz5OfQSM5dx+dipX4KDgzkC
oe/KkTgwdvbPBKAWHEM6HATJk10vcp+ManiCMltIXNzmcgqoy3JtHYiLb65pYnLL
Hv+j9SmsLULZVfj+YMqukVMEeGD2lP4Fk7eBYKNAtkeGAokGWDPmrGbP4MObUbtc
VFRjNbh/v3WkBCBBYnzjvkAMuS0q30iEh4tUTlGzmXLiMILnaLJmDVsbuBJ/4bOy
h7zeQVVcZ0B+t36kc/VSeA903tfS/GF3VeG4MR9S81MJnFDZrrYhVoeMzAdzDmFl
wq9sJSsx9pcw13HHFPiM4wE4k4x9h3rA8qOlEYLhUn3J8GarMjdwUiSNis8fNMyP
3psBSDL6Z4GPwDDqgOzXF78KzQagAGiVdVQG6E6ns7VrAIkdb5QacKSVj/dc8jDp
6hAmqtyH7GytBmU/JxwZVKoyoXRtRZ3u5z8uVWRGjwQ0/c1fozXvZBimhKt2IOsk
5O4A9U6s69mDhVzcbQVoC42fsSKthEibFLPdrXWN30MXhZ5OU5vKaiMewg6zwjcb
7CvBMvPcipCjYHhowh8bhmwKKOYClazdTEtCX+JLK3HU5+n8hZTITYl/EFSjnCMA
CmgqupUjZvVQ49Ey3goYbSQ5PmjQ0nERdFrA6jKsnr6ZJ31Ek3QDeqauLyGHJSRy
MUKa6Z6gZbhyQyZ4Jdnbg4QA3/BawytnISrJe98CS9EciwATj2PdYO1hVjSTTiE2
to4FCef3h0EezSPLBpjG2QLQi5MqU+v80phzLS4jWFeWw+vRvT58SFOSSMbQyprj
OViSuXEybvKcrwrlM36/DJ9YAQZM5brtDVx1kDwQwit9AW6IQAjRWuqaqKUBaQea
7mGTYCmByVmqpJlM2IbmiV20XTqHKoZgwE7AG0y7fcuIh3AzH0wHOOn1PGooqrVt
26spBwza8+tsumsHkE+TkTEHWlOB8+CRw7zzOKPO7jekLxhC6vlJwBPs/azpEKtd
Md3uNKkBCqjq66yf3jMelJhFA0Yf4CeoHRo7K7ht6fqza0uw4U5qyfZpaDxTrq20
Lhl/zX5q5r+BoD3h/J3hS71LV5DhV/6QhnvUhf3j25x/rdQsyFzjqLTIG2IuOkHl
fxDsD8zs03yfMX9/JEGASVGRphY02B7PIYj2Myt5R8/NVIWpuf6u2NVTJ3oR98PT
owFn2Mc4SLH+2qMzA407rE8RiSKcTCv9MfsI1m/17KYAy4r+A6hfnULqfr1vyGM4
KuK93DI8x4xkpNoS4n3dTAv7rUZuUnsmqoBwVT9CI7Lg4T/2bIfamULlETBpQoPZ
LL9QPSzFPCaWV4/HWuZx0m8qtR386O3Qi4AGDjXIC3X5RvfzzCnvFr6AcllVj8vt
Tbp9SKN8fWqwrWBmHw/iCgFzrEI6aSDxy8U7jFy9WVv032DbhWgkd2JgIaslHPGS
36AFiyiOyUgIfTWGjXRCNCJUul+CmmweEavCIrEkIjg1yFkD+erOIgY5L4Iyp+95
qJ4VYpOXKk50pVuUDHO5qJOd3EbCX6hSxsh5V7XSzhl77LvATUxnkSlocyHB+qTm
heR6og2av7SrSABG9deSQy+XYTPjs6HaA20AD9GqnH+Y5u06k0yoA2/So7/K3kCx
wXJOd+QM5ZMn1AZcvz2R5JLEgbfpMmBBJ5du4EuzIjNqlKnqT64Y+9QTkkh5ohaz
xN3wF6rG1b03pL3NfyEAhw3nuKXsPSRpmLbKqFkgrywTAuKuybBlqs08Du/2dEhN
BW2NgWsyQGBVgkWm5u9rcaDls3S+k5PW4PZu7GjVmzgT/RbTwIBIeIWFPTBDiHFH
e3eXYxp6TrJTg5RBDcvW2CiOlX2naueMEDDfqHN4LtVsJQ7IfqhEqYwWDUDWIOmx
rn5my6fyuWrYDOp+JfgxrhMOPq2F/+0M60AwVk5wM0wympVCDl8sF48kLg9VO8mG
3vVHgQWESXN2tnlxDVm5+/0tvE+slP78yx2bkPP3j6GAxq3eBzE2irYZ8vUGEkd0
T/spPdq+COvF2fMbIrhd/LXW5BWC7nbl27bG5SG8Ds4HNLerLxN/DAjSESa+q6Iu
tq0VJOef9a90Dw6Ok9OoRrpQF1lZXr0sQqEh6ZSQm9Tsx3mYJf+zXVj0Exrgbe8p
4WbAhdvxNO/80EtKwtxhRLj8ZhAiNe1iLTLFKOSHWuBVte32jnII57bqiW4sFjrH
2UH2PGQR0zzqAUF9I4uaW8s27PFnbG3TRk7Grpp9wJ69Cydg2DEYzI4HZhzMrlob
OQAQKWEXwEKUrQkKN/0YlcdvdlLz4kmxQMlzigDLoirGPF4bErjOQVOJTHt5O5s9
kzy8s4asPabpPG+QqtsW3FthY2XqxyfcmFX28jmFbnVgwuOGYGrQhyNlJ0P0n6IW
84O5I/q0y1rxLqNivVQWNYh2u9Vz1YmUX/LbPnDTnAy2HITmLkzuY815dXD6cf+L
OEs6c4p/zypyAAPZ2BCTujMB0BBobxhKbe6Rr/dHqCUQhNh9Vt1SC7/89AGA2KR6
9/qzj0ZS7fxmEAESCtVgkL9p4V42/21WzgpCGwvpkXXnSAUIFwICboy8N/JgOxKq
nKQzbjKAsaKHUZFCPW0mWFQudtNnwXvl3CVw9eJuLMAKdrUzschynnTaq5XhwUJi
O/f+n0mcMrbxmQxRnhS79CeOW+DPHsNrXRT2X+soq7vlVbWs+PCBD1T27WKvKB6k
iFXeGDdvhCqzDuCAyoDhgsLuQDC5CAxD5npl3ppP951C9MYLxrQiALPg4ZJctr4E
JOhcZe5GoFKhCC4N3xqqvO+xvyq1JDUUrGsaAPlXjz/BbFmvDuZ6DYzQUd44vE30
Frz6WEvSVXgUh4Q7jxQHLBM34OSxVWrZV4QUfUcFU08r4vYD0Z4dDcRIztwjQ2KZ
FapyJDqQ9w9MJmtvusbDT6nUv62UXwXMoWnRcMz5+MVDn+HJqnHk/eJBowi1ISNX
qV3LPlwRd+A3haiUp68Wl4PZb5xRmVxQtflaXlYk9yYQzlkZD+5p0+bhKWk5+X51
GwPst/1paC2kStN7Q+nnXKwC7XFYqDwkzzHuT8pdEPyc4Nf/hmA0wKSfOGVdRueE
eQ3kzKP3yxwOTjXbiXvOa2HxvZj9qNZQyXSh/aMf9CZuEPV3IIgqAokglJ6k1KHc
hJdF3OgkLwqdNeZzT5cMkxzvzHxOcgo0CwFg6Ui8ukVDpTUN5cjx2MX7neaAq6TN
a6AY29CKIwvdOEQx8hxef3NeSH3s9eTXyexYoSniV884RWWJQoD/pOe+2elAHcGV
Pn8Qlyenc4e6kt2GNG97T1i6U4cxpIL8f4F7jdS8diDWMTxi7HmDFvOdvPS7Chpd
z5l9p7fMXD649VQ8n+uOjWeBqDsJr1UERrDNBc2D3P45s1sB8YsT3oRwJzD9Lfi7
RpRN0HTZucJAgcpjPFHcYn6ePir7/yRhMCk0kagjo+LvTB9bMc58HCzv+HzKiVBp
VaYtOP9nJ0R4bObhHy9I4g7tjmZdH+MbPDmULuW4gY4U+9PLtRIT+kQRI2fNfWIZ
vHhN/ij8QE9ieHnZM1LvinSPyf5hjr967VppCdMCt4bRgWdL8BPCIUN1DTWmXs8l
ulafGOI+SGQsatF7zho06MznQi1h1bdvrqO9o5YPoag9uc6BVil5QhvDiYfOQSmr
DI2pjhat3jQb1mEcqmkT+BajYQPBaOtGB3GqTPKLGGnQiX24qVzXfWWK5nR+zDC0
IIKo5nX1J5ZotqP71SiqI+79Iq8wEF8gcQGcm69k9AWHtK3rRxdoNGZVGoCbkFsB
PXF3lo6ZasmoSaBfc4xZRJFYQMlu6ykBUGs2gqahYJ5/9+EkLulGCW0NNqeCdmWp
tKtQRBBYQywLyFF1pHCwYZhKKlgpMKsI6jwrqnjxYX9DaaRx8K2kf6xInm8wZ94w
zsAGJKjuVuta7R3Gk9Z8Ww1+7oe6F4wGUk0Vjdqk25z6DWe/9VEuGoFH8tDtlewn
12eRkl16MucFHpbpM6vdTOCfGyC8ISBN1ohQFHApmUZ8JAMJNq3SF4WKNODW/vi6
ZsQ+CrD8ShUigvF58h7aqFTXDu5N5LGJTYy5TgG79YAiRfOWEwfbTPnduj9oSFtl
e0lQ/OTuuUI7Rw3AZUC0W3w3gCh1drR6ejBZj5+jcUoE7BuwvAwQuHI+rDT5CH+I
dY5j2lfFWh1rE/SR9taJmFYv24smVneR4wC26Kg6XQ/jmYMKgy4SYikp7jLmspDB
hLMt31ZMV4O9qWrzn5o4ul3O2XewGkLiBv8xNcASEAfLfrEOeUxvrMtiEzqkfQEH
AWdt7ZOCy7FiGhXzp0Gq3CBW3+6Ruud+GWeuq4RF4xRLmsSjLhCQJRuMC/f78Nj1
UKeE/ARrLaDs3cjH/+Z9N3yzVeE0o/V931f6jD5EQs1u2hzENg3dmP7ECV3IzkjU
Z+LV4aZKGMd0qRgQePay4OEevh9B5MLgRLIJx6xJb1ycK/O2pYeGNNnz3SFGFfgo
5BaoPAQrTpA/cyC2YafgD4jDnQBpKRzQuW0MYS6B/LfxwVs6YUgPOm0tFYtIDhX1
nQU7cbxOEreP33UlM8IPJo2/sZK3Z1xzeCrrw1/RAJQG/U39R1+/WgtW29jKr65m
gFxy7tgAz86lR6Yrq++xhXURrItz+Ra7kiuofaqhMAebq3MtEjftJMJmuoKiwLGi
Vj4Edz9xOf7SekdGOZCgTu0Y+Qsl4ZIrcaaFH29qSLlXO2r9rV1dOuPVlI4qYVS1
hq/krYGRpsjnaeDh1/kblFNjJNCPIQhp6aSZzioFYx4Hbh+goK+RQsMUDuAg95MS
pBeW0Ci1ZHS9WAa9ktO25DR/qjRxFXmdf9AiQs+95GCEUi0ElFIx3Jzgc7RnPoeq
j9vA6PD9ornJpd7tIXlrGTlWSuQkRcRM9KXMaD1Okw45iEgiL86D5biDMXpyMUuU
WNxsUOMQqQa3NCUl04hu2dLMt4K88p2Rp4VdODb0ZkO0ZxvgMSXeXgEH97zj0cbT
FP8B/9o9ekfRJx6MDRX35/ursvZzmFiJQb0OdKwIo/Fs0MmymJnvchQpqgi8dysI
0jWRWkrke1BsF9huKJWayXRbvCsxgKhBZcTR799JpGCdxumBjrE596y0ze04XSJI
dcPT/jYGCnWZ973/My+cK4Q5M2kKJidlt3fqcpmEnVzNAVAXT5VSPcJHSuPBBUqU
L3090BKI1vYLydfdCCWSS0ovexlp8G3slGQI+UdTosKejIV9Dwd0+JWJaCmikQ3b
QTvkUu5iZI/5ZK5/NrcnjhDzoJT8KcAJ0Rrs1CkZ7r02XDvqgwqNjSugtG8omG2c
qnm3XHOtEEr7JXD6kms40PvOxoA1IF+k/erfGQByxZRxpPIECby82WNshiVbJRM4
DW9lQ28SHgOIX2f7Q6/fqzqjJPeGecvoriKQdNo0L7qTecUM4uTCgSmRYim5nKCb
9pBQ9aaqJu/RZ7SNk6XmtrXRyS9cdNHE9plmN6wZbdflXJCMLyWLAT6iljTjcXI6
utlfPELAWXWzdAypbF9tEBb+QashMprnJozJo2z7cY1pmaFs5ckhBBHkEa/72dRT
799/Q7FqgO2Hv07CLpjKtMW28hm92iWX+fHkWzdrZzoFiyUrI7anHgKE1P5yZcMr
HbLo2l54hv04lkHKKjcW73kqakr+Pj7pB2Pg5vZ9csCryYoqmIIyfH847VqyEa0x
xQC59ajhzK5P+j1fJwUIQCiycND05Q/OJ+YOaH2D7+S3oXPDFUadcGTWowjSnT9P
Sb8fYZwTLmnxyILshqjiXwGcmcmoOGUdTV0vSlOZr99+JFqg8lVyy80Iz+ogGJ0Z
wO/32A3vtR/faGp8S55hrX8+wCWfVhwEZPZHl5oU9dIDiCfigHVI2SATCNC8fXGw
/pQYhWMO3XbsSTSnioJY1X4SJ7le9wPfba4Ard4m7+IisM4g+Ou3hx+Y0VuaWiDe
cNUSlXCteSPGXS2+QLPvXzg1C/kXcyraBDYWgiIPvH71zSNLIo+bhfBGxI/gTjhp
cTjRsHw1vn1HjY9ykQXb+HgPqJDOXFfmFGVtccmraRffsJXe+KWIijdyEncNXOc7
I+kBb+LMnUO6NVo9j2dY1gl0TiGrfKJfqvL+EbaOMkq0LmsEIXuYu3sf6+sfKvVt
T7DRAtUFlg1KSkfSPtwSYHYg3RNrdhRYLpEKGKP4NW3Kc8BvP6KRg4Mq92XS0Aat
NxqbM7EVr7KRyrwUxaVxDrQ/szijhCTN5zjiNZ9pjybKX4imOaoAYd7JmcCiftL1
/wFnSh23XvdiPNRxrS+fXXnIsHNxPH5B09LKavaShz5yZiM8yd0IsisP0dGQwHEy
MoVOcoHvf7RUKEe8pak+ltXfALSR/j3BEQeKDYzvsxOpUAYgjlX4H3JKoiPmXE3h
8LP16eyBYe3mDObS+iR2F2PRs0ZaEF8ZN8d51ozQ2akpSaBOaziJzf1QL0kINCJ0
vr2O8in6TQ+a7t5fQTBA+gaXuPPjtRfquF+9PyQafkDEAKszzKuihxXeOSbxUaJR
xwcKAzVaXCWBaq32Y+BWBPvUf16uYaDEc6rzX8BLhgVoVQA3eGabxfjlMAAPocNl
iToONAM2HVgvm6OlWFGUmpgt3cfFR1wa0n6Pc6hqlv46tbfoTRX4Trf81jg6S8k7
/6Y/fhO+/Y2H0kg805mTmmXACo4rJ58Kwt/wsyvoQ8BY45SBs3RLoMG0VJUwDTud
L0KjjKvoPhyl0PCfHXyQFxgCDYKH1RDuwV6hmun9WXKPp9b6ULXQEPOqyAX2/Y/Q
u4bT3tlW/HFlbQ3+TrChuRnUu+KVyRYnGJvdtn3+w9sssG9ywBnyb8zecc3zzdDd
OFRaZVaCz2TfaS8Tweo3r/BmwDaNvEYaYAokHpGSDFxSo5fQ7NNqBKyC+6OUOPGL
NekZv9+cDgrxAV9R9D3yZ2PB/B829cW3lqdt3oEj0Iw3ENA/UdXYSb2oGJrfN0/A
WyLYmgy5TtjT6OzDk23WOgSNJczLa+0+cAde4XXiDJMr3rvF7xRuEpwBV7+iObwd
5b3duM3CwEiI/lFs+VLPeE4e7YMISJyQBehGXAJxwc43mGFLlNWHijYl876RczAB
6siZGzgWF8S5CNb0A7PF+U8SpnMDpYCzEq97hwAvdTKjQxT2SE0I2ZquesoLyHV8
CO5Hp+dS9KY95HA7WpQ/katxvEs0xmHRlIzT3KWQ9MwAm21Ptz8sISljC+HOhde6
t1C+hPyoynjJDljDO8Bv55IWyn2mWm7gDSFeBjK3APLRzuTNkuUtTanlNmhtgkf1
SSCHL8RmN8mRok2Tlo/Z+mji7jg7zB/yFK1T8MftvFr6lrwtdWQuz6P2WSV7U8xt
qpf7Q8K7De860mHqxv9dcZlJXeXOlkARodM3Onfq2Ai1+YN03Gp57PL3n0UG5q8T
QMouuDdrjgYRMz4foWOuQgVtPM2zv/2PawK6OBGroUzj3X+NlnzUUDZEvu051OM4
eEJQDqp13+7ycvtdIrEOWung5YqXtCtMsBSL07Yo8FvBCUWhXhul+dPN/6o/94ES
X8bYjZSxlMNF0Gq1/vzBSzizdJ8gWDEpc67zCh2q5sz0yBtVcIB6NLlxlmoLghvr
WPhGk2bKur5t21HiDKbPpwxcOWlu84UwO9wzJcti92OA5hF1XQX2Ob7Sot1DKCPp
HqcaCMncg4x6uA7nyLTKzu8WQ8P2li5GCVsE6vAHD005Popra80z0SO4BE8hCk6v
DyG7BEC6+a4lDD5eNj73YpWjk912GQWwyXWha81zuD+smiJT0TUZLljlMQ+NAj9e
ZDKVjGbn3L3xiZznKECNsKcy5sOWWjhgRZBvX3B1y3fegTkfL0MRAaRkm/kXx+bW
jwlAnzj+Hc7p2KKSHX7ClSBoH4N1dP/vuh3+/oagGHMm9qPucYV3pSJFjfZOqaw7
6Tm+Gbusieu0NLYEscYpYYN/rMlTDf4Z+nWZP3caD3tJHMezT61KQs4mp8T7Nbwy
OQCneTL8o59ID3n1Q+ld76TEwtxsS69KLrQBXskkIsa9EwQsSWBR5Xp0BtSbn8xo
UgA2SZFYhLVoBR5bKlhPj6CV5AbqXFLTia91tYEa9XMfL5g3h8sXu0gRssQiUg3E
ESt2hcuuA/lGTKtT8InwdYpjwpO5VZzWtrq0GXzuZcQ92ys5SdQ9MbsGIwIgR4G2
4k07JoWBSSvcx9a9rPUuZ6yNsxEAjqsYaDkx6XMfInXn7j2pDE5W/Lz3qxMnzE38
/UX7PBc56i1nLaFq5NywGYOQawfOEukxPZF4vIcE/kIK2kaCCs+Vi7sbQ/3TdssN
VvxcNHVpTDMkTye51lSfdCdOzBkFumI6ivqvurRsC6CK7yJomLFbBCo9IW3UYVeW
wF+nKQmSVsYqzWsMaqv19RuHhCfm7AjiJUzYfUNLoNmHAi552iN1pFxVTwMakVic
PBaRpo+nNFuRzE2v9Q/A/vmOgArj/7H3gGYZVxuSm49P2cP7Dx0X1rim87cA8H2M
huqDCt2tzbZZj82hnu9tbmbKYF0JlTM0Zbq+QBNqSNUOjVaF0sxc0DPP8uAiGjLi
GgeORXuAhmyXY9lgsrMDkVprpo1aNddgIdcvaGbjMLaJOpnvrYEoEcb+2fqSwTES
FV0Rmajbfq2i+qWrnugpglxi8ml6oA8O53G6JIA3iSQG9yNMgcJzbSYE+kzN3QXN
nmAWPRX7wv0+2S/igcu3j2XupakNYRJUY3ZUnbiJo93oywKI1AZ/KvvYV7wPttlh
QgNGT7kykFPI9/0Scm483n7waow3N1z3twIssM8edsEGb7zVcrjjPdyLV5tlQe3l
LVUHp7boPbLvgJXXFfD+UKXRN8dKxAx16ybswh6iluvbTRFP9sTGCyruhO7JK8ik
BKQO4ylTJZab4NuYAP0OvaA69KmejgMYDHDig57KnI9NPiApDjUgzY52eke6fMjg
hzaZ6ugtM+0tKTBhwRtxf56vU/VAtqNCbSY5U77KkRo8RzG0TZmteoPLA65p9E3w
8hq7I2iKqirmVC4TVjHnTCG7h42Cp089LthatCuF1feMvCuRIn7z9eV+hsdkg+Xy
Qir3IP2q9ayElWwJ7yWpi+PmMe/posL8AD6GIfOGqX4M2sd6aJBI6e1tuoFLfe1y
hFVCcfP8vUcc+SGkooLpYXn4woSagO6OIuFTxRVdFjfT8r76GtBV/WtfFOROeGBy
9Pj8uhnjn5jITTZTsJgiU0620kAQO5e576vDhlF7R0cPF9GBSywDJVQBel2BgqRo
TN5MoeW9tFkoCtQoCK/fbFswzM4JEZ2VYPNoNgdIgghzulGLi1Pgc3Yfg+Qe9j3x
wmiK+U5Efl+zfpxzaUoVrOpapwhjwpsYjblwJvSClPKRT7wVlT3D8V9GkU1aJ/dx
t+vJyZLnxO1dbmEA0CON7UmdRWwAY3MsYR41q7szXBsCkZ6Sv6U69wzQQP4d50N1
Ymrwd3tI4u8DnkPHVM1fIcEfh49TjJKIa8z4DOHUg5xgoietO88c9B2RwK6dMGCd
IBtQBb2VWQSmONm9ngGGi9qTXuKN1BbtE0SX7nId2vqVUhyrdfuuUgSzEwbyF6PL
AzbCKbMpUMlq7LVgASMk+nkvaU9SGgfC8I9BM5pS1swJypu0kXkU82pl5FQ0QvNO
kbctYfQUveOHF2C209UAG8PsaGaJxBxvdiWmYyH5y0eslarw07mdV24vWQDLqUjs
0bdHJMLdv5PyQ5oUCc3KHXPs/aHNyNTu/aBpb5dt+WcnGklOo2jsc/wIn6ig+NS1
vDi7OwPMWurrXwFdMGwobJ0SaL3iUk5YO+DnEQLnKq6D0VEoo4MYvdadqnfjQ25b
7PLtqvoNX0OFMl/3ljkh7FJgjCE7DgZ+CGMb2Urol6H8uNnz3+ErMdfFcsdxsq6P
yuWDPJedQX4fNnQ+Z/agRCzHhVbfl17m0hvgCbE8mVAEl8FULp69y+avQ2DONyV6
8Q4PxXP7jKGFo0SxrCA8rUjI2/FoBMmNJzZDUjEpYM2W4GzxAt0KHWnhFRlMfKP3
4PVGcPHoouLVfs2BnJ3rlp276M6xtwAXpEPvgy8AWF4+eBTQXRaz7/bBdTmpaRmk
JW2Ny8q8OJDYFZOJrSu+8fzcPLo/kYafhM/DxMQyXmgVRSYnPHjAujgSqpWNFdIS
Nb4RgR/Ql6c4htUlHXK7x1EM2FCbfPkNTI/qyU3nv0qkXHR+ggHEZYWVuRwzf5ms
zp9OU4zPkR1aXFOMkXgMYAlqaC1RspEL5A7OQ/RMtdsdeps556nqOwhgUG1d34c+
ui3i065PTP0a+YKIl2bExvs7/47PYiGGIAmjqJfpu+OEoXJv5o7fJFvBN8I2SF+V
dc1UhCSqkyY+EKeWOrSNx8lr0H38eVH+fmiWZsY5LX+cQxbBWCt3N1Hibg4Ir6QF
4ZxaVMcfbd/GQ/Ys3OyCBKI/YLM33wln7WTpQ5ucFR1G2bzW9qTHzq8cfng3OE0Z
+ifImkc6gzmpFQmTcXZWrrJgShwm17K+32OppXM0tAlFk6XBxdohbmKcWu/pMgFU
82nRPCS/6CF7t5+JrGpl8StninmHSMLes+p2xLRPlyUDLWV5vGf29JLgBtQzTXoD
JKDJkl0jzMCq2ZnS0waqaJIbLxK0qV6M9PowjNRYMvbyBa6xCREtzIwyfqmGXyVj
RpfT/sIh0by/nP963fpZTdMOnsuu2bP0xYsp4yVZOeNOO3tD8/44eBugzO3b+JPc
KoIjk8LpToqyNHEO4lc3FdmPGtmixlf9j7bxTnm5bC1dqYqlv1Aio6amLFwU/LuF
wq7SnD0vzzfvsAEmi5dIdx2NJrvYFZ4GcTxCNbxtFzMWmxCqHEXeLxwWBA+GNzVr
uO9GT5laZbJrKrk5xXxXe7Wc/F0hP8QixYNAWmwNp5DRqF7EappKnnBB+in1FWlP
V/umzMHgXncQClb5m8hNhw==
`protect END_PROTECTED
