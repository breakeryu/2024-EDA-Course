`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FI8g+uIC+OXPzasVWPHsxnOb3JWwTggp2yRTBq9uTsnJeMtq7rrKFzq1xCSZB4ow
o04y/MhbTT3oIv1lzd0tX7Fg8mHkm3kC6daBDBIO93Cdj+jMqwyrg/vJSt+/EBXl
ZPv/VqHqX5nFWl5ey6zaPiZrNCMxqGtrlM3rnOpXUxMHLD7FSQ/PQg3zeIvewF1k
BUivZHkXiXAibXikY7o2KF2vrUnyH7MDanVYO5kGIvfDJrdWDVZDIBA+vJFJvb1j
pPqSEsqFiY9avnObr+SWjOsJK/5JkHlKrPLiauXepkSNBNtLza6aRgN1oUkFD3G4
JPcIybyoLLyvtE6a1Vq1aVFu1mu8ibwAzaShIIsKqrE0sFeq/pPy8wgLbquCNjM5
cl0Ioa4I/osXZI7AJS2xlJTupT/ncCs+RhBsgCgacyhiVNc+/SegRSzUwf2zrwjk
56bx9sF613pzVNVMGtgctRvOv0uHv0nLHV8/WOPwr5Xh3aruubQih3cQvugBGlV4
YLoBRulpbOnzCuqcKEQS87YvgkLFm7YhySq6b+jO+H07/yynB/Hry/48SqJR1WJS
51rWr5gTpeAuNq8mjfP9gpH9BCud59klhv/tuh0+dp8DCQt0Dr/CyRJHmtIjz9pP
eb3BeVs8WvKeF+lxpUNMk5mCFet97cENnZdBpJiNPq5Mk1eiDX9DJczKRXo/0Zdx
UVFEBGFtnKfNLENLe6cEglQwGCTB6PyDecWhW2AxoCgNIa0Pn4iEBM84qMNhzghI
0/O2dZUEXS7QjsbjmPunAF9osxN+FSQfwHZlGUFd/n8tlYzM6ZvqCiOdKm+BLvSp
8amDzZvdYPq1fhzEG6VQubEH4y9H+mUeduSi7njLyKHMctPN8/752HrfGtSJiCu3
nqyZYnlKC3rmTHUOYz8pL+Hx6+tD7kfoC0bY3bOZYEdRE8m5L3CjeR8xCXaWnnST
3qHxx43ajPOlCYAvQ8r/JTZqWODTtb9AkJ3mFwGiELsmtP8xCeywsiGbvp7GJD6g
9Skfs5ei+d8jKlaT4JRYl/h/JMF0zd7GKEZVuWwpTdA8aPIXyI4Hbdqj4mGYeAuz
JSgNbL7yqmZebs8wT1+m0Yp8rae9vmHGWXp3d/pozeUsV8/xm0uwmzpGYQ062pAW
mkjINjmUFbbxHlUB+kX/Kjv418vrPCwgaJ8FL0rznuU2o7KCxlXFExc+M6C1aRV4
YvPQdfC6LykoXqd5KL/zbpGJyfcD39V6CKJJZMAkCF7o7LtbplM6ijgEj6JleLZs
HJH9EQVU8CTySvS/mq/d2pIlzfio8CMRSQ4D55F0GlBhTjDh7sRNXJVDn3TEoqAK
3YaC9dSG9FoD2WkwB27vlpzh67A1U4Uka8Uye3mFASynrnJNFckY0LIGBtP1i0Dp
OGTq9uvxOe8LTKOoJIJ40KLMA8BPNmW/5ocLfwcMQDA3AFwrEVP1ZWTyf7ERGhyP
AmNFaRNgexdJr5ibURXJ94t4UofQ57a+Z21rcUqA21D1uAmRkNcOKsgqTky9Hf/q
CxPnQs2PTUxZSoLtg1CqwA==
`protect END_PROTECTED
