`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZI3CbxJ0I3+6C5C6ss05oIThzgF9TmX8IZ47oirL86AzKaJlSIs+JKUscpeWX/uC
vTNQmx50LV+UaHYK7Nr1VHgw819ZnRJJBjLlvjJrdXCFv/gbQAs1L4WMjE9J4Dhs
e4cOmbODTS0jSm3c4KLwxf8rUh1zWUo6x1mdIYf+fbZef5Q3Ia3uvu8Oor4QeG96
oUKwU1TLTzbnxHcBe9a16ihk+ZL3t7Lsnbm+KKEMVBHPMPrJpQEzHBRBcUTzflDz
f+/CT8CokmolfgCxcsZggTFke1kbvuGBIiDPkIO9H9P652+kammsEHMJoQt4bFmn
O9KdRFUO+gQdd1cuuuqPUx6bm8sqo02XNDGGG5uG5NOLODmeLZeHvp1buVDljnKY
krip4GMHoQf8eMGov/KKvpOIpqxBBSLkOe6p6KZ4JRa+dbZMV94byS7y5zPZOfVn
l+HWZlU3AhuyrbkbE/Z2fRSHJq4Lm0noAOKHdCM1+sjOGk5lxjmvbe23oqMlqt+G
qnBWhIb1D/g413XzkAOpknZvGF2EYRe1mOAnBSim7/xZf0w1HWePwXD7cm62de6y
mIJmGlJrqMq+rAWaQK+Dw9zyrY9dr3LCBkBuB1+Rv1z+tyVLFf9+RvWln952s51n
2A9e3T+BlPEaCm0XivQFQYu5o87StsewxRta1tsVkmMHij44ZkmMXDoZM9WJvptM
F0hjQXk4xGWnAnQRZSbCBvEslaKFoooBgemo4Wj28OxDUcRxo1D37VcaBUIbdl7a
/LBfa67ol1aFfY2RjdRIDBVaOM+tpI6gvDOPCGzY4DHV+buijLHO8h3Gn24AItBy
f1rugIQICF3hdekpoC6Bz2uriK8PtonNXseaFEOxoRcSUq1k9XblCwkpdFwy218O
66ttqDtee4IM944tXubhgrQwc+CyM1xSPiJprt8DssaZhr9KNTS/COPsPOUb/m2G
W0FNSutAgfZF+IddYBA1NPEhMKeHru1M3SEfNFS4ccJZYV7/9sKpkgWJRUgVuMQt
mtMJ0mfIEJYc6ShjpVw1B3CQIjEU2FD5ELDyntCK7jB8IB4asIJqWA6+G0xsHHiD
DzUtQ22MH9ISFhTA1aMQrT8SplEifiQBbePer+SWQjTll2VatnLslMCuti+EqfGO
P99T3H4GgS5ttCNZWbBBq3PE6DXT3boqLKb6THzpsOXTm4+5bK16jwBm3Ci4pNsm
Y4Z4S7w1UqyI/GbEexUh/S7gUx5qqWv9eZHOp58K5AjvfbtK4hyBQhnBKsAvbWwl
1JTaysjX2ujo0nmaqU2Y+V6xKHsYqgFicxuJR7KCxLfCk6Egdv5j7//GIPYzbTba
mZLOXPKn6LGfPaI/uV0D9OlBb62+emxDNWdL4/kG22L3sPCrSSDXT7+W28jcSGrO
+lBHBQbnXBx3g/ANlBvSNO9VUnFE5RBKkwLTu1ia8EzYnatWXCjPT612WZXMIFdP
kMLQI4B6QVpdcL0k3rTwKQHMPpUbfRVUrge6JbvAiiaDEWf0QcQtTGxqSVQTzoEe
Jot6j+j/KLKapnmQt1eemg==
`protect END_PROTECTED
