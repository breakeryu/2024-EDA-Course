`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFW4ZVW35HDdAGlgVKL3vBcKcpY7DP7MQwS+QCQGKuQH3oxc+qLnnON7YdzvfQja
U8PKc93MX278+M6iSpBexkGPoSeBvvSaxEtsZqeN7UwG6OhePPl/xPZmMYezC3HG
XjhoeMe3/yvWoHNUbysczxyygap+FlvpMjz/mVtPs8skIGuXF9SvGdjH1Qv6tQoP
mwh3sdjm1+f1mY6SRYPMBTv7rAKq7V0cKQCt1eZYi7IyN4C/RUjAu1g8WvcNT16w
XtVYox5Lok0rUEt1mJztMkaVtaF5xYjomfgVlzpovCm9J2ZX5B1jaEMhZDCxqQMa
yRGDwFKHXGGHIJaosQX926jYQ7gpyR4RawkB3VEwuBLUulpxlzvY2wrDzm10x05x
pRLTWG7dYJ1wdQsZNLiSZPHv7Xq0bODHyHu+KrbW1nK8bjm6UyLTBaqPP337iHOh
iBAh/JRUCsJeIfFaxGRfiQCx8rMinUi+cCZXEOfBF45ABGc5GI5VKTah+3jnexa7
q5CeZq8uoVfRzvDE8nJeL74XXBh4QCbytqhu/3swm64uFiTawe7w+g+8LUYmxpwy
pU1Z9JDwwKkOY/Wxune0yYMM2Q/0TLPxqvISnjBJcpqmsXFCsPUD6hZizUeBcXKW
/AocHy2Oyq1UD3Ho9ygTeJQQqpAx5YKLNEezG9F1O9Xa5k7zmfksQJCbG4QyMzC1
fiY2FjzV6YWKOeouZ1cdvpGxWQ89OB4MUR1qh57Dg0U=
`protect END_PROTECTED
