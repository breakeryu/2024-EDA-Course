`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKobHqQikDQObnAy5oyT8js0WzKdkZ+opN0VszT+p1F/UUTfmalnIi6JwTklhuFC
2OTifEG0dE0UnnUTES8RGXf/+FFkD/YLDYsuJIgMukOYsuYVPD/Ozss9Du2on+5e
tWVFjX/llBzyHW2fLsnKPBSMPX+qVJFXXEs+KCOj1yMEopL+JqMMTLqjaZ7cxgYS
z9ziqYzp//agwXR8YveyuvigPAPE1ff+FPaZp0bWOas8p3b5gs9JtAoWMsoIWkUS
RWoYrMg3/62IKrme4tEMuQASNig4G4aKnKAiqy+GrCKPg8/EpLIgVJ6CYssJbw+W
Tgioa1d3k6xaNK1RaJWFixkgdBZtELYgnFyGM79SOowWl6e35GCscZT9e9ZikcWl
5ZGDmOHsaZFPiSjKRNsASmoWyVpSeNZ6cr64s7aOl7G0X04w56LPFJ+kpfCwoLjP
eSOkUOGfQeMwqtWWUeGQ+3KdE9sei+3cb2ixxBl9BAqCp0M/rFs3OWje+Ig7OWw5
IQM3pJXi0qWBJZfUCbdycUwW7RNt9XshlEkHv3t22jntDrfmrOT0eWId/bO6O/DK
IdoeGPIkzCNHZoHQB5VoH44L+fbBIpJHsOZJG/vIXdlq2EAVH7RaHRLXV7JEquoG
hsFTP9xnyCJ6p76kFZRuPaE/SGXMAD940ARMqk3MQWtdg9ha6y9K5Uhpk72drAg2
QiFqa3WyaKRtZ+mD5WrSZwB9DDp6fNGSkIu59BlvzUvZOL7NgVaub2m85VLBQ+Dl
X7zCfJvtoQ9Yc6VSOhHJpxUkpWSkYEGnO3j5Yi3MBP/r9FUo7H1DuF3JL0nB7vZq
zT5fgsWO7I/AQ6YuGKZd8xBpXXbYGNN9b5HoIvjOOUXBj6J9FYl2DFRoi8cHTbBM
N4f5jGzI95MHOg02InQDOVmawZ5YKI9HIoOnnY6Pwee2ccjZ2wCvmRfeZo9rFfiI
bPck37BppOH4z5+9PWm0DG9/xJYxwETm7ujpromUQPmAaawS32Dn3MAYrD2iN0iS
q3fSZ1EnPRj9dYO+Xje++sFb+QJ3ueEoRt0WaFhzuuUFqMVFrfWYAki6BQ3/W+jI
rnF8ihXlZBv3XGUtUREu1B6aAEVt2qMzwT6aDHtLikKy0mP/SkwcBQcMHHP1uxMH
vWtq7st2tMG8n/ilBNopHebzN5eK6KW1IKvpXvswVgUXGSLMPe1/gxFlrE29Ftpt
N4nmZL/VZ91wdGIwz/QLWmJ7E8RHgyf5lImYH3eNYe6LuF2wPdKXcoi1qUfOncJ2
O4sineamrGDCI3U93kQveRWolfxFrH5ag7/8SWdAOjVQUfXxTVroZ0M5hQTgKIEF
OyKFq/qkxyR5XP9Axu27njPjH6d1cVEX8Yp88U8isidra6DM2eK+i6p2nBtGDyKu
9CtbM0yeA0Gi5GlPHrx1D+f8dNmU02o9vC2UMXT0WxcwC22HkUj42JrIWL+GzbCr
hd7wYNHDlUXeVynIQpChThpqUsb/dOlrAcym5Ve01C/RDxqlUU17lhb1CsuuKfza
yqZxYYPcevmGruQec9Phb03MlSvQK92Up7tbD8lgKGOold9rD5yMDCXxuubNLg7S
B/vWM9m8OnNczmNYvTrGbind//MERusBeIUnTT1g23v3SuNyRy03HxKyFTiD/D8A
wr3lsrdALR3b2x2QJhP7/QUb4k79MRGW/UIA5mwn3Hqqz+R2PKMWfUJUi/5wtwmV
8Ds3FYfwXQTTIwnVzh471B8FWBttlcjm0aVH4czefKPdqJq/hKqM7gi5RNtPsa8N
9KsEMdcMq72RY51ZRDz7Y0qw+AySXzHgQBugRYE44OqGz8d7MZ+8MMPueQGSqHVg
x2yEXCUSO0brutDByHZEm1ihMGQTTavpDE2dPpUBQpV994VTvAETiqv6swv79inY
kZRSGhgpkErNcWSqoVE/8KFrghegN70fmnKyXCXg1A1Z+uigZNAVl9R82KuB1C3j
zh5C826Y6T+QX2DMJwbDlp7aNSgiLPPzKHO1uALGzAbrdyJmkl7tkeTIqlXF/rHl
mvsjueaDhQ0uchWcpIbCngozTydxRFU50ZHV2HWIBe1U9JhoB2v4j+mmw9/kiO8D
+HgeZEeOgqqESJbNQ6Zs3kJilj7sxb7UpkmIY6DuPIvGRF71nfSVp7FHlpMKEDUv
IfqT0ai9mLCzmgz392OyF0mcK3inK98Meq7r0pFpj3AKmcDWYGEFTqukBwPnJRFE
cERi/M8GstyQN04EtHbgXfRCC2iApmxjSbsxHvI4Dcr9bUGdGHkbeuwdDPlzRZH1
2XSLUuG8E9y6e+0inalS201c+AKtbjtc/MiS4zjRGmK314+CQ3bAG3p1s49TTlYe
N/ZE8ebLXSL49S26WRvZ980D0wWxxlQAbYimEX6Y7rLao6emIDDGfj6pCB04PP9v
dSoxF+BHSAQNx6lSoVrfuWQmtcjF311buDodkoHXuFIx6nvKDIf7utdJyfMAcL6o
H7H04uVjDKst7VBuF8OpolL1TMQvN0+BPCl/Fx9Dgdo0zWIuVL4mzx2fFXCQ4RIn
OW8U9B1mJ1u1VLsHtFjRkxoREpNzVYBn5AKUcEjtBJCHQl3yZ6+15nTetpOlbXbK
OkzPI8Vu0C7OpLVu7Pu3nJbMonnD5vtcqG7CyYsjyT5zM4xlRWsPwl0FUFGa9PmZ
EfsOTinT6zFURCw8/Vlvs/n7j6taV6U1uibP83IYGJHboAxQb/mIChTIH3ZINBrX
BTKv+cBnqiMeswb/mCtdeILi3jihqsDOZpwr5P2UC3JBtatYYXRl3hicIipKhrpb
1XXPQGqVpzKi8Jta6Vr3/NJRjS2eS4rwhUcV1IRazqwV2EA67athnHeUbLrdJ9XF
+A3mLvgxpNKBL3Q/6rIHWsvODo6hIiX7A+b2jl6FkYGjRlSBMgtui+1kPNEsi4t5
Iw83JDhD6KjXxJMjPrHdc9IetG+xWRJOm4ZCLwRSAWYxw8X1+UYL9ZRC2hI571qY
dh3DHyOg/YZAacjUR7im5zHdt3Uk5EjTMcA+H5QwtWz32Mf9JP5PNAq85NloRMbR
gXJOyofjuWMNi2FCGF5Fwhfvl6TBUVFTMYCmnXY1Hjf1uVQq6314I0K2j47ydmQr
uh+UEw037+cZ4O82ijD1ZK99aMKeexxw3mYuuqpjtfXln3doXcol+hCDWuQTXQSr
hUELVSeUvLr/lXzMXi2XLp0aVE12A2k8BCwcewESmkGrglIXiy8SK32HAEX1rowr
1PbV0ZkMrYvsODIZHNrBLhany0B4FXs0Pb3Wm2+NXQNd/yXJt3WVQ3DMQpjULzWs
OHbwBUvz1TASHAXWHxoXmqC8bBD5a2ae8q4vkYFLAUHs2oXJdvJ76Pce4A8zgFoo
Hj5SbCFqcc8D1W+vor2cbveSS03kfHKW/mfgK87NbIcLzXtFYeRhL/sVxiwq1Y57
DxpvW2nBFuhZKCwjEsxb59wD4aYa7fZd5cGQh/x7nwYkmCBRhojgSmn/KwYuD2iM
maHVFHFj9qWMqd75dN//ttzwDlCet8AznYSZ18v08SqFvD6nPvR4uS0bWzf2usrX
3DkbbkKiCP1PZHCD2TUpbj/NFLZq+TWFwCPWGqsP7vakId0iJPNDCA1K4ngfSkfm
TMX5q16DGbHNLGWROzmlhd2gTZboF49Ucx470dUlKCwDvAd1Plo2s45XZUGcSPVM
6knk6dqmfmTVXdCOLkRejG2DzrM76HOg1ahtBpKTjDjARKNcNUwZG2beE/ioyQ/p
UsFGLHugcbBJAeqGrlCNnm7qg4UDUsuvQGzOUFSPuB2bjz9l/iAwgvHV2G/NuTfH
am904gW/ze+v20PKK6+J+XMtySLR/LiCo9KrcDGD8bMXFR+W7oI+xFQFBAr7UoqE
+8KRRyuh2ZurxPAZl+/JsbGgNRKkJ34vu91dY8LLuWhZr33aMWKGDvuRRFkg1iX3
BITvVJKjJltXg78vnHJeklQihp01bPG79BlkRjYbEGi0zLDsMkSm3rWUngTuSPrA
uLOx7rI54W9wxoeH4gwssERKAdJDZEMWOMiFw6BgkFBRv3H0j8KpgWw5BsD/w5Lw
OMqoSMcWAobVGvW3NBKLNMthbP02JEvvFrGXRIn5y6qVMMsvtbJmJuyow7/PF+Vt
t8W+rhkDbb8IAzYqb8iJZrvas7miN7aYqtZ2dwNiFN5MeHDgHjic1J+jDCJdcfis
glFsVsAKOOGUdpYWatpxvBp5/SCQcLkmY2UCe1ICiyOiTPV+xfsw5NN5uYwlmQng
lucurIp+FKjLbSEwLVPp3WBDl7P5SkSzlWNFqz/IdMRC5bBdSv+UJW+eY+cR8zZE
zD6Xq+ALltDSBl9v4TTlPm/UtLyFMnK5qC7N00LkTZw=
`protect END_PROTECTED
