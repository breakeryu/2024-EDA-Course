`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ym6VqbOVz2F17BfRl3WMZ4YqT24bYFIHhGoneUCMW5H0Dhz9XNj29fqkhSByEna5
fBg+qa6Pbx2+8lSmszH19TZUYb2Q/lqNgKrKAJVCcadpkSHC5noqS7zm8/5l4pKh
9ljpA65A8djWeufREZv3wMB71Q9q6RZbIJQhBIxaE/z3YcX88fq85r9jLW/zB9XV
Ff7oiZk7qWrt1DMQVgyw/8m0ZJb0iR7ugYN0jnvnom2iY+bavn2anD1dKJLNOntg
mlkHMxQFPOrFJTN54l4/gHvYxN8OghqsEPX6f647BLQVjGTD9ELTNpesaHiukv4s
m0hkJXNnwtorGH52LTasU+7jImFeTOREOOAzteNK6bizda6k51V7pV2E8IMVkYC7
iLmSw5SeQdpAkZGVP2x+dHHQSH4loUKbOz5etf3xb71cNCDnFnIbl4sVpOvVAsYQ
hY6z2iLV4ISpFfby5nTATWYH1JwJBOwQZlq3s25qcyrVOmWKrrhwoXr4o453ggZl
NWWfku74Yysn2nzwAE6jvIADXayt+QdnnY5ILuT1MI5NRzHFNFAEcWooKi86+DES
BUNGdEatoEWI35/CTiZDsHPKAtFmvDnf8Fj+YfgVVy4kJ+Z5g8ehcW2ZZxy6ohTA
vf+uyQAGFR5loseE6L1ck7zSMLquHKnEmEcK1Xg+g3ZQHcPfkZnqzDLDNrxwitMS
3Se7ODSCOGCu8lY3GA4hXR66Oh1MLjWsRIlDKdrkffWi7l+z/6/BSshGVw8xrhxN
VeC02XIRTtWfPaqarOMs6kFlA4EX5+HQsgkyzaf42TmaAF/YstSeG6lZpB5p4pee
t0psRPv1WXsWJxspTc7GkBg+CcWBY+dhvs+Cu+Q3P2cVhdpAnCUC/1JHtVEyWqRX
SjpbSUsb4cFRjqybF61LbezZEVlRNOuUu6e3U/1oM8trGnKjpV/aWLlHc2Pgzm9L
ffsO3KCEDlaGXiloehSmfTYCNlvTmtHGU+taBsB2+uqChOB4WknW/ObzzepguAjh
b58c60SbwfuGbcaXaZyZ9Z+DtvxoDwzYl3UYNy0GLZUGlD6bulyV2dC7rpuWJyxl
6xk/G5AfN+bv0TCoqZmeM2C1JhqMugxvqg9NpI6OCiiDaCDBTiL4scR33FbQjG33
5n2mkW/cum5IxPdbTCHP5diKOANusP+AGXd3/zGFrk/2YAsyFy39QUtSOoOwc8nt
fJkebHxokHPvF6HNrpSOv8Ra3qF/UVA8otqWNtqNVAoOl3/qLEcoNB2DxslbsQh7
`protect END_PROTECTED
