`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x1mS4cpdEwKzjD8JTLDosW4k5Q5qhQCAUwVym20T6iHl4jAQFEqr16cjIzTsPIPM
3XPJq8iOqZV0qiWG+XdIHT/WiLl67ssacV7Vx37SDK3b0c8xNGWoNO/GTIsM3tf2
vrAIIMMdYWjZR/AzWyGfKW5NpQ2GSlmzajvGrQEFv1qcxONCCjLZcm3bNeVH+v0f
rUXxxIZdOpMVIdVCLwwFsg==
`protect END_PROTECTED
