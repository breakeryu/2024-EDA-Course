`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+oKpxtRpubYtFo2slLdj0wlJahQ6PaImMvYgZ7oWYKyCULUwFKzz0s2zGLDXhoY
EJ8WHBfokEDCxGU8bj9aWgkcqH6IqldDN6dcdbFaj21wH6odlvCEnu23Rm5Uu9jT
5QsNDZIH65sm2fbhO4w1Ge+1pdVD47f6Appynq54ltzCgQHEv839XYzmMaNTt2EK
OMRjZlyOZliYH2azuOaYo4TYAcggAfNH6MpGy/umW2kGCuNsptiee8qy5A3zw5Tx
JE4z7XJy52MA6rxIvNGVCH9AjeTnV+9qIToTPmXi9nF0pGOgNvkiHEa1Yi8w+KCt
JHOeTQ6NtgwrUYogyLCNJGJTobEgHW5KuwTaDwRa16F2xEKaRwoMnTWIbJJB7a/U
0EtPzLe/06knzBUU1yPEXAornONeig2X0peYW8RpOAfIf8dEWWUxq5auDIeYRiKP
91OvwdhxIU6eSZuua5pnET3ZkZes0WCPsEEytaprhs6HyTP/SPGf0QupU8yEqOcv
HP0fAzCeHAjXB9+SUyF1YKl29bkney8xWRBwpA3yN9ROnT22zO0J+PysrUlZsPBq
Gp8Bl+BGlBjBC3oqMASfsKWDEW2dI9RewP83+P8kGRN8qPTd2lUVORlAGoz90t1Z
qjeaNKBAlB/AXl/FJ+43/12qxxfVhLg+s28UBNfrj69xkxIxCTwVUNN5j2m/89lW
UuccafZOXalWXI3h3aHNe0ndlvbb3NEVoVP4II4sMrOB8d/CP3JHiolOeL0XYZZ9
XdwNJUdv1indcV/EVbyEdpjt7Q7hLRDkK49uP2CRvUDobysfjXyU74csbN0PsNsK
s5ZODNaw46U5EkWuQH95LILvjznLDHAbAezdOfCQXaNKkptwcTfgl/BFURh901Qn
mjPGaHw35I0h309/XWqp/rWfPurkAQlFXdY7k6jYkr9Odu7E7Td1ASb1uNDFylsy
sBysy0ME4RM2qPLTFZ9BUx++RpEtAHPN7ENDSUD0cvcfZfyDx66Yi8ZbE53FWMv1
HB9nx/iGHmFvTALnelt4onDzu5tafczIUX9zn5LYlEd+U3aTrqSonXjtjnWc5Bx3
ToDlHpxHlElScHBa8izRg+kqw3IAtsJHNi5GejKbEy54UeNYEpfsBz9td55QW2bG
DaUzxU4C+kQrwdsiE+ONdRlFTNg+eU4Z0kuh6ov/s9OSaYk/n5ObAw7nd4n+dH/S
kBtpBCFBMFP4hrx6Iu4xtgXfTNvhZ7NUkSSm7rYm9Ck7qClSbOdquJQUhLdBprMQ
84ZwCkVMSRI46lmfjae3ExBMv9g6UQ0mIEM1NBDoQUj+2cc67DPY6cD3XN34rFtu
gjzb2gAMNZJ376rL/wh8yaa18LpFTTdvbNmRjv4sNiW4gj/boLJIAcanLTKYqj3f
G9K50/LeIBLcpv/+jkLTuM2BtZimdSAVS2UFdZOVP2A2FFm+uqEOVbnRjr0cZxPM
eg8EzBLjudzEQgGMxkxYe8HQaZg9svuYgIUfJTQTdapQIK29MDexzhtrkblmzq3E
hHT53akaWwXL1McNYnynV+1bvvKnPtb3Ij3Z7gMZctgpbbhUaMplgkuhgs+Mhpq4
NybwEwNwxiOk7yWkBtHt5uPlCFwfCOGkS/W8uIFJenoB7gPfYnHdfkyH77pw4H49
IZbehygC6BhmW8fdHAJ6Z5CcxaiPyQ0lEfFxBVt0RnFv8mbMiwZgu3ybVAdq1SCP
0X3Eo6hgeaaR298MbdA8CYNvbeJiu67vqhx979gQUE3NWqcVLBeMcbxpj2cLWTXr
cHZaGODhdCI6P6oz7l9B7g==
`protect END_PROTECTED
