`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cwLyNQ0j7FMvMj+UGF4WS0kXQUDdSt/3mOrwQ0JdxJriboKI9Kw/j4QW4EKT7nBf
9bpbByLPqcDzdzq8+5y9xDBuI3IQPfggitinfTLGSaFPEJrUlsq3AGhip8lahJkh
KOnOt3mNkyMvg51/ivob9MavOXd0yPO3y/SpcPPAIS92wRgcleLNKuLC3Qmt/XgV
rcQnQ/AAuyu38NozSIu+XRI0yLMvzv22bGZZUCrobJ5j5Dm/OAI34V7nfWaqtbI+
KxVabIQabulO5BBtCavm6VmxZzZ4dzyEG/P9N4FPIjMzaUTd6hFtJKwZSKiTMnBS
kkd0DLb13e2DEnqisLKRtvf3rJbelo1LUperh28KhGLCpxbCum9c6ZnyDfhjPCdG
U3r59hkFMxawFxoYey9khDddhT9r9EfoutP2Ib4lvYI2dnlrkKszf0q1kEDvmiui
zvoOkSZ6GFI5HQ6Ju3HEE+Ut0hItHo9XyT/kwn/meCdnav+dvPUp6nDoRinDJ3Ob
SZjqR9MKvTmNqMROFpwUiWsh4+it/j7X/YSrSeXlQ7d2/05PpladYoM9NYnLDdvc
msTF3qN9dfRSZhgyKTmmS3oXK/nYbFAfftU6T3shKHoU0OUXgdnEXm91whY3scVd
q/2mp7ZG6XIwpVZ9GPRxc5qWrWh/jcScDdj1GYp1oB0UFp+hIL6UfJhW8QVXy6Ct
JMgcaEsUS0iWbHMRR0Pdsdc/2rDcuf3NqK2bfQL6ahfPPm30u+UHPGowvUt6mHpF
OEbhY1eUbohe2w9Jh/TwOxfu0GNQzAn5tE982Ml2CWpevvv7PMJn/tJ3umAmIqEq
d2hu0X9/scfO6Kj1ww2+9mmYEOz5nKnFxvPEzZ9CKD+3YgGs+3l+YMlfC5Kg9LPW
dhtddBXjF7Bmfnn9fUXvpIFB9QdftzyoIll1YzkwiLabpvfo49CZ5wfYXKnNAgJU
7qdZlVA8Ok0kOdLrXFrzlrg0ZVXuzHIB6xTJzhmSwSyWfzfIWR8Flvb7sWfsrzeU
9uq4f0BnitdFwFwmaQnUnd9l4opx3UlWCSu7f6A4IzO/b6DXXrPPKt6NMB1BSnHS
YnJnD30JxwTYAPjiePDwppcCjcMjtF8KR6iVQR3abI7wMrpdHKtUoQoFvlWR5i4O
FN/wU2VQTF67S8s+U8uSAqXv6e7AMFn6QFNUEIjSLImKJ4eJxeh3APh36qkXUdc4
CNDCBMyIj92qqvaDGAdTIXheRPvg4fCOzhiIAFFF3LDU7xl5cxw3ri2+BYuGUVl6
`protect END_PROTECTED
