`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XqXVNIAjgpxfJLMlf60i5fxGJdTnTHgxRekqr0Ok2sZ9cZ08Ya5cDMefzb4s3JGG
dXM4kuKcztBl5Xzn0Jc7h+qEOY1E63FM5vPei9hRALGbSikCkG6lfS0fMpw0+KLV
nX+KzFf4md1nXFTzGPUV8iG9rxRl+BfZY4qZbEsj0ClnrCx8Qk0BacvopTIXGRvK
iWf8jRHp6XuXi7HdDV/sMpCucNfEnXS/tz1o3l/RCIrzrD26JQZyjbGvkTv8kdjA
y9la+YXZGm1CZXY3l/ZByTf+Urn/amp6BiJxIv3M9LI0aZiWFoN0vKG2DZw9Cpmp
MGEXIIni+HRF9A4wqbWEzinLUNLvG1VeU9eYtBhDt747nDV/FUtn9E7rB+siYOlD
TLyfrwtAoOTD7im0YDWneG293J5wxGXN+pgzbxpenE+0VKLpIltzyVZWhNIN1E1U
ccfxrrSCb+WKB3Xvsja1nNiDQT2wFk5SM+BVscPcb3Gut5npl6d8m4qMJp2hhWiB
hTVpuuC3ZgWQVMLRqiI3FLKTsg8YT8ykgEW7knQahkpjWdINYRwwaKgQ7vt4dJuN
dEnqFsnWINigyXuebWtIgB+7uUEpFV8sE+R3T/4MaTBSGbAmyoyV1wutfSBKePwT
igevodsc+XR2mEF67dA4Btxa3LWywa5rvl7FKyOflYYPSlvfEo1gVeKuSte2WrNJ
wTtrxCaLjqFBupDH4x1TYwNXnkLFyWgoJWjG2ZkteCwNfmw93cefly4mkglHW1se
1G3IgZLGgLru6mOK/fD2T+TeJj6zIkwvjxWg/U/adQ+nH9GhjNJwAzaqUaW1EUtQ
iclR6w6o3c/aZFerB+EtMAvR66IhvBSB+OPHxlL2ADTzdDJ3bHW+p6B1JC4WcwOP
7/e/y94qNvFB5S/kdCWbT2AVOVq+FHbb0yUm6QJUC6swghrqlqoARWKP0yfbaPbP
1abe+3zFperNZVgA9SltM07EcD1ddrgoMhP7ZAL+WErC2rKKDudFkGisTVaY9VkA
U+60YU7PzAdSqNT/PIukX1FLmhpUy8ZMuhGuCZiQ1Xl3YzArkp2zm2QA0DpF2TKI
ZNCsR26iTkUv26TtINWraxnePj/XUEQ0D1dlbV8HDvUxJ0cz+xMyL2TTlu/g1BEU
rTEMiGzXRqeq0v49hyif20JSeuGEehGyuIld2vaHU4qcrk6Wh4OichFnErcXTMus
lWinN8w8XumY4i09+xNGejZ0H+ZRVb+wHhbVO60uvC9wxKnAh4eTfLhIVB9hhqn9
`protect END_PROTECTED
