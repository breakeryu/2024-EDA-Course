`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRmOT/ecDyU8TQG5yNOGdFNEQFMk80Aa96uBqiuFhLlkatcuTLp8lfg1THbP4Esa
Sr5fM+R/mOoMnriiyGMkRK9zX87fCq14SZEJ2qjA3TAwcwM00Q5u+K/mWvoUWfTw
R7EdWJK90sUpzfMOBSXb0w3lAHweiV/x3P1BcjYji69lQ8NxjMBMojVjrr2CQkeK
hYghyxYmTL9X/SJ6cu0+/FT0/WQzpOcowtHv2+lznjMc46k57ANlFto1WR7bgcSn
a2nyHLLnk81FE0DLhyW1iiZlFQWIONiX7aD+/LX7oRc1sWaxNWRq1vDYGQMEf9be
BLV0wKTfIN3dcx61toybm0KkUIqDY46c01prbOkeH6xKlypxhVt86cDEiDTJzo59
cghmvAYamf4zsZ3h8Bvf+0V7Fm0tMUtaloQ+t0jlJL/eWBQArBEkSi5NQEevVQnx
+w7hWmThYn9d9zsXhtN3og==
`protect END_PROTECTED
