`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yZ5Cd5i7PHzla2bYT4A9hZMFo8JXwr3x2PnJAmzauhXc/Hjur8IG9vYniSaFutxR
7VbE97szXHcF+HWHrct0len+NBsjwwSlDENJ8DC4WHVlQ35moSQ2ghPvS1rWEUIN
zIcw/lQPWUTyxCv5/SysUGGouxYn1iFCo57IRAq55R6KYX06+xfnPCmddeInVLLN
`protect END_PROTECTED
