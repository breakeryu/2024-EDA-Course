`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5a8IDNi6T8vFwQuyNYjlGLYRGpE1RwEvqL3+QSiTBagq9ljbdq3flfKrP4MvHUVL
Msre2ZyHpnSrZbXj+nkaWgxxeo+bdP/hmrK00eJnPtEv5nasbwKjUxmEuS6WpMYp
1OurgZUlQGUXfUY6IBqvqP0/3F1ALGvRSCv4U1k2Zpi8L4xJJL092w30QR834bVK
Uy7wxXoXuFzUZquzio2r+6IkL1x5eLFrlAYlcWyMwxPB/1c77SuB6XqL0/gcaqBt
TO/HKuzToDfvrEha7cwA7e/cNYS3yOZfrOL4FjWD3TlIVcwJtdVKj0QfL59VjmmX
xBCsecISXZa4Cird8sabeMog9PRn9NCCHseHd0QMfsCrnUSa1/XTL+J66VOOOxR4
NExxoL7BO8jJtvpIL18h2mwoX8J2iQpf5MVzK0X5l6PP/xiJcdDrmfim7JAqobpI
T5/AhlK2SRtH5PojiLX4XTgArZzaDIX7UE5Pzml8bSHh+KOTzR8rY/5QrfTfJOWh
10WX/e2UBKAb5kaWGyxJTwoPcbFl5kmJ/qfkzlOX5hq+JMuTzOJA+zWGbDmjiahL
dEkB1Lwu9IqgytryZLTA7MQvFbx8LYc31s27UIFGV/h9o8ZXK43Wfez0Z7XHEt/V
T124Lj5/rdwsfuMvN6PKqitnRYGNW6sBSoxG5+f3ZGl3cq5ifaaHNqjUIGhlt5tK
NQBvAj7sNuj5Oedu9ieQjR4s1I1OC81SAp7D1RfrFd0gXGnZB2d2FDj2oeu92ufy
UKQDrVL14C5OfELJc+Pyt+cwCY+eaYLjnWZ1zgRz9cOj19tRXjH2WLcG1+EEDAEi
zLsYlz4lilw7/5Lsk0n3jVh23z3JzmamDKtitmATqqUxFfnT+3KxyiJtIId54Gi0
cGtf8xbnquhtt+rLM7MnZCQoTM32KM77lVGaRe+vfjMZUt0Q92kR5iMNFeh+Xv6A
42BSLR13Niv4eiEmrNidDozEZGrQH+C0N8ZISAjA1Yy4CMwklOe91GdKa9MCW7aT
pNg9OmeCxa1uaJGzf9wBBvB8u0iZyiSmqb+fAmh4w2MKhsR79DJj087hoK6e1JlJ
+CXnKcYd0zBzqHa5Dseh1G6/0k7Uj+f9RZzuYbyhSytYc6efQeCj8uT634IaDuom
ILE8vB6RtLfQ3fGotVykZ3x4Sr1fSJMeR6ZvOQEKIFUa2e65+0wjISLz228J9xaj
Ac5CRBqQs+cN3TbknajNq1e7QYG3wGJDeXeLav+/6fs84nfJzRCZadkP20enDIf9
8PNo7wLi2qlhl4Rw9sHeV1w0zVzOyWC/eeRhbyd2IFyh0/ZEMn2/Yc5XSHXJQjf2
qic9zzbRmoe6bndMOEyaoSAOAE0hikoLXqZYOFpafLYx5KOoy6wk7Ok/ukcMaQ4T
kUFC+h6RHnq5E90Dht2gD30z2Dzf7bYCOiUNaQN/V0UvY7kiQOWU4i9TaGBKVAbC
akKjSRTdrmd0CjpZ/KBMY3TKrjqx1iJA7SWKipjONcS7IfyB6B9dSCIb/vQ6qfy3
c4wfchXX+XVzCXudFQD9ecCoEn9w6PGnEQYkhyhdvaxq/hdRirEwtie3Tt9gQL9s
ZBbfrB46HQszOwgAI/KhnwOaNozqhfK/O53yPtXB0chIVaxYdzSim8KvC8ko60mV
lscSAyQ8n1MC5Bh5ww+tuSKIfVQlGng8xEZdMRPWXyxIoMujCIYPaD8GSP/09D0M
V9BaiyQLFkVOqzuuqXlPmSmliZqSVAiEyPR1MVefSjeEgnjmGB1Blgodb95fRUNa
IFqvP8V4//fl7arf4sP8iW0uNRFaeCr6WXrn2E2Qrsn/OYLWVPcEfJ0P8u3kRebC
Ot91MRhBaqd21d2jM1uWxmz9ZwQzZAifilwGqbV3/IkKD7IrBebmGXlwWg9Puw1f
EMv1Pw/rDJ2rWlJldlwgYAd0vkT2TbPWDZuZhrKFHbyKuy9QX8I4RtUDV6Jceror
rBFA89knlIW8kWctfTxikDa65byVUTatR9pJlHYGCsBhwAhsIYBVEAYQZP74eHUS
mySbB2xnoMcKMZfwAsHrM3CYoIVPTfNEbRMtgHDOomXm7vUZ1ZWVTrR+htU7EjW+
QF0CxrcZ6HOAF4qYIIXj3VG8l+pzz3QTxDnimAI56NPM48iwu80LDhMPZJY04p9K
hLivxE0BHT33IcgZbCk2JHEolmFKy/SSgZqLXnOwiQ3ECu6pTF+3xTCnDWQArOqI
h0GezicCXASflHDgi9s/ga3PIkIMXy4DR7+RyGjkCxReQN/jKgn77gVFh0VlcwDb
1Bjboqu2/+lAq65RWNWxmrxK8KPv1hHr7J/1TrylZh1RGd5Fsrjm/g8SQWD5SU5N
UGWiwJ9B+4UDBxTtBPSztHOh8OCBjXesm1hVAymjAP9HRaBqmt+qKwqk9tlvxx9J
wcwFN0GuYBwx6I7nEUNpftjNAOqgT304AD3xycRAwHRQc8GomXc1iTy57fne/QZT
q/iBB1IB0D1dgNwsQd3UcEfrANTfAZjpKZkbLErs4RkCk0nX0uLOrOHxhgo+gFM2
/oVOuODX58fVzytWt5Ph4x+VqmC7gMm7KtgMVsV3kTfvI9MBLwX9fVQbgb9qbBB3
xzebxBaIcqVC+RfgHFmOqT0dgfuIVXlSC3KHU0X2KOCsvt4pcB4sAcdx24MB2MlH
9qmtedcbnbtZ/zxk5plCfarjKujzxohCFLPpAJbytirVUwaEX1SVhRv65ts0kGJR
sv/I62B7YfqaS4I+AY+vxVanAeXUFzCbBkCjxs4BUcOPg1rtPRm+YDIWj7Eli1bk
hojNiwi2R0fGd+qWANNasO8HMCBmQxro9YcWjgTtsPVIRoOA1RHs6qcMby0jPY+C
75ftBnhIXlyhIQ80YJTh0nB0G5yo5OJlX47xk4+Z7XRd++eOueGwuKvMehYflduq
muPrLfdbKA8VKa/tldR90rypq0TGgcRjhR8BqewUHAJWn5dlS0mgRz65D9NkF+F9
rM3BOCfp+nPoE/hpIt6EV2xcwJKYBfkUT4un9VRTqahBMAJ6OATRRISbpk4MNg0N
fU2294FrTsczAfHtXxtC5yM08okSY9eD1ZUllMhHu36MF+hbT9E4vSQWjL2ciP6L
+gxVhO8yJmmMkVauyOOWF6lTeKw/pqvvnamkpcGSOoSOuYHvDfciUEM0udWdGg77
TVS35NPtB2NZpA6JK61aCpKPrshEm6nOWR9l6x0+WgqDJ8gTIGmJKHaBFEcqGmMd
7Kv6UeJuKOC+PMpKVdYocDD+wUpvZ1Kk+iwUdiMFutbbVKL+/WUYNWAo8Fi2wogF
xoxFDfGK0l0enGu6TkHsUfUnpIO/RdTzfI0XWZW1ChykEUSmTJSFESq7XZigJF+T
1Ei6MvPW313Xhtuz/mj7KUk9VmCbDvjfr4sKJ8npqdx1ov2g2p3gb2fJuRKU4hpm
uyqPMI9vLqgdm6xRbxPEeG5e9PSUFTXQrw7HdacMbS0no57R6s8Z5d0U//xioavf
c9sZO7X241sVKeVNqWAFk9GPFRzLIU8qhS1Rg2Y93g5Ri9zcMB6iKVhb9xoxwIby
w5SvAaE0MoZOC5rqACOqW28TX6x7cok2uh8NZXNR1N4izHbY9tkTA7OH7LySMbyz
v32mcZd0HkTxSsB5Y2GKHBs98Q5h8T/Q8iW3TfPraPAbR3Wu2K4rBWj/MA+xyKFO
OisITWiW9z8UZZ3rAPJVdTeVcAwKCvPclUa4c009VleE2dccvzYWQLD3crtNBwiH
qzJF+R9Pk7LabCIMTr6oU65ajUL+rzSeV9uSPmDKixpe9egwGI2UKuLU4QCCW+4x
gsvP3klQKOSS9jZISjwlgE+PAPjvP9qGa7KYukxDNK7TqRtjywknjiOlR/eFw67c
F8Nk3tThTkd5hlN86CFpqTSrwh4raRaIGkalCnPtN05HkP0Y5YpeZ1W5joKTjIDZ
j9B5SDuQCs9sh0QS6kbYZ6QvSDnfSxrxOUqp1TNw6izeynle6yE4D5TqBXTVZUxw
7/wrGd7F1JSABJS7q0wRec7Y8vzaLMgsCBDp2mRkJ/Z7KOPGvYLLZjthW66ZphP3
1zBwkEvsNdUorH2z/zAwp+HwUtiLJPE7OC7s2ItMsaaZlZb2CYWkbFUJnzS7t+2M
qs2UmFwu7orJDyCpaeW61KUkHNAQrbuq2ZWl12TR8m1paWtO7Kn7r4j9l52RMOc1
fvB7eNUcMhF1YLHGvbckOOeuRnuFW5MTA3dP++H+YM1Ugkr0DKOkAQ9v5nBnLh74
VB+iqTyOO0HkUV8NHj0Wy85f/JEKelkQU9On1Hfn7vHkpKwAbAo/yS7/nSe1lAaG
AE5EOeokV5YL9n/BxJbudoLb4GDCNPuZWk2GcldEblQjy1/0ruvBo78ZzLaAQkP+
wrx8o1Eid9mSZBs4JvAYvLenW40V4zc1Lz2thNKFG1jeCWrcLdzE0cEHPqVSu092
iA524eWxncROR9kG+xMW+p/4oq82Gar6DkMCz+hx2f3EcqzgNApJCoUMqx9ifD6J
B58WMBscA5jvOdn3np6FZU1EIkMAAyUffLNFdCi6Blttssd7Rje9tcbvr8nWuKSB
`protect END_PROTECTED
