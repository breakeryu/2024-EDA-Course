`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGRa/L+8vUYo4UfRS2bYzSmkE/VlMFzsx4c/l0qavulXiw08gcflfboT5YgEN9Av
MmDWZhupmLvdI2vpn5iF0FWesPXc2vkps7RATo2YYkjfshEQNJIilpYnC2Z5LeLV
VA3eLimPJbHBR8Y46ram5C/++ZuKWSXUd6U/W32VkuZBBmiC328114Qe2+nfTa4M
X/Qd6q7HKd3Rgyiw2kLbv/GVoEL/ig5BKAnEFU+Z02zCkwgiwD++ZL8kv2h/DDq3
tVD/m0ehv8hG9KkWQLRS4+u8NT/XcCJf6wEhLIwO9EKW1lfLd/usi+6S5MbF4rjx
4k9rtTaPCkbIB3pgfeFeP9n/1EKSioW72v357sl4rqmo0xStPVWpeR++U9Da49EU
UZLtw8F/64JqNgGjS6n4JQFJFBXF93q1zjQNCsHZa935txEMYVBDlRXsuN1XFOLT
kWfBs5fYoShOgr0iaVzqqCFswzNv+XvZHITsqsQJ+4g8nVTVDB0fkv+o7rKa+tp8
PuzRApBGj5SGbNgEiRqElnlmcvVi6ZT9dqglGhQH7jpfhSQ8RA71d6gbj23y9UtZ
EkSHaqNuoeY4kK62DXQd/iYUvaK/dBI8yjHhY3zVhYCSfSJRwgD+bb4wT3f8XhJd
ROsW0GdEE/iyUbQOMtBr0Xd+yEBqKjNFdmLncUGAQ0OrUgTCP2Q64PilmGbZFuVz
p1g0KZ3w3Fu1pDpl3rXuZAAfZNO16Rm2Lqni5Qf9QwPYrVAJJHWoBlN8j1BIOP+i
kK15LehroM1salNdWJ6ZfEPqjwwQ+oZ6cdfhFKMz5rzSU8hafT23P/IWRGw1pQMh
A+LJXciifr24vGhmFXsvDip9y20UybtkCxc8RDj6L1c/xi+qLSgOA1kVVk0/M8DN
WP0sgRT8GMDxwxu7wRsCJuSEC5I39ULqyjzqxrzZSE+r6k6Qw2WWHDzwlBmcOXnv
2uX5lWdNYUwo0733oXtwuJzYzuPUoQz6Bbe3vCWJ/Xr/EIUpIFkDUwxZ1/Ueuns+
BOAAaGS0WcX4pjaxJWJeHZOsxGTNCGxfuZveURGrI1hCTWlurGeuQXrgyPdo3iwn
3hbLSiGJSIXRRFhov6Wo/VX6nJsRcmakuMNY7wKoivRojGgrWRwd9Tcb/OIEdWUY
YFfvolJjv9qArBJVQYDSucgcxIdfFXXArqOWKzMtAO7at3aU+/btYpjoPNiIfMjx
wwtyar+bjgJ4bxnRb04Xl6IFwB6SrSLNfHIErUjPcrneAY/trM3BxwCReYNG6CKf
Mi8QvpKlX+savq2hMlVfuxyWVpA2df4TjOO04hDvFDJVTW7glEfsG2zwExKaCxMF
86wPuEHULhngrVPS4H5crSpVvtY9MAIKj+q3J7yVtWH4EWlyz2v4rHitSu+qQlZl
ZAhiiWOSXq/UUGXFprVb6tvcGGXX7wxy8jdywnM9w0zh684XP8S/6js8hZjzH8fP
hIJJ8ucuinOSFzZTL2O5RyA1qgfKLnvGWeSITZpIaP4kVn2xVyrgwELz+K8eUgTk
W6vXf2YuWQBljwpXYFOhovtXDP+ks82cI2NOdapk3GFJO7uNNHHR00xVHx9E1dSW
aIh3HuoJvzpjDZQmihq3KD36r3SOglrr9gUPGO1M4wL9uXqVZ6+LJCJsndu3+FMS
W35KyMwg5CAzZq1bUWoy+ir0avwm+UVMTFFpkG5dhPN4V2AlkaHeHsQu12+l8ez0
bUIa3GkuO2PQ3jF08TCmf2wS0qDMODYKLplJ19SfdL9tXzBjv30m9uE6HcGee7hO
`protect END_PROTECTED
