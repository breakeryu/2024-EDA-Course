`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W8NCiDz4vmdH3nXwsGr1dsp2XrzvEDNFsKb5bioyuSriTGCJis2Jci4N14Vsrpc
KAy6f5nW24wjnSWuMZq2uvL3jsSXewJLJGZVKUC3NPVaQrkd/encku03Vv0bd6DU
g65iJRAkh02sYwYTCkqoUDNGrnC4Kz1iAKRZaL9y3JBan+eDDWOjfh1sYoexgG/F
Km05oP4peput+JAymM6UzqX+ZMEiy+RiYl3+eEG8Q4u+vSlrkkoZ0x7lV9UQdov1
mgMgbAcjr/mMaOJld0zt1Kyb0W25r3BjLntLcWHyQ1zJGeX+LfTU5kO7oYZgqr/t
9EuXWCo+dhs0Ah09R6y4SBrCde97dYGXCeCXrmZDTyT9UFsx0O4iFWPnVjdqbaYW
rtvyhwdcwLOjZQwExuD5qZ9yoTL5HVk0bNgX+BxVMl9Gv8qB4ZmnQnIbctSx/oZm
bLFJSalXEaIyQLDBJnp6Rl5fVuSnRcUDEtvM8VdTdocsiLJRK8a8YVYAep7o2LOF
9QyLfcm2S+jU8yFG+As143v30zxCzuwNBVjlktAoW2kDcQ8eozs1W1pmFJoitd1n
c2qdvyXhJtxIgvCTI83X5OCP+Y7XN+C7wcN4MuA33151JUfQT4ehnuzh/wUtwJ1y
Ba0NhLMCiSbnos8+/B6irm7qFtb6H+V+5yc2OEHIXvVjZFCTFw6CU7YY/S9sXzo4
Aj0JFWm8wnYsYCHxoZeBgDa26t5oBEfQNT+36qrhOPBltn+kANAVXkrZGMeho7Fi
zWELM3hIVNb69FRwVlpm1jDchYzaTYOgdFP+sV/ekT4YeQl5Rg7jGF1CVZ0ffGNr
X4SiEeyuWeCUIxK7yQ+gd1yPNiDcPrP+vO/srfvpKECwfESGkwy44CdB9OjGrQpm
7XbeBHMLQG456Yv8/MYAOZXj6EOaEdz0c7mR3Q66MdIE4Lrgn+2pYYqWXbg181fY
ka9CURPVsNcdRfj41Z9r4jWPAQGC6Praldqpd4YPO+NqwDjU0EwrwhLRagcmxSsY
ysZWtmvU3JYzqZTJeMEjxek8ezQIFcb1KihlOVSfdS0AFA7zksG42iCAitrKXgWO
hL1UXzt+DlnV2nSJP4sGmuRvnVHBoJNLVXc+P7rdVIgxxL1Gqdxk0jJ9zOXIHcP3
ePnz2fhHpU2SXw1+qDrrGQnqIWh80cX6zo2jsjOfa4UBOBVnBL0wpwJ6tlQsQazx
bC43U1YEpjmR5o2FD08kOhBVJLUqUOx8ziZ2hqoUA5z+sGO3LlJrqJ85TS+Y2wnF
`protect END_PROTECTED
