`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVwF3BM7ctbedryvzoGFoYojz8mfn3Lu26ALEk3NqU3B9VacmKff4rTbUBWxt/83
tnBGF9cLKHsxl2oxyNeLnJ1PCyBj1BMHzR6RDDQxxZBoaFsmzaPGII6JAxK2Ph53
Ns0wDQ/p7aVNVxqHELriMBx6BhfhjppiIYCMl2EbOmBDVHpbXu6kDM1zP4RFQrbg
Z6nWaBDq2BPXuh/OA1dtItlcFzwzgK93/QkrWlLWLrud7UN2eNSBiDoFk27DEPN2
2914V+YZQF+DlFMIFzj0zNhXFpHk77RLuoxhRzD81Fx1mDMvyoFrQrLZtVoYzJE8
rCMTkYVdexONlncXrrZfEwyQotvBEC5+gVFAxakwj//Lt5yplXiy+dywVTfoClSV
Z2HiCB5E26eIpDR8k5GzUnVQYvNKmQwM6uKQsQWnTVs=
`protect END_PROTECTED
