`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DR6sdtGF7Wl1hun0XinpEZSwEz6i6G3f/k2cLgOR6LiN8FLd7tBlZg9dpVo9l5yP
TREVubPC004jGqw5G69E1wXuIF8/HSZrvA9rfz9iOwpB+UDLQKlz59LLfLAsASxY
aiTO0LBkbaFjOTdFdPby1EABHHkBMIH9nU+GxE4aJwrjTY4hLvb1ub4RMnohK+cg
AvpCycbb+1gtW90YNFbwUTO1VAZmd0oKo2pTSQaVSp2qO5qQScR6RtwK/M/Moaz7
MQCnqwVSJ4gIRW++LBXpekVamuxYvQFXz2NNeZn69akXhyL2ojVLhGZIQIa+ccnR
8aqeXNgIIqrzOTQfLVQjftRwkgXZo1/sjD3sYMzutQ8r5AoljA+DJxAvOlMBLIh3
e5MEPvmDvn+7wyNWTam+gXn2yaIIckxNwwbM0WShLrub5jtFJ/JzMO9h5N5M8pAG
wrwDeby3Je2kLvkQXWhkRHv7J6p+stR2Che8xfoOHt0ybjZ/M1r08aXzFn2sgc2a
o2DECUjbu8iqRiYiuiJG2G55zFmvUQ+taqqvO5tnEami5It99dHCnQHAAZPv7Lue
5tqWGdz/10EpSRCbs25SHY+54Om7w8rKRvOX56IC5Dkr5sumIQfOe7JPor1h2sIS
eM81NdkXTGD4pK2q/kXPj84SPdigwfrKYnBoAPgTD5c/6axAzz919sUrP56CoSUx
wpDJ+YbV3+ZR+R8y6e5GNnjWHssevPSA4cfH5pJMgExcWxapzgKuzxR3g45xJMe0
PFT7o8EfP4tZ60lLEuG382iHfZLPJAqOROckv157uhDpSP0Knim/G2zoDNqo+LpR
McmK4wzlPGZeQv1bFW68PSPWCbSXp5PY7hfx8YwZ9tUMh5bSdnTF0UuBYWn86BMo
iuCGsFm3SqXHrsNis2WDGNtfc5Q1ZykzChRFEauBsJEU/SROlnnzUxTljG4xbdQt
0w2G37Fayl2/x0R8Xxem46jELE0N/E2HWtD/owA6gUD0xZOkshEs76n8ihmoRJEf
3/jijGClRoO55MdwsNC9juQu25Vn5NvfpxnNonKxTETW5fLbez7phCyFRufhejdQ
BzAHVRlhpLfzWGrPztpoSurc7PD3XNx+txpr+2cekyV384HW0znW4W8I+iIQk40O
CBnU+f+U7s4ZQmh3LvopMLef7zNpL09w3hJPBo36+aGIcQZmMhIHxgL8GBz6BHmL
bbLrwVU1PTaGGD8lgix2lSFWR2eoHwCZ0qWankQ0/5tFBub9Q2M1uXA8HKyimcG0
DZjD6CqW3htHWdvFKrTh5ls26HBE73CoQTu/30m0zWZjkqKUimeVz+/hvZI6H0pI
KgslrI6Pvz3B2G+0Te7Po1b2XXm6A4ZFZglBr7evnqyxpFucw2hE/BAi6b0Pbp0g
LRAUQWUMZQvAeRzmMhbQocOkxCSnQncOTFo/a6jKMGs/qrq0XDyj3SXVoeJ0FFCG
gHQGzUSoqlt52Pi6ZRvg3tBlEBmu9LhK/qAo6Swpaqv80JeYrNqPS1NLaryNmom/
SVDNdhczdPWBGoe/W3WvBLiWJ3kD+CejU2mhzaxdrur65CF75wVx/eIjX+YR8EqV
qXLx/eL/ymudUozop1GLqs8LtngC3EjamENOwkkoHjXWsdLTx/xIdgIVS7U/Mehu
nYvnUmLVIhPi5q+XP4QGAJ5jAnMukYuPabwVPTl8Ch5TSQfSTp3PPXhbRGgO4aEw
KY1XtqFBi8ADf3DzR74HeF1QfCtk1bIWY0JyCqztiakM4V7DzhKhX6tHSC9NpTiM
`protect END_PROTECTED
