`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wuLfnhi12ozFXhRIipDACahtwYhAoSn3b5+5t6xF0w2dKCIXCLwyl5XivXwNxWl
SeeKC9+k0G2W4/95S2s/YvqdA6Jgw6oz8iPeqjfw/B+wKgFxNw3g6xL2gFtwHy07
FPJIInNSw/C7rDNN/goYZ+enlQf+5gH77A9Q+sTHnxxL0UUusQ1SoAuf8VCvT+xn
EIaWVoMR5WfUDzVadWUOa+yAmPQswJ3mx+/7RouP+ICQefQI+TBnsX1c02FRTdKg
5Ixvft+v3ZwM4AaH2jP8fYi2JdE9/3AKCpc5LbJlpQCkjewWkkUoy/pX5iBhESmt
H1e5ETBqrNzoM6GkGGe+y4O8sVZS5cx55kj49zC5aza0jHwxQYEazcZZOj/Lpat/
aPkyp7PH0tXm7s6JYZ3/Wn0V3HH3Id9v7CITie6A4HzaX7Xaa0xPpDNl3yFGD/Wv
etCiJh1aIhogOFbSymdnv9P7fpETMEm5kwncjkdoKX5kZRNSaGvbScemJy+7VT2z
ObG6UrAUbY/O0Dd3BN4SJBJpnZAhgrnkJqRjIvm/UzDPNMxBrthyTZAlkxfKc//7
K+iSqjIQEPhsbOQ80XCfwfETJYQr0CIhe01TttnU1wUDJUloDMRXrEYdtRGFrYLv
TvDM1UPQyYoPsaUYX7LHYlh1QHWPulnglLbTKXcs/rpI7tpWUgLSARpHiXkplkZy
QxE4MmZYUaysQD4l6EgYltqJuHK4cO9wksI/VhKkaU+ykWS1hJCjz4CrmJayxM6l
wKo5YD4rQ7M80+lu9J9E87SV4AeincqF6miKieAdw5+7a/m5Ye5nXJPq3TFEx/7W
+O8BRFpyEut89a4W207pmn8K+4QwEWsESpiHLqk7+QnTbFJd4dPA/0kGlKivJQYP
mx2vBFV3lUmd/q9Iaq42Rq7foDB/Qftla4sAHIQ+k+1cfXVBCwDncU8K37qW0Dxc
+Te+v3+ajy8Zd6t6S3gJm0G0HlSSGpg+DbkZ4ql5zW2iz7vo+BZVSl8ZCIrQXotc
lin+uNH8ARYiMP/VTsnNUk5gBL6xWvsyJwDX7Axn0dDi6jvDOhpJIOFQDwEy8Y56
M18Pi6io9gTE5EoKLCCCrWs9eFRdkeJpCOuyqvmY6EvVqLmYgEuN6bmiVYF2b+2s
T/gIRQyVa5LpRxfZDpXs4R23fKJZ+9Hw2RQt+H8sqqhFn+kkmiATm9IbozyuPfvY
YmsXzpFdsgMwOPNIicWXnoC5VIESQ+wihY9O23fqXtKgaZc0zHMSTcEwYKfdA8rK
HvOqDFKEEIJH7GUT/Sxa4yC32a0r7sHlo0GdV5bpeuZ3251UPNqXQiCXVHYeKFuV
JhBSVEmurMNfag5DIwnbWRoXVKeHGMHb6sn8ynmM5m0JubBU8XQVuTW9wApfymck
FXMyF5TSJprI5zfn4dUvEkS4wXAFyMiY7zZmGFd/+m9JzMFJ+rbMQhkQypoVqA4C
oXcdoGQfQJy4T9VFx+fZTcTiNoGvGbUNdJrBeyFqQgrl7sldzmuLUGzZxisYTvBR
GmYRY2uzJx33F6xEX+vgpLP1o27RnslpSfP/gnM4WPdV8jcApIBDpCLVv+LDmpUQ
E7O4tRT1tTSX2TDMDTSCbF2scVEu477OfasLKWwWYsXFN3uAorWw8zIEqJeHIs4t
qKwaSALa7TAfdeYvtQnoLI1Z1GRLG8iJQ9O5u0hfgw3RSAPtfuYu/hriSVnOfNj3
h8diHqcyU+XG7/6b+acNwr/hJ/EZTh/OQ9W/G4R9UBUY5p+aVcTGyjqnWxh1+5/X
K4SL9lq2BVsrT3esjCzOoOnFysSgPOrcQuAGvkpRb34z0u9NiKM74eeTTXulIubl
io9xEF8RHBCRnQ9K68L5ozMDfSZjGhVBw0x1SuAk6S05MXt4d/kmJg9S8XSeWJ3a
bGbGhny2a7yAArt6sdT4WDHOsMTsjpZMcPqiIkdQjO1IKAJBF4WnrzJWxF1af2/s
p+jvWiUUdG+tTogblU6T7N5vi+opMIQQPgK+O34HVa5HbfAl9niU0sULnnLL1YJT
9EhpYIyQrCkLEBN1nYDVQbBSMUrOhb5+xfOnSeE0vxnrvvTkx4NMyRClQpOvMC2R
iTcwOMuhSdckr9lNq+gR5g5EQT856Ipfg5Ch+xwN8pbXLzxB8SBkkoSgKqNZ4gNh
Fdl9Lor/mcFJH7D9MVWDrzq/nlmZevmVG3U4uPUuaHk/ESpjg58qJCVUNlelDY22
r0kHAUqb/AUtOaPZlZjj1VDxLSHiG2rejYHJWr2TOHTi9to2OwUDOyqQKj8bQJVL
ClHBSM9YsnE8tm1KU/+hhg/BYly2Cl78NwekGaaXlUAUWS9f7ReV5VduPrmno3n+
dI5qW7q0A1Furhkr0NY2B7sxs/CNjxT63ede8t3cmc7VVHPRPwjLSw3l17vyCDa8
PqDspAgHKfzmyEF758kXHDyDbJgJV7B+evmZ81uPYCRHh3Grd4xLYNhcKunCu2QU
snscm3hL8rTTXHk815j+AT99ssFwZFNKp/SL8S05PDEO+aVayIfVCV6W3ReJ89o+
jliUxkdU4pEUHzuIQ9hXCo8EpSEByRIkYhWUoHrf8BDZZWpVhb8jjes74LmMISBj
kSDzF6+42UVYHziX5D3GBJ9yS91QfJBzVysALrs3P8FuOCJZjjN602XC9V97shW9
TRX7b7nGsfEVlexBfv8lbWu+Za88+DfmaL8s2ysZ+CSSMLYq4PEue8ckdCNO/HhQ
QBNhO/+c0ogb4v/gEY7onJ30UJoStHeXo7R0wPjSbLOo1iWSMMzhlhk50HkPQIH0
HDqyJXXcdPOc7LcRP7LTC41E2AgbU2DuSL+lFaJ8h6epzk2azUXUQpiwDGDaSiGL
nm4ewjF1t8ET8cqRMUjEGWqIus5dosSq2rvcjUUQ1yPozywZSt7kWyqIl5kFJPI5
Re1CMQpnLii/xDM0PDEZziNCdDzeSyJlDuBYTNBXLnLk1Yag+xP+DnLKzLbr08sD
Ok46u/MfUW6Xd/OEwR87h7SfYuT+95968jNa3tWEDBeuQGQme2fWSh7D3huU+twO
AcJViIUYFENY8iQy0AzvPj+90lNfKEKd/EQupZq+eCeHDj2lvzaCnPJPsRKeaoGh
1VFvK242h9oY1+MIbA8HIjbUWM8BaEjv2/FxDY0Y0fCDvAERZKz+zXm6+tDiQZe7
6n7SQscnoV5pkMGDc3owxjyKNDomC+FsY1baOHGvwmU0eL5Ye0+A0tbqDTvw7Pry
q1608arHNyFby1HfOtSrAb79IXeBB927U1v1O8+V/3JRMJT8CVM6jvV8t0b93eFD
uwVKnwQWMrRk+YCBztpq3F2rb+DaZXJoRPnRhPuet+wi499cRysQ4pXru6Z/fimn
liK19IHw3Q2c++xlEg4ODu5yNvAOlEgLSpgf2KifW18tdRSpMhud7fO1zfrkAnr9
PRp5jPzurgtM7cCUUof1bLZyXrd6e9wgwxcQLAQA0zeHDFsYo2wc6zdsKE41eZtC
rx2eFcQvQQojTroSlVkjSO/8RXvlGyqwIX5QAhlY61NGGMfsKGvqSpie8U9G9jh9
bf+9wg2zalVP+xO9bQKN33JwTv7AtbZmowZ3wn+lth6KTwtoZ29D+mwuJJtwarCK
gi9JBesFtJck7NxsFz2j/3oT94zLoug1QTCr4t1eRZiQKY8AX57YwfCcV5U+9jd1
aZXW4+vqlBdnGS4jdl6Y5d0bPnaQnDvkPxiAlMemqVc1/lKGzFTRjjgVrUugKCYZ
JibDGblFxMcScTE8GkVtvgDvsT3Do3V+KYXAnlQ+4nvhvXv3o+jfQTztoniIPTnc
aO5SVgsLh6mGGju/9EnWRvBANdHRJVvuhfa8zr8eZYwE4v9kvkuKYzELHMh3/ntl
bRrBayRuJDFtDoTbfEgsownDbhdFBbaVz2SpUaz3//RMiSo0jw2C5401U9r+GciH
3DEv/opQ/ChHN0FmdO5zIGaiqdkRKJNbcqAt6dkuqqgmLjvU0UCdOPK2sB2pCjjP
xEBArzPVOdar7pmHEZNP3V/9b7GEh2LEHqHqhaAP0JekfJWjXzID6Q1AN98otT9s
3zuJ69AoDtGd0Y3gNHwLy1OYE3ZOWu6HhW2uhaJX674FHq4wz5VaKZzaWMW4ZhBg
a4XcavMi08Uy0Eufq9vu95sSOKrEVEIzGHjtEMM7NRZoH/92Xd5uyd/mw4/QXkCU
9Dc+JrGBsYPOru8SCiwaEOdu8aONdhMXLYW4YfT4IyqzEcqWxbEXlwhVaeplxTJP
ms4S2/5K9udJ5kX3LfLPUkZVfyfspEN/ltJl78jcPMVgeL/ev+0GYNTRPCspBoA0
SL/gCCKlFF9xVKmXgPaivocJk8UPWPuww0BFBbhmKfJVwC4opDSqchvdymNnr50c
ZNBu2k6KPrGTvaUDS3EdwcEZMjxcPWwM4oC2IQaLqW0kiXc7SY7c2wt6dbeyG0NI
DTeIsQVeHVDm1RhGqjO1Wf4j/zMR2YGm80yRsl8Y34glMmGEh5GGkRt432vpVn3t
F+zQGsat8+191udClq12PAhHdIk220zNZGrgrVqcl4t/B3bJCFnSxJLUhnM/VKE9
4LVYRDo0wl7CRY4J5OfejuEr1MZskb1Mdq0fVslOyDcBRj15gErgPf5pRzU4TJzu
fQmndaDg9/mhMDLsJx2MTzpv0H7gd7Sb/jWgE6G1yiFib08RbvTIfgv+hQxYxgQY
vQ1WS2QGM3RSC/YDnGCcHO5abiQvgs1oIWmH9FK6ab8p3pom/vrdJCBTjEKZWIxZ
VZWS4IZfXJJmY9IYIny3F/W9P32E9/vZ6SIktXaFj2NAyA7ALJ9ehpMrBOLRmvNS
ys5ITAPki/MnsCXQ708l+EyUdSawPOAswtFYcRJsuXSX4vMWq3cvXNfyOrQ9eKcz
GAcjEcGc1UXV0ltvJJflbOYNsXn4gJ14Hfjw9MRhA4q+3M5MmRnn3vNFDpOPAQeO
GClUc1yYMQqyjEyGZe5DxzkgeYJQ6rlFeZP9J2cTymrEJ+mNScrdiCuURvQKsipu
ZmJWx+SRDB6eJAz1XMjbvojb3gp6M90k5yIVRmrT0MthYd0EA+xv4ZFTxGfGbo6I
jakZZO7qvEbENzASFYsO7tudEqFOnpZAtghtpfYhsYaL9q5u3GZwSclI58LtkByR
HtU6fXMni/gUz4mSeiHhu1Vb+fPGX0TWae2eX5WtnDt0dtmQnNT3Nas9H34ngW7m
gqqLjI36tBZKgJ/hpTaU/gOxmPpw9uoUjUACU/iY0f2LLi/LPRXfCGvy0gVrBGTX
jdZimQpm2SrC2X8Pqe4+tVFcC7mpRsTNqT9a86wVbWpmC9r7LIE5R6VojdzjsC1y
c7ocxYIotSLbL9uFgmowrSTuTO9ES/jYOZJl5UXHL7N+ICesd2hVCSJW8LlcKqsn
wzYRluVpd/sQpKLRO1jo+iJgF62A2ypHDZBQW8BO7hEvRAqkx2J4iSXGKJKLudHT
NSZY2ngVNQqQ4BokU21DfrWxIwo65a6MUIDtIzkVBmylrOQdk3OvoBF4TFqOyaB9
qUr6cFxTOCRs+7YqzscNPykVkpKoT1OjvIJaH5ty6juBjEzD05uJCksPVLATVqEX
ul6H5owPLZIzvKnnwM1K1IXIvf+vjhy9Vkkm+qNPJqXPI2gCF3LXxSljfqblT2s5
0QO5he2kIY7NtaCrTSCUcxpcYtrL0+wk6zmeJpcFOO3AoyyWCr3dBWvg0f1lxDs2
wzWzEF19f+nyO0mCV7TaB2NbHsIm3G1CiJV/dbINjMBz2upqulNjy11dD/619gKS
E92rZhe9CuAtPYLFrJJFL8UPcDyABlCnFZcfC18t9RsghwI17As1dojWWS7k4sCs
J40DgpnVNXAEn+D0iqkDhyhEVarqomqchsga7J+QnzVQxrdJMFCkyjlWWrbhxCKK
eF3ZjeUFWIRXFTtgmx+sdUKiICdhd3dvWZ6FmCxbZICLLNY8RsOLJS+6v2eO3sd1
iVd/up0fKGKUtmbwWOz22rFJcCEBrWO+1zNg1nNg+7qxWUxYcFHzUD4C7UklN+IK
VUTc8OrCI+5vhZ7yGs6+U94VlQMTOXPCeuCfLgyW2+fJSOASd24tY9e0+iYAQD91
nnq1UonK7dn2SPvgcywSoeXZP3Kc0+hix9esWdkzg7A1juaoKldMuYKZdxSZTZyS
Gq44Uy1FdobdazZU8GeVf6W0meuQNmF9/YktW0ipUWpSBngFuxK57Uk43LVSgU6Q
/y3UdaVqNZyLzuJlv2yVor1XVkVt+WmTR2XZwZNPBrYmYB+2OtCz67TuL3sLKWBJ
fq/UojXaMQ7xetccaUwaxEb2wjADtdk3bvQxE9cB6YwoffLBFyJzfFUjxSrT7Qmz
f0CXrw4+QCIKyNve+zBjTIR7DBgQuUvsluQhltIgIvR7lrbRZSnkCsa7qQrNCQ8g
npL1t3F8mmkG69F3ySTTFJpRGUNiAS1QroU03O/V0BKfz06qwjq3WkpVNcEaaaOm
1f84EZR6w1fsVOwk/Kn1LLy6xYMrHsKkKlfjw73v1CyIHwcfWqYLv5bk9SFqwWam
IQKC9OqkNWE7a1WFYO5g05ir0GR4yHZ6UqV5uUH51TYxTRT3C1cE3IeYrn4kCCcW
W0z+uXEleowBDCdlz9J9gATZg96mNbSkBLUofSL2JN4TULjF11L6PItIZSEVxPin
BxgoSzetFa6M3nBpfyKASW0HEb9TMHAszCoLflfnbwX7TVz1HeiezF88wQ9wqDwS
y2vz8YUt75+i8IOCLEODCtiY1HMPUooEUAEEfGkYGdGtmAnVhEmpsFhGrlwqNGVv
oE5in8QakGhUZjWHGydIY621Sz/NzinReWTbIdKQnYy9aXiGj31juYjdBsol6e3x
K8OOAColmIg7n5OVKtbKkQizPaWtu6Wzfcds3TCq+QFd2vWaImyyn/BwRki2nB/8
NsLGvI9WDOzuNNui3H8CdQ1rCaQYwbJl0UD+adzKUMjd+0sWnY3dREXdPWBlAg7e
ngPwZAIc/TYSzmDdMHO+on3NZPulxfxNd7V7ca+mMiJmVYjTQyr92oZrFdjuxpCv
7if5qg0E5sOZFQGy3qgnb7HjBswo+eRvwGaT0TN9v0UPUD0JD45igksT2n/hXZLH
6CvzIezr+6aOggQCwO02wuKyP3dmyBJRVRQJJBdBTd8/kMJCZQtjpZ3Gs0vJ0oep
Okm2rCniZxCVH0lhxdfzkCBsbwnPUNE7Nvgd0gZEqJ4AQpm/CS/paUQ3qJq+oHN3
jXdHpjyOUtCkr4NOCm+oUuBGl/uOyfQ/KSWhoks8DtA29xR5IIMxcNDz17tEmV1K
cbFzyeGydMj6eeWjTJ9u8CxYL4EyTcxFCdsV5b+7rDHsMC5WHdwdGFkJS/d9BDDt
FBiNpYSqOaMVpmo6t6GbCTMDwOPF5wWlbz3LqkQK5sfA1Bbm+eDuB8lkeN12SaCn
jmWU603so5Kxk07nVPoXBd0kMMLIRiiwRH0Q4DxhVYv/Yw0BMiCScC9zVIVWYPN9
FF4B0TsfrH7sXyNiTMCWDf+AaGiSO1CXfEX196EGIM5kpLuNDKhZc2aeHSakM9Dm
0ULdCW4gkx5hE/qaL7Eet8ygOwfjSGagVl+OTiO3qtCR7UFjkCHHEZi63+7fR/Nw
PjVkNUEAf2UTr0p0zRiswa3+yBdZLzyc3/q3hDTufv9PtfhuFbwOeBOFDaMjWAu9
L3UUAhuI9NuGwkBIYhaJpzgmYkfDPnjsW3JqqpkyxQvlLHBJ7IWjABU/3rbXFewS
qi++9NHPGa2om1unFQHgJ2xgaZpnq3WxyrTws4zTHtcwqJBtosWdPCpYRDgX1TIU
ilDMCC8WTe3RGBilVLAED1jBLe+jBm3epJBmO5J9vBVnNvtrzJoaGCDIpV5aEbd4
sve1M39IyZLPkyl6Pw9L5ti1H1wFF83osemh5WipP3Of2E9gKYMYVskyhu2CXl/K
xcnsUoaa8Dy63qybAK4ZmpGo/C1m2oolE8f5+x4U1+cghFjgJUql3Oxor/fQC9HT
kMhfGOJ5/KUo5aIbu81eL6mZAfUtimIu/ZWdN/MtFkSJPqvvQK6lPZNvSmzVT2/O
2kRYi6TRvDHm1wvLIKVJ4Wf7GDPwSNtUqyWBBRbY8SfCuxT9glT6B3Ajd8Eff0ia
+2o7sLiaA2amp8h9mJfLM0qIzJPTNntS7PR0HAxyxlRsTIfTbAJ3SguWJFPsCOgk
AsuNwEzSlJb4QUMiHG3gj0KDkcKyagLHwTf3k9+xS3FE6M+LckZw2rvCfUpPqbX2
eR8r4+gDcMqzqoDZK2c6q3E+y5rH/1p7k/UtSmOmWRnI0lv6bPEGZWcqwItr3SF7
V5Ylaob0wff9HsS0/iPYTbQeJ6TRuke96oOgfq3W709yzGND5/Gnd7+Qj7NMkXfP
na1ZOvjaJRyFGeuX9c80LVjdhNM/7CnKjWimtuTYXtVI1x7x0Tz80qYOmweFfBbc
/s5NX7z5qCf1ugazlvhsE9kLnCupskWPqxtEba5nOXo5s7BhA4uUu1uqDqc2W4V9
rKK+coBq7liC+TW02+pn52sP7AsKX/t3ft8yrnGB1fLOSknFFwVfeKe5Lst3X0lA
XaknLrdrSHYXjOSBrY770ERDZds4KV0gshpvoVvXsEhb5Fy9PGuuiwCJ0mhjZyXd
KwKdaDSots/R8V2he/8SqdliO9bIbiq62NXD5jRsfFtV2oZTsw2gqjJMOshjTarv
GsjZJ/hRtOVkOvn0C4wm4jwC6XHXRgA2RY8P+p9DUs9CVrAks2XvESssPXOEYOqR
QJm77DKXT54r1DbYUvbc02dmR2Bi7MmNOrmQo0411WJH2Ri435j9VE4HTLbCW7hy
scygilKAO2sAC8lTly31a+Dl8Rc37yS267EuaMtZS+pczqkyrUQkT70Qoell7SAD
Dx99ZzuLuh6B1rrnrlxc8rtKCXMNgtYycACD9mvHbo9orixvhVHDrMzKOeCxQZZf
j+LV6R9N6MBzoH6r0EvyTjBSKRgRZfktBRTg4w+HkdrNEtjvZWyIYF3gCsM41ZJi
J7ykSrZptLbp47EbQgXZ6Y3vS4VXhSBOFxIpMCKdZvdRdRM1TXAeiyBysQ08OOfR
CLwLcljks1pm5rMtLWS23qtT8M51BsYktBPkA0hWfyuSykfjNgVm4KZuB15qBUNq
+HoYRBYfi9oYrkdkTQ/q/XGFZAVgBJgDDpawB12tvuhYntyajrQT/HyoY1rCS+TG
k7c6jHFrlqtZATtMmnTu2i0UL2PyukLzF/8nOPGVrRqa3MeZp7bXhsuDpJDvpLXT
FdCz14iTXMN3nS/cH8/l/infCU9jFuv7vzeiLDHb7aZA8PPQ+5ymbAIYn8c38uYQ
XgO7XQ2l4KJmV8fItPZnVs2zWk0YYELzJXLijIjd3RCtLGwJMlpja2KSFUTG9lxn
dlUlwjoqQ0KF2MykMJOGIXDSDqvWUhe0aUCESRWAwHzALOvYAjsxFrL1xk5jEzI0
Dhx8+NtoH/AnWgHTjElQyjaxQJljw9tGfrkAvdZZkhh2D9MgU0UMHr7I5KFsomiQ
HFjKs453O/xvzFqqsKNA3fj0KZM1zZtRsfB0GTTL64OJSUeq7qU4DunW7IRg7w2l
mmxjKA/DXx8cZtxZLhMnSiTQjmbkcKCmDADO7J916zwaFZhiMC33nmXPWdeOI9Sc
+m8rtRqmXrPdAjbIStasMkDy9X/DHO8DBj56CDQT69Rk1G455E2pntfcI3NTYkeU
HdfxmbGUD8DdrEMt5RfCycInX+I6cpfGDZPjaxpymVfOu6I/OrhHuv3CrgWvP50s
StGbS0BzR9yGzGvypNq9CihHZF8Oy2AeDmOK+EzR0jfy9cbQ150KnegR7H7LjpG7
CmszZww2qnJLJOJ+uI7rYTw3dnf7GPy/e4AtDAoxeLDIuhl5Wb/dnLcAWKiZ0Rdz
uiUAvsv7572Js3OBYkq8gYFZMauEgRmN8Jtk6hP9c7Yr9aJz1OejbvddUSC9Jrp5
FSGLrwyMVAlYihmIa/4NczTLv2SwphpozlGlg41GvefjCkYuqQu3aEBH+vnK2GFj
oef7pUQLd3/LjD3WiXZTlfrZMLbHyR5qnt+oKzQDf6/uMWEpUkJtzAOiCepMF6N4
3rl9TOIlJlKTE1KF8fQnp6iTeHprR1dq/OZsbZPy0r/ce6ylduOOpQzbc71Z4zwR
kpd8H3kpAPA5urlIKchFb/GvZ1vBwwpXajv+MbEUjzNWaWVHOkjwluk9JXOCXc0o
8Anl8spDzfVBv8v2ebBTneByZth4I6Ox57b3tlAg3hreVMKlJHhDu5v6XvvkO+GJ
UcKD0UInOEfLm45W/zs9dEymRhH2rJAjuWx+N9fsRNZL6Ymqtwn6FU3GPMl/nnpP
x3gBo6HYKBs1c9JIMIMy/fK2HzFHujYDnp12fMhBDV2LaNLvyMwPXEpq3sOPfk6v
zv046b55ir7QR5tOOviIIZtKBjuUA5eYbYV63VNYZIs/0mpIUeqGEf/ErvnzUMNN
l607J5kemNcfpOqTUSqugsqVLKliEYxmcrLQ5xD66f8CwRxPqUO7No2KLhkPyudW
DUnxwvTMYLtV79H2xDcO1QtGcHLqr57tohJZTQT/yZBRyURQxDEq9Yspqaoc2RD2
NYB6EEkSJOgzMUQUsaseAf0l85Q+WGClKQpyYkCantEDBCQ7siAlwV39RB3EuhCT
0mJmz8JZbSpBiDrRPauxuY5uLntEIN6kvFJ3dEsB6I6qpV9tQQua1oM4Q9Yn1iDw
DNPo0ow5arRDdsqYWZH4eiQz/55F2XmttCjqVXVRhazHTfhRVeO5DMU6p/gxiRyt
yZZHgiEnYnFbdD02PrXGeZhFuzVT8QvY2JO83wu5CU0BsYPJGy6NU7j59ep1KUES
vlos5nLbcJtQntIrN8zuNEr22MXAliyH4z+dnp3k2G98eWyRJBSvxn4upd0aVxAn
lt73x5UYSRNkGmvwBFuGvCGjyUM3Nbmcfy6odaBCPms68o5Y07K+PZe3q4ahR3+P
ZCOpjppqU4d91Is/gyyR741zvU4aAj7EY0pLhXtLmWNdRIWEDG19StEzrDmTrwBw
eqZtO6263CTORB/bb5U/f2w/R/lzRwg/c3dtNHfDFrZd9dovSRf075Agwn9vVNc0
hKOuibH/LLYXt0DGe5+XxvFOHFi94EoXHnCa4JkZLeS7ahbmdmKmYPZVEEpr4dX7
yyvT6Csam31YdvKR4JcyBz6MX9L2ix2mDbievX0myjCx9UR5dySEb7NCTYoVIoTj
yiQ/QpO5FcSgTXKzUDgk6cb7rA5jUiKwRt/G4yPPmSRZP9UloreY+TShcxdnE1nf
lNOCs3IA3Ja4DkYkiIueaAL4UpgFUOfhtYEd4K3lKU3iYexCnpySjKdMyiKxCMXN
1WPePxG6qNYaQe0QHSC9MY7BvL6RbrKSRsUvH/c+hJIWl9gysmz5GwZos1kYqJgx
4zW+jZi9OZqm3MLjIRX0lnygq+je3pxSNfsr2RBtabh62H/jTOVJHiTGvmWoZ237
ijzr/MEuxMsu9RIWyC5cNzy6XC6ukB9GIITEbKODNj64iYk2F4OBqGvZ779Yz5H1
ocAMYUF7WTCviD1RToJAt1g+mZjEOeSeAgDoCy9p8QCgH3HvrIan/r8k8IvJtkJn
n4H7Q7ORy3peusAWroKy8X4HU4aaatXqGxxtb1pZSzV78nCw9YILtjtC2I83eU7Y
Paf4q27VOQrlZZ7Xk33gUtFGnnY/sAiIffJ5hw6Q/YdK+j1htuYJvtjKbBdDYy4J
ihX1Dni6zAn5EgCwUsu0IPUc2eBYBrkPvNeEqfzIoAxN1q96qQKfMth0p8cfqELk
lu6JVdTX0efxjvp/rhGOzIvO9P+eSTdMUQABwP1PxHPrED1xLkiiohLhP4nOcvWD
idtAQwaxwtb0FKeJkEuBJFNH6FV3PIBVmQRrVorbDQWpALbjG/VjeFfmSKQrj68K
FXF6xqiiQjHLjEQ9aMywu3zrIxEKE9BuuOC+SC3h2VafQ+jhEJfnvFs/DAp9mGvu
VuFU0NIOhIimsSESVwTBoNz57uPUzd48cTqU6G5LmWFvKnXuwNHHT/A7UNUhvWZz
MJF6VbPzIaxQKYQ5TFq6tcfs74iHBFKv0XH/ZLQwdm/lUJ49Tpb0tg5k3pRx6SuL
Z6vFvDM+k7/rrmPcuRGaFGOqXzWA2Aq1GuSgI+B+GhQ5mHa3dkzct8F8KxN547lx
L505YrU5FKxz/u1NNZpu13y30gXARjqZkjXp8T0/3jxR7AnLroYhTS/4RPD95G/d
y0zi6CjVSkiat4/evJ1aVKZ6608Q0YxHEm602Bl1X5G2LPc49hJ26ur5mKaB5vun
yt04VZ2isIhQWZr1gXAgiwEU0UXK6tqD6HhXrj2LZp0JMt5vwBVTUHBs+ayFk1CZ
erFh5X1GHOBza4a7wWzwUY5oUZ6xj/vpsvfDu7HLtVs=
`protect END_PROTECTED
