`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTCwyH5wC0Cy5iqJj6cHEzlGO8mrQ0ecLtHk0m1nElOBR5W/9OM864V9VV6BFJTW
KnETZyLi8c04ltUbDUhgNSxEU7mhwMKd23OsfcFhlMGLKltlgOuWG+Jy8lVjj8QW
0zxwPWUADnY596nTtHKmdHsXnf2Vn2X8EmbU8zfP3heRRfeFhBrL5HRFup9p1/w0
VCgjvv9beQTpv3QWqwqxsgtTF8otSg4OtToHRGqLZ8ahGZ7Ob0n7nmw9TTK9hWlG
I2+z+MrcYQ6REmvtAFqGR4Rcgy7G0Hu6GvHW9Mx2fdslbYiUHMuAZBxNL/lZhyK8
NV3+8pYmFwbHUauf36nTCyydWNfwtXSPNNKjGJSE4W3QINoSXHkH/LEiTOIUlvPx
EqHhT1m12FwbBo12uFfGz8gyiy+NN2fLvu1I8QtYkY6s1tvRlP7/8OazJVeXGCsP
jvwiuUZxQFxDmfanVzXdISBFlIAxl1BbePalCw8XxjO50TOjrAFW9QrwoPdIuMte
WGuIaJA1OuhDj6rNkrfFSD20dmNUnI8ltPpdYYoBHXzNIR7vHezLBko8ghRolrOk
oqt6nocDfKrtbKC/S//ZFV+hB1x/DhA8c3g3V7ecEeclhII83cUKRm+YYQI57tP1
EtC1dy2ymKh+jz5VxK5nppeh4JMM7WnxM789Sc1zoB+nwcHtZWcGYeH4nvug+LR0
sXrjEMeNkVT6qF0LNfaon5cVA5A/xFW0Ci60xaDMctNlcTICkGlQU+c1vJVBXNra
DMIQZh4kk+fQT+ylpH3rKYyPeGL98NHgX6GX1pkeB6B/Ioc6beic/ys6ippw5XRr
+XiMcuxe0wQuMF+fC0wwqMzUhnjXuegAkc/ffnSu4em4cpIYxP/0nDEJbEDuf9wU
cDHxEKOoNaprJu6/ISqfkYSjJTTi8sfjWk/7FtywKPHfZGmag3LGtJSZtQgOCqqW
dInolu9zk5zlSdtJx7XHl7Id837oNew3Lu8zXgmxxNEUt1XUok9TBAZsA3b+Xjy3
D9kvQZ5UgmTqH9+71FdCGBPgw/8MIqIYAInXdqUyQx9Xv58mVRSx9dNxOu3nnSR4
SZQc1h0WCLIsBiu8e3QAkhQwvuPy2KLB2L45TFTKLTAL+0HOk9GARwvIP4X0yv/7
ypcOqSzeBoS5npZzdubkwy5kiGN85VqubQSP/SJuPm7PTBLDx+8FR9Jlm3yLUb3q
x4Fus/UuNJsSrt7ffwDzv6KPC3y5mcZ5JqKXQty/W0Dzgy3fi4RhHycbSYCLeviK
XC2KiVwBLkB7/Dv1hSSPnI50V+TknEsA/Ov1/HQQg0KNmcxZHqwMKkf1frbRZchq
iCAfxvQzaAsJdU0sLGiiLcCWYgHarh6MmMwsepKt50hOIs03Qcj28lUunUAg4IOM
FYAtWZkqTG3jW/n+KKUuQZ2kUpOvA5Rtwbdw/Fwdit2hdkWrM8WvHjuXyEMrqTCC
vd2xGiY3cmN1P9anGHa0dF1MvLalLvDb2vSxVkMMgDIKUJkouc1+dt1cbm1aIcC/
t9Vh35Y81lvSXz6ZUacCp1KooZaj0FnG6dt3igPQZttt14YaGUB09aWIXpwSocPK
Wg2r2PpJ951oltsGXuy9UTlvGRgZ8Il3V6rdLLgT1CITp43HvJ00JK+HfzShQ7pY
CYPVxf0N/JbLJLN0Vla+jlkOCKg9mhHkRdgAzCA45Dum+SR02hASpHBACskbP/iJ
v+U4+tc9PQVPxLWPlD5rT/KYWdR3bv+UVpAGKfgG+89wsXvKZIx2xPXJTrE36Zzy
QK7dkSWbxWJE0UBXxJMQMf5UwszUAxypdMd7Dgum/dxssTprg9JH3jRHpGBOourz
ABVIibgy6fV0tBvFb0spZfjC23XP97KMvvHwp4cNzN1QBgEEuOKXnUD2q2uik9JT
aoxVaei+RBjUlXvbSCDWi6K2wo0uE+ptDjoXEiZ29iQ0HaRYTVAbO5xq8p1nkxg4
l4k1vqT2y0qeUCmismg9CJ2nBiBjTCNDEb/Sceu1GgU/hQ2OIkDbHrRwX87wDUM8
m0ryg62+5oG6zEMzbVnDyd7vRE01IkTgTJ0xJhYMh+NO6pm5hxX70hn/pigof83/
3p4N3cUKQ8mYamJQsOSReZuHCOqFT8Evc92aVcjn8RWZmTVFYH927kwActQYYJ8c
cPZsuJciDZG8wv7R+71qVJiTJNg+TNE56JLiWF0hZh9xyC0uzieqKood7TEhTryI
I3zRe6lU3cS/xkE85yyQp0RAxZ6XOBBewzeLRepQ25f3f5d08XeMSmV1uIZ1Cj9I
z+5k0sQXTlPqKkPbhKbA9PN1sFHpFgomHXf8mpn2Xhe6QM1P6tGmc5o6EWTZoBAG
M6vJc5lD3+TK+/1FXUptSN0PFLM+S9f6erXCbdUjb4NuWaSNjvBG+6f2bFkpVDjS
2jKMjOU8ukaT9fjPyDXEYMQ403FfoYBia+HTWy1kxemODgL5HSJuKCakB1KVuf3L
HHpFfh4jGS0zcMlHh62im+wJq8WmevbkKjrcukdmPAaYEzofWFVTcZMcOsTPb3lt
HO/5sjNB37JvhE1/zsjvHj35c8EzoWlKqk6zB5lKZbkMNNBaXIPrmbxmIEJ8g1mt
f3UlLNad6UDQZM5l35MiAPRi57XZEVzycbuDDRZLbLOyltcfpAF2nlB01k0qx/y+
6GeWGn0qi6N157EHaKMsauqGe6/5m5ifeM0nckiQKH8gIsoNid1OXdhpcDoNO21l
frtSjEyw0KLLdsQSNQsHXjs/UJ4hliLTGpubcW54X4QNUCyZT9lzkU8DmiBOaHId
lVE2Bi9lPMSYTHqDdqIswta+ICIL40IVQqa9YOEZpDnjp4TJDygSJqcBKThXGanm
WNjq4pjYvxIwPJi1i9UnHRG30yaLsaUvGsqM6Hc+K3q3arx2UKep/5vx6fSpHQOn
xEm2WQOpUmxPYZRpY+m0bFOQPmebXc8Ir3xdSPKKpDibhVRC6Kv/GBsGCkfRWsVk
MeOL+vVyROk8rNxU/cNimN+e+5a1moAlr9JdkgGFBcqb919DodijrUfcovbYkm1a
rtQcR7XbSuQUiPVrQWIlt3SoMrPWe3x2R9Y+0+OfwErOsM53z1JpxIenmL27FGUd
KKBNpKu8L6EExlezU2Nr+KR+4QzzvmefVBrAbSevE7D3VZaJG7C36BWa+k5eDehJ
VDPfHkpwsyXbje+nSzoy9UbHFGY2W2moJS2NJVfNOsXH1WtFHvExVI+9R+ioSJ7y
X6/IqvqQL1XWyJJ8HnxNtptIoAk8AkG4uO6uvJf3mF95noZXpCfmo3+NvVzIYUah
7qhZjzRfjiBh4hqO+gaiIEtxQ5Q9C4Skmj6w4PtoPlxiHABHTu47bS/OfYcsOjj3
aLO+/zJRsA6K3cbPFaWM7J8srrqiLtqydtKqcJwGia5qpAJ7+YiJEwLDAmbGk+BM
IQE+psbk4vomvG23uoX17AyPPGSB5jpmrPWPAUnunTl7pMWvW7qxgoCoxRnzuDUR
MhK5Q2Szp1WwQR4TW4Hk86g1/v1NQ7MF46gFcaXuFEdfwzY7+/UDpw0DYufrok7U
o6CK20d6XOmveTjgbiVFIsN5oDjgvmiEnU6J1OhyRLqwJd1NRrPCY/viS+d4ANX0
gF5Vj33di60yTtZkjCqALBv13Nnc21WG6gFLEpLOMWztq/ggyK7EI5xxjIiJu6zd
obl+50/EE8T4clOMdt696HC7DIjhX0m+ShbW5GudQk+556R3DbPWJh4rJxEsOlHf
vDj85+mOPqmicihTt9/9980BjSzZnKqF9qdXPjBHF+fCdvtDs7A1PqXcDiD5JvsV
1Ns9SaawoHvYgG/f2H3rHVD6Kkh2co5A9YVMShi7VwYooMBn5o7DNYvAkoWmwp3n
bEiejU9ZkenOXDJimOUzdQMg2E63utUDUjShkt0PP5PltuKzVpMdt8jC+FIBOMlm
8XKQATILc/oTakA+f6bjRXUNRmeyg+JIFJejboQomZIGn/Y/JQc24G8kQg+8t7yO
4EPEYvUpszM/7XTaiX5M+kBfAroArVbmZNCubqaz/rNIDL/ypSk0HB15hScCpte7
m7fwOEH6kSHvWmn/UtJM+pDQS5kZH7tSTW9dNnlWwnf5lGmn8tg+FGmb0Yi0MCLO
XnxxBifahUOAYnQWWmZFknI2s8U0ol1mMin8+IjhCMvHZLSceFY2/1cVgnjs11wZ
JZhkz/M+8Nyux3ylctIZs2cpe5R5XS3YmP86O5h0JmtEntPsE9DHRUQ7GG5Z4E8M
aJpD7H8iAaAuS8dxDKkqSPSc6vx+d6uccHkAQc+LaHKF/5ktx4iQdCbA7F9tdOVJ
ZVHFYacwZ7FOeiiX2YY1s6iyFoDYI3dKCd/J1ZDkOnTGOTMGSRkdI/UKjbPfZZFT
4Y2CbcC4Z+nMW8irv3c6rX0AlSbEDtfupqaEyO21sUW9uaODaa5qUrXhAFL3fH5C
dmU/Lqwe9HgXn3CYGb5zwdO5FRtSaDnOzFeQjRyMLpdtSQHJ2msH6HtX0RdhN2mu
k2DWSdbPg60ziZVEzq7BTvI+VsGH3ne7iWenr/9Cs1UZpqdt2FkffK5xb3piViNL
OLNTdVec/I5GX4oWvF2ZHkrqmtaM42Wm+Jb1ymhYjVoUFSKtKJ0R3z/qIRqvx1q3
PkFBocQnuV8+X88HCTyVPSS5zhQiEVuXdCPn+134PjCuquu9mBkNO94ZN6jLWNnx
5llvWbFqB4OgyvYFhSjdQCsFmj2sUBB6NQsx5Cp6x1D74//Xy3n+fg+WI7bCdLbt
NmU4IGr+IJ1W9nhvTEtcem5k/j7q2De+HFWth3TFQO2o/pkN6Ia9X/u0j94a41t0
p0eW4+yfSsgsoq+Md8pWsWXdyrrxcK/v9tcBdySu5aBRjKOY/H77GFGwqw1dvYn6
IXjUd5p09mh9qAfDrlsZckZZsRijdBuh9HoztlcubFloOcPj46ikFk0eZiPLvJpi
ESe0oxW0FFQM92Cnu7h5SSn8aKKPi+/sZ9S04L/UTxLuVbzGbvpfMGkg/FdfbI7/
TFTL4zXCW62ccZ64o5um+g6N/583gRQJxfCRyxfB5cqnd3emgcFug93VR2GLjSU5
lSfiSnnK4O++hC+dOten0lP3esaeDoCdH/OQA4JfjZ0PvQfaN+byb5pVuuOUmunc
8n50DvEME1p0s6uJEiYV25wC3KNvlHNdlQuOUfV9hboxDdtMDVCIBJAN4b57cZlY
NqpC3RoH78Kp5wHqgvuFrklt8vYhRt5TNbG37axtmfVsSCdxycxfepi8tsiUVEmL
IT5KDZJ39TOBJR8bsXoOvevebvdzGOc71Yxg8CVoOFXVmI3Wd7Amu693tt2XGhcj
S9AvoU6lY7WaRZUzeEk/fpHXkBax78q6wMb7/ZrYqpw9yJRxYG02kOMu5jkDbFv3
acslOYJCCfc90UalnFjupOER2IIUVjc5nNjIEstsmXqixIn7sLoo0MkZOPa7TJuA
1jhyHLRqC4wDyYfu8uT0LNEQKzXiNZFU104AWLxcrEPu+s7RHy3qV8xHjkqCg8bT
mCOM9YB5GpcDH/Ptn43RMrTQC10S8jmWnQ2qKmNt3tMGbSa+HsiJMOOxTdxV6bcV
DrptGg+DCTlwG3BLoexsQJLTjMEDUTUlQgfq7676jpUfMcm/qlhYm/Dksa10nVad
K/w6mxRd+lhtfpVHNFPmeUfjbvhTabNUygNrXQ6wBXDPpN5VlOrcunugMyWYZqKI
o4Ji+D9WnZ79oy5Pm35Sag3iTM0BkyNSC1Ap4A9OXirPEUlRLxO70RQzS7n9Vz9K
GlS5AJDHTpLhdRfGK8VOUBGYxerdkMCda9GJFaa2ZxAmTZ0XVkHFwmzArVWkmtPC
zcweM/LFHwCBbvUW10zXEZVFE7EmWXOSXMdZPWlu3EvDjjJQWBPOTj/xrGzs+8z4
BomMK8a5La1lQ7wO//wF8xIjWiX7W/X/b+kLEJBTw9apUEEZMQVgVO2KzdyZjUlK
5Krbw+Wds0PjtdpkVD1qi6KDYe4AFGT5T2KaRzQ8H92GOE2C+UqUq+wiTPAtsg5C
h0vg5huG/w93a0pouWDx/wElk8p9lrV6dCt83sHAk3cl0Hf32TT6NjAaRZZ4mOac
QVd7E0+D1p+3YivLbsQSMzzCWg2elqrlccsfogRTbJ1M4lAhkNEwRHdCh85t8VJt
w8r3Q87DrX8rlyZGt4fBmzzMoJw+mAwD1W5HoFwaYbEBlY/fLm6jP5jJh2AXLPqI
lHxJKL6WWNYn1oLaCW9SMVluLQDSvhTAo85Bit7Xv4DoKEnF4I4vtR04Vy3ln2Xe
6eZI1H5P5p6UC1Fe6S9etZ2yWkehvTDXpHrQ9Q0SXH+fzAmcnnu3qSjfPqTjJ0QX
A0GxEzozkFXunuAQCFmn9/51MQRxrCsAHhsm1DVuuyARtH5Rrpv0u25NoQubMDLa
k/86zf1m9/Y+QPd7oYbfVgs3cttNF4O/4BYfjFJWLrGqZxnRhZDwTqG7CySmDr5v
08nWzLdCunUdIzGzCT1l0x8ZSonOhfaWWSY7asoEH99u63ZA89NEWF+5U6pIwrcK
T1YA4IWD3jh926PSOuMcFnuzz3SpHVZG0hGFWktP1Ce9rK7knum1k5H12K8BQvuL
GoXq8qxj7OHp2lXJbJUgpgUcXTD8k/5l1o+7+4ivir9mdJwLTeDUCnNbDt5yCYJ6
YET7PYB/1mBQjc6qG52Nz3jcJSR4QstZHrgZt7D7oA9491zYRPp5AAEKDsdyriLC
54N2v33OBVw2a8v3+8PH7GAwQ0+h+Nq2Zm38c8WTByHylJVj1xJdq+5oWCBA74jW
nt3rDej/LAEEgH9uTnisGAXLh4QmOCDlDFrceHNYfZMo9c6n4SnDOs9e+9OIEBS/
BQlrSbsCBZo8FJIaZFd7+iZQwWtopgUnSttEosFUm/WP/av4PxqgdgF16pYm1o9t
G3BQA7yB1mKN8zCmcpuG/vxLN2EGBG4almX9S+xBIkV8weyfeniKPJqHyTOEXLWe
EIOzBoTyCkImksHygX4MkYleYtnU3H3+BnwfJBVi7KmqPgiJlGHdMC7++2j52jMA
cc/gzspTh0JlPoixsQ9T35k5fEp3FEhxxSL34F+f5tu6j+Aro1eAvfoakhBuWUhT
LalzAew8RIvsiGF18pVJ1us2A+L92NdpEbNz5IGeSrI85s7RTlBUJnnYgdNSsTjn
nn13eIpHt7JcBybrs4w6jqz8lxVDf/9V4G71pa9raY2uqYqm5q3+KqfpoEEs8qPO
/daY49go8Dsa6rn8Xuz+0fUgC2CppOxZuUsOhmbJIffGudG35ezMmnE4xnrHCTH0
5E4zFk4N841RwQml+Qs7V2ND/TyKWammvcajJ/OGBTO81Y4AYOad6NlB+CF+yNzD
1ujHbEafP27uylwKNd0I4i+WxVDgTn9hxncP4JaJgtWKDsvqmAxnAbTRUGwp69Ne
8t5ESUSAPXWwOXHyGpGSOC7c+KC5hnywo/8KkRqqkOY8LNBN2E1T861emBUE+TRj
vHsIx7hDKkx7dEqGuMg7sN8ohQ89t9NmYMYr6KxcZ+wsjrPp9PS9pYIp8kJhM7tr
l/oAms956ZTXOkh5oZRDcthxryyhbnigEPCocGosn+zt16JAaR9ZjTfScgYWVhOC
9EKJbZEKT9zOYKzshsP41krSsQmettmGTj4kQ6fdVQ8bhzRVTVhrurdW/yxEV6uW
rSt810+SRL0/+sjDVK3DruelT3/kwWVwB0qeI5pupt4zzWYu1DxOi5oqHS4tED4u
OXu8YCLOpUhksMjkHxRLNsDPv4GlZZrM/cfI4Hv6S+hGPePIIeDkgz/HbEVt78iV
HUekad48PpQ8uLHqR2+uRALXq/my4pkRBPhG2kXulP4JobCG3keMteB7ktu/o1NF
bKHb03hVTrJiIQBZHkxk8mSmRqthLnkFTyGgyRtb0g0QFsucjQnWPWV33vWH7NCs
63oO9xbD7Wd3g+sO4UQukWUv8yrWv8u3SPUScMev+27BrqiawY7QEWlwAobsD5mB
GQWFmCaqVV8ygPOQybjfHSOjwYTFn9IHbElnEKRybTW3yPX7cYKB7ewHdirhQF6g
5HfG2YieKLpR60alXh2cQxaG4brict+Uf7GnZtI3Dss/v4dvo1RMNW5zoRXEAFGF
IXSSEtL+rfPO5bH5pgkE8GrGuTkALt2qJw5OE9Sz8YWpnt7S96mPSSSdmACUue1w
Lv5jw33IXI1cnjeXj4TJ94y+DtAFQrZmFd48AD03yD2qgn9ssA0sqV0uGdTbK9yk
dFnpc3kstdQPgOL6ztFksjLl93bJwC0aFLCha3ARNlQKrZ0IeUgV3usRJg13e6qf
OcwYKVz3N+HGJi83na95MBhY49cm0kcOsHygG4lmbQiGQ0pUaW2RqQYhDa9dJXdS
0N/QFDjssvp/Wjce8+b85uK2+0PRiUU9ZsRaakE+sWJTU6rnLzBHZz4hqXYUfSJz
+1UT0fXy38Yc9kgfQNI9e92T94t9+woY03/Z1ntycIE6v7Yp2Wr1ipX04rs2SbgK
bR1Dbf+D2OFV2+ZHmFVYCNkORvIJzAjP5iZFoMhuUGblVYgFyWhj3AKmE9bwyiM5
E8EZtezR6mB+bbsM3i4yS8DxdVLdYUo1f0jFJYyhbkDVkDREeFHh6NcD3Uhq5zlR
RXt+u8LLeM940w/5SzfIRCSV+u4bA5uxGZGdc580aE5Zg9M/gVfUdoBBzRrn9Ddl
/X2fltqTNgc/U9rxxs2Eca+S+5nfQY4n42dFfa2gXJrvZaURb8K6GM28YIr+7SLA
xecGT73EfTH0ri44dy6eagH3aIgaqkAH9MMSNoX+gvrbsV8vXE/WHmG3H98p3yDZ
eqiOZbphdWTZDg9BBXB3G8p+AfhV1epuqCKjQk0yxOUxuVvtftD2YaZfqFVH/F77
gnZjpP20q64rJp1/Woz3SxKCPP4NxlDI4+OgncQNezsRqU59fYLcBRWBC0jbuM9d
MIsCCShVTKeUU3/GywRvlIyShJh9KkZ898jKF5P4uOJdfe70M+tB0wlGGCPRFCjB
m9TZLgRUEZqnoAEjFsnq4fg5ki7PIveqQpdnHN98kxYLCrPz04eWiPUkwVDIx66e
fYHUoVkdjPxKO3gYWxJieMci0uUHIzFyOtDu+9Z/flX9P75pktdQNpWgZYod0vH7
7vLkzoIe9kUXpI0mR8i9u6Bjy/HkQXJEGUJFtUHvMgeZR7WQZfZsIbmo5ew+iRKh
R497GIG1XqiOoC0lFEwDGuTN/FynBwoyYx8NKx+UziGN+28ssJrhDbNYcwSjreQu
NjFZaF29SmIR0H2H9DZJUO1gW0vlA6Oh73A/aaHrjwtI+ezhSSLqDBuZGAgWI+KI
BLAmjuGh2nCKVRtdRvOoDR4nSzhU1s7DjdotPNW6dr557L3C2PrNFCDEQm85+BBN
KPZtaxP58p5Eresl66JEM6KdJWGnxle3G3hRzrEDXF6RUaOO9PKCnPU7rut+S/Fi
ax9jD2f2RnFcWaU/MiNNOy+f5p/QqX0fBdgsL9ylDNFN+AHtgTDN1dthlxy2YNC2
0VMkUBafLpuMom+V8uezy/PGt9MVgUTNeQVf2bK38Bn2AK5SVvVp2Ctd8Jvcpxeu
u7FNSHOP/LQpNhT73d/zSWIwRn82Whste9O5S5aaKdQvYOw4gCeyDCqi9USO+xgO
1pxHx/210iRParY7zTSb2AWokiJQBK2lAymTMBbUoJPDhGvjUz2+XS3izmmw7Oc1
NWA6I7SiusxvZRK3R1YF8pURTPM1Jfscy7GnzAYHRRRO3mOJ4or7uX3jeBZ8MLr9
drv8Y6tZEU0qovjpNev1s0AIDRRkaXgI7Oy1kYW8F829ELMK9MF+B/NGNrVcnB2E
Vn2zAZ1yJ2zIrR7oQJbUqXmDyxWZiu1ldET8N7lzrKxj4dPLTiCZOWbwSXA9CAcl
6GZDymxHB2OvarhOkqBnMjw6N9Vb4ALDTrr0GHRXhpniGNnQh1DxQcu1MCTz8jf2
9FX6I5SNiS8uVxlgcuihf9ylh4YzLER38+QyBIQI4E9mbkMl7nuxAjhfHIEceuZy
0wY+PL5PNNzyDDZfm60fDNUembhQljHZsqL/CL/rxLEoXAfqRsaPni+sW0j1WYK9
UCompiPbf/cJGEqhEg3llWWrUD64plNHs3+HrDPFdl9PDkD+HFwFY8BgMuoz4A0K
I081+1WwtsCEnen+tumcf3R2gmRphUtgjN3xcpNGQ2biLqcz9gOGvA2lVyisiaI7
QopWMy8+subAKS7k5zhX9nmwsItpFxoYImKzEKqTwXoaTkbpZB+3Nrah/wvQ2Txl
tNJ4eP8OqS5LDOFdgFZfOhD4yHCekdWRbI5wTBZhl5XvrFFJLRWKjJH6YPlhQg6l
qarimMIXtOiZzADtUDb+V8bS22UgF7T0cltAMp2qiz4bVOeIO0xSk+2NnJGgjJh8
LryWcgmH14l5hLD+SoC+syRQRrhfvJD644S0m5TJaHTPNz5fQEwkzfCJCsPVvBkQ
z7gWEhWcx+WCrHFKMgnajiyp1FbHA7BQ/ZdiOwqcy5guUN0mNve/FCqqNVHNUEvh
jzFlOd08osButok9lEbV4sYWPS3gn6s/kVjQT5905Va8Bg8JcBc0eYzRTC7pb7uV
wDG5dsifKAwjIntwAPO37wWbXjGfrQr9aKmu1eu8iIPIc90g1HtkZYk1iB3Fhm2I
FnCmRQXolYDutYrTSvE1EdOHscUXDHeNdPkIjjsdqUvbiYdHwaWIUNEopDMpvdpq
W+2ylK6LsoVPaRIqD7amH6E90GZmvN+hU7nwXyXjVno8mD7p1mNxrc5vu7U5auat
AXkhEqRw8hpmkrCMqEzBSZ/25c8aCps1dezWr2cx4w5fT89xygta6TUXmLNwgL9l
nDjM8KCawLEwouqRfwV9WICIZlYw5sgpsDVRBTSQZ6KUW+xfETiB1jM0+jfJWyWr
WsXbbn1Q3UPqOBj1yg51PdtWcUlx/bkSC+z5Hlrc2xhiLVAi+9TbDIFZGt+hqvYy
DnGQDVh3K4Fajk1j/iTx0B/Gt7pM9G7PvZ1Q2Kjud07Q4x3HONFzFvnCjYNayqoo
rIQSHmNj5bpkjPsWO9vs4TbzH8QWBIJth/bSXGc+JBhBQf3XxeNO3qwn5v799CHT
MDypBUqj5+OCGxAzF1aeLyiD28zTZw2b3TTaf+uygt6d+hVh0g780UXqJe5cwx8h
ryaNow/kYwWl+zuAOmZaG3ADXlyCosh+h7lHHerCVtues9G87f45udgv6NyR8TKt
wH9wGjIoi6AJhaJWEXJOn3j8WxgF/jjyGJbanwgbLrhnoWMk3rS09wwG4dEbDSfH
6y9F5mWn3y2qE8NPGh3KmFarj6dv5lq3NFPgsgv+iOXcljZHcGYVbmfxfzeVg34p
BLHNzZF2AW8sUe/otqRBJEuYscsnk8zD4d2CAioddX5gAaBx7L6YYwIxMYGckS7F
SuXFnrPG+Csh8xd2guluIxOjtIJqMcZjZ4XHF5G7zl6zsQVySHS9PLN7ONXdUsJ5
eu80Mg1nqDCRHdgDibR0/MAacAtcAP1D8EeIkkjew6U9eUhhcv+xUt4ziPa4HD5F
5S2u3LZlriuWhTqEjQ75AuV14P+vKimPaCcT0wUKgakToUDJ0nIw8hqDPDM63kNO
c0Eqs1YehNqPJGjH4G8Q5E1rdUeEsvUmjLR3Y1syFhpt0epmUzSreFvpXT/z4v/X
PMg7ZSx7QSMbyWDGYIIs9IJDOooImfLfcJV5QkOSSnkiLtkqV1ERk0l5qFtcnV3F
HqVMwyVnXBU7Tel7kzwD6fA2objgU+jujXcAocq0sHj1sd7s3PwKjyZHxvxIs6u7
pLSj5WsBcW7lyvIZpdT8eeBqh/4bOTD9p2rx0ex86j1jHOekHVPR4AAJFUQvH2Ne
b+hrwonO1aMbLua/jO4fAZ89KUiOJDkjGrCXHjiXwrGCH7mgpYKB7G+0Te55KN2+
oQpF/o1Rchp61MKHlYwpRZDEhCQ8NDUZMIGf3uP6Y5y4WVJA24c0tN7nz2w/zXPd
gndDJweLzXSMqVu0KEOSssM08vTb+Ft0LtyUNZVat+4azT7z126WJt3jS92y8ngd
P85Ih1o5axpsP4s0y8elU9bPaEVsYV40cVn3WTbM3idFEzpTDklkKpq4L1PZ2NS+
EJVLm0/GJvdlz47QGM9OPReUrgtnKCwliGgXF188rgD/Kqn+WMMZzJvy9EtsDdlM
Dojv4Tav3khlu/dkbyp5+YhV0taEW2oK+nFSIIYplo1QolTDRoZKRSXh+WRY6nxi
2AYYvMGZyL3GVL6MBa33XCCNiTBfmv5GBXdsCQWXHbeXgbci8CAZu6Z2RNRh2TYS
UZel6uoPz8PbGj+L9du09xBw6wWC/mFX++tODf89LYE2Q66STFNCo+VdPMfcbAdt
i0gx3YfcppQQMRRshK6Xti4/LMBPNDucFtpNi05K1n4=
`protect END_PROTECTED
