`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TAhSAJXmtw2cTGE63QOyqVcH25EDCWKoE6u2SllSGtHosK/PUFaG02kel9vxZPoQ
nMQvVzYTTQD3k9KgNjWUOAfrYPxx7Ehps8SzFGAQOUbhSP4zSTfxffHaaQbMMRpk
iqnHapRkWPYMVMcwr8e30Kxr3FDfc4KW6i+p1YdAo2J8lyaYLl8zYNwa0oM0x8da
6iYIIQSjWOwy/wUI5maNAqPuc79pqlzJANNfxr1Gna5CCdrr07JXkdAg8MuscZ1E
sVfaLmnxH4pzTcOVeYhRcZDt1EXSDbLigdvl9JfWHi3XZEE0vynt9h9ZNy+lDWSx
51uV4pDq2ZZkuRizXbI9vrAVJaHwGWKmYUEU1m5muiiM1Fk9ovzF6tMZub7JLg4k
rfO4RNXubeTvhMvpV/FLMnmRBPU/FQ2FWRrz41fIUJ37bp8e1bxoB2PsTJ+R41ts
wvuXzaJ7dG8sfFntrpDIw6eFEiMdSgrF8KzTjE4NFgOSm2wOE3TwVDW4UFV8MlhE
Ut+GPlyniuS5BYt6RwhZ8U5CGhYr5qepvvKUc52dF4MItNaGNwzFbJ/caHYlTsRf
SlO83v4VwuB3RG1EXvgTYegcs89mLdD905BQqgJplELQVykrxwRlwiIyBqha6HzT
M4ekKjDXfCVBk2DlNdAusiAHgyUtE+wjxrgHdCM1kP0cUlC0C4dxnPmN954TpPpl
yg1majEBqhRHCTurluY88FDtazi69MkwJSzqhN8bXqkc1eZns3cCRxJ+afMV+vI2
h8Dw0lSUa91D6aGqgN5MRNlHD7bYCZS8BuqyaFs2xSkCmLxXu0PG/4nP3KxNwJeL
EZwL6NOgPrtBW6NgdA24HAVr/ygJMjkuth43kLyki1Kpd4Dvvbb/xvZuQeoxE+Rw
sJC0jB6H+7wu1Dewr2vceyp7J+yBM93rGSyLb0lXADgSg/e1E0jCDGyroiw99NrJ
FNghKMkiDyOe0Fp3H3UVC2w4psIQiJ19ZqQ5/x7bmTxRytZtMyYN0pVkmDBd1zA/
MKyh7MTsiByerLs6FA+3cI5tXTPeg1kBSJ3+v10XOWxiuFD0tgsyn9dm8EuiaHtF
zV0GLc3pcTOBlsd238dSQQ6lrdaHFohTF14AmXx4jt5RLD0tVa98Z65Zi4ViJIVX
DZ5KhXRqQS351p3zMyp3LK8heeKOG9bzZIdxYeSZhvNYluEzmUIyZHx9FdZepNpA
hbd7OXnFZCVE5zi1CySp+dGMCKqIBY1C7vLM/rubIp5SesF7vQp1L4dBm+6ivDXr
PPq7MM9GAUbTWLkM1LGHibr9um2SxjseaS/1mUp3KaiYQXRFzbCHWycl/MdWYN1i
QScn6/cRCpf1eWhhge6TAS7pjeKbHJs2us9RzEZzhKYZ93krmPUEbVhap7qN1hPM
hHt6R00pUxeOD5fY4rwW93TjKkHbdJuIkQTXkFhCH8cZs3OPjBozOP5HtBVzhz77
4Dg1hmyJOUNSckl9eJRiQpERAcNG3Ec3A6/+vSf8ajTelNMHML96TlQaXmF13+tq
g8/BVYALORnndPZXF5kOoMyN6Gz3hrScVaMaUS/tqJrBCIEpNnM/uev4Zi0XG3fK
9Q8TwzAa2ifE/cIF9t7w/0E0sBjBCGZANACUTgGh44SoIPhmk7GccD5HkVvG4QOp
lPIG76TzMF5MNru9IDbyjgwl1XzJ+lV4/NzKiomo7dCwFaibKduAWCK4SODF1qhZ
qonjchLV+l4KNpWyLGUg8uU7Za/+qhAB7a0s6lhp9Jr2UEIrDFXoPJSxcXQHkY46
93W12xGov9ypsZmLekRFOPgtTM86ne+FPVEMQVvgvYy+ddEiDnQ2UGVTnR4HHX+/
0PTsB5l3TdUb5IC8Xp0vJGkTmTmV+XN7roPZ3N6MAwUbPzuILAAqRBFxHasO6vU1
X9827Nxt+WerXQ38e2DLXNeZcpzOUHDwqkr9dLl0v+ad2oVMpH6VqwkXAiepnDTd
qBa9GIBClRxMixYOHFmf1Zk0WKkHWaG35ihnERVjuT4Y7gHfdoupscnjR8LCiABZ
zr0/er4YoGqtKA32xPFJrLGdD5CSL49KBEvmv6JRIgUA5cdDMupXmawXkNE4hKvM
YPKoWYUAgjLMUCkiEWbbL2zkWXjOX0p589DsElvq2OQsV7R4POjc3YZb2aPWKCFo
z/m7QiTQBFNS1z5m4iHaMeXnduIFQtO/HM20DiK0k+EP2cQMOESlpUq2BRiuYmlJ
RUcReVbqtBadRFX/c6IhLddZmWxnnkrYcCAExzRnqnSdpq7S5GQ/SS2mj2foSXC3
SKMf4JGTyuEOUft5T0enzU/AhDJbKPOl8lxEKN+wMmTQR3xADUtbPSLekQu4pUg6
PwiDo88ftMGdYvM249d5wzzBi15hvbregrLUH/stSLCRTL3pbDbcGxAjLEnektOI
cRiiira0OD/ch6efZyz42xi92k0AbXTVSYaFfZMvampkwRO/cWtlxfDft4RdWx+5
mChNgF1yyYgH4rDDlWJtuC1qAGBf6kb5MgDPzR4wdCOlfz09t3WUVEnfCYm6YJ3G
n0dxC4JHZSgOxKcps4l0M3l5lIz/b0PiyzYw3FI48BsWRSEYv+SCDtz/UJwUSweG
UUN/6ggqAmdalEVFmGmElUyzlxp80FByzmMN+2gkw/E9zgic0OQ/K/iJFAe9JCj0
pRWrnjlv84ZyIY7nWb4B2uMor6Sbj/rMM1RruPbITmcMI+GhlBVaHRyupzsX3Ybe
8/I6v/+sS8wRj+0cyFFvOaTLfC2KAMWqmPrAcCLwSeUxIBgPXRJxs3r6KFDwCVAj
RcxNY7+i5cv7fKpxrnJAcU3/VXrj3kn/mt+ozgLYK2gNjayrcTxJ9kJXjdy4csJO
w5TLKGxnwY0GBln4BTc82bl2wa5BtGZS26LwTBxi8XMIOTJ/zhKRCBz/WeaN1jjM
Ej8atw305iU93zKGA7Uf2XCJL8LAQIaQYHsa8JLJoBQnPjrQomVOmqLIvNb+s/7O
qIT/bgujUOQfGCLEErQouSdfrOIEFdQY29m6Tusm2LViXXEI2yQaeiFljV3lCyQB
kzdcdHFHLcHRdzfQOAs1vpQO5OqsMbEDRI8I/6/nAPlzjj4KbJNDrNID+X8fqRg9
tOCHV9e2VsjTVw0lSQjFeuyZUWxjM7n1D/RzMKAMtG+jnQxcP9bGAPixblZE/o40
Fdt5tXG6pUf9wD1NywPvIzX2S6YQN1Y1ufo8sMjgNpnyeDSgW95TDUVtC5+ufmki
nhgstPxfem/wMmRbBrIR00tguUuoRokofIH78HS4+PSbMc+TuLqM56fxhtZ65K0L
Oj5q/DMa+zFq4cxE4KQhNO7IqRdkv+AO50YJyJk8HAUG9Io2SEn89MMQfuuLg4MV
Y88a3uW5sEEA+sjikDZtlag4VP1IpX6b8Puo/F+c5090SHS58f1Qg1v1gVyIvjaw
2GfCRUXyZBoK9PrhNcfMf3m4zSv3K52o90songloirBIVQAOgBnfB7r32KOZN5/O
RVGxDp7/RVLOM4bh6ahZmvyxRsbJCafXpe53R3auhgNdKZLm8sn+rFPTGtTzqTrM
tyV3oWt/7YQieIGUEIM8aBJ5h7fYaYF3VTbyjiAlenluPNDw4AnRR1TQ6oyzi7HX
F1kMMR8xPrsos6BDoUx9dt/efVmbfpq77e/fd8nae3F/c4I7OM6ofwCXh2JX+tqB
qq+fyzMhfJ+/a4vSFGhz9T1kfrzvy0LaQzXCOAsCCvlU8pMJ44R45Kojg7q72olp
JhSTT/H0osnkIbYIr63BtCZ2SzUAi7oT8mlixxCI+nucNYTZULLgNV6pXEWtZZ0T
Jx8wd7i+OKjHf6o2j8F6jKmzvkYLd11VezueFzUNYkE/FR+BB1cSQwlJTHTEzrMM
GcDXpVUCJH3b4YwFgG4/1OsdQvy1iEdLFkzvUzTwwNFEmzSK2aGIMekIBdIAab/B
VPa0vNl9HJdtOJeLVw1AIObjWjHpjI40mOLkrUk/oAYf33m6Y0vJ6VcsEnJN3L2p
w3UN7tIDFkM2fRKhKHcghugWAywEi1jrMQQguPYT0BIJKQne7MW4yhgCSvl5K3yx
4mjamr7J/X7mf4PAQeqTroiI875qC4NznxoTHERPtIz1vMeS40gvW04z2aL8wVhB
kuVyz69YXFArhyCQpyTFwWQvQieIGwwi/RjNhbL0gGVzNlKng5N9DQjp3n1cnphF
MVQhS5TU+PzbmWYZtV+0X3u/W4JVVt35gn5hRA8Ury8p89MHnupYcoQB77jmWBlG
qAUGOaKzvvHlvieMW94JmjGw6ylUcOEYIP2Z4iYQQjX7iUCV3DKkphLq7VLPjEG0
U5agjJkw9b3gip3WLjx+RYijuFvg+1sC2872+6h/mC6U/+KWr17poRz2D482MBp2
WYqW7/Pri7EHEZM+22I341YJUce2WReb/P4eS52fBbf09FrFctjj4hqAicnq6owW
KV9S4jc6tVhlfASfTMuE6ytRECOUfZGB4BIL5lFAFT1h5c84ZpFt9Qvuv3lSF3gK
/BKiGWo5Dhf4Ha7Eeaa4UfeXDoRo2bWAemedL6Ip2Tzi8PoWAU1ak8/fxy45kBpK
bSp9oF/0QjG/KAN8MdTYULjaJURxvh2K6ME77+5nbknxxBGJbty0D0npQLlJdYcd
C+dBJ7lRqbnWK6Cto83Ng4ecqFJ2onuU3Dvh8DrdZJrykUonXG7Ksvgouf11VixR
FsIwQ4QTM8gA81Sf9egJ460Imnq+Eg5+JEkYzcz7tGWULIQv3t/AYRQOBaUEraZ7
v1LgVfdrVgBzKvwy/QS6ncR5JTiT94SJSh0NCFMolVu7a7HOvNhH0SSenHgvZQ2y
SnN/UNHW3bY8/5phvSy3k04Db36zvKzjWeRJIzwcLyTbZUDXogbq0Y7QAQnd4yn4
4w1zjrFYTtlZAJkeWcvt1zzEPHFgqC66c1810U5xbXDt2I1Wfw3+XblEWyjXIE4H
yJQJPSHm9NRANCsOT3+z41yLIiLYpo6wlAlFn32papDrxHTmUez1HvYbyJTM0jZX
GCsPW02xRDfHF2YQWDyw6hQNE9w6PGMM8uUNbvkN4bEKtzqj96kCUJdg04z9PtLr
jtoLnLOspgPouv81QG0oWIlulcPLd/StmZFNOAHZJtMoJIhG31208vPWcW/Q5JGf
svmWpdRIJSVQyyIkyE32Cj01CEcrJJEqrksLeF2el7+NrIMEaG128gXTsKHhS71f
ETV7XwFu0nOIHt0F3SXLQB6WjHTyxWeWBlADip1Ewo9N65rn4JB+fZw8ErF23/cO
ix/J8kEC3KKa1G0rHj5gu7pdz63TzDF68SrKsCYv5/FAJSFrkz6k1wixAsovSyfT
sVTM1B8yLUwNTnlywU0oVjmiPp1vAjJMQoKPPLN3r4xNlTtajcEj4KUEa8/0+oFt
ktWUQBih6wmzt9I7r9O/4vgQhDmgTXB9vvlXjneK3GSTVMous3cUWgSXUpY2Mt5u
EUq3xolTI9tu0mz/gA+7QeWRAweCir9uFntcgLqMm3vlQvTLAMACLJ13Yeo65hLP
WyxFBO5ZEyilEGTx/NBnY2C6dtjxx6QQVpBYCbHCtlY3fW08cuifAfBEWoLRg+aW
k+mhJIBwGVaKwCKE6kX2nlU1J9E8Tv062oJsYchQudccxl1UFVs1/yv0fzngCnU2
sVR6QUDvDhwANeDsBsXy6W8lqCUlIiLC8SGKovB0yMM6khXm8h2h+X7YhZ/J4bz9
A3VvIgcXkTHDeIM84OLWC0nrDNH9bPwi5+KiQNPlKMIfpuTAMKUSg6L1RBnkBoWF
Cd1G7YD3lGnv9J+EBBBq85V09cML96skppkTw+44wdJvZMmOJ0gp1z8mUGU3bJrZ
2Jc0LHhMWqti0d+Nyw4B48mgYexTRyDqRNIDw9Pa1D6Ab8BDWZz3uRkLePZrOHVt
FeT0F4Di+sjtKcs1HgSN/9pQmyqPyJYqTzBeJpYN6AxWdWt5m0wL88XRLaMG2nVD
HOg5FGBpVM5W/UNwvQ0r1TEFLaBbrqs2CqgasrXzIZsu3Wns9NRz4IKTF81Xiztt
w6OD54i6/cW2JMYo5Z1XwONhRieTg3tXIUu+iT4A2Ndbjk8JZUvvgO5GgY9EvBnh
/CbqjjaLxhSTf3uuhLLxi6daEzFMw7gMM5Z+nzJY50zMLA0Qyk+0asFZDjCw3XdI
AdcQ+grFIjUf1lUP7ALksIABEHZwxYyfdvpWT85cevfYZuU1Ta8FhiTRvvgdND+G
fekJmg8MDZLHoYJ8VTgr+DZK61pjELoskx0nI0y4kF8yUjCGNzkDk04Xkw486/hT
om8jUjG2IvliSREvDqfgBr3mCX1uB/LBEond1u+OGfm15PmoErXWDxF9TG+5b/v4
k0omE6E8dI+YcxUptbEN8KvTDYvnYdiUUzH0LmMT/oIz7FXBP0oGwDb8d/8Jwbgr
7LTdz2wg/4gybwhzMhJREdCl9id+W/59xCxPGl8pejkCYAo0SUTRvNEumFaYZcVg
1TF2J3/3l34+9cIZXXezjudESt8rNYBWvGbBQelzqYYVowz7dBROH7yxemh8ulP5
0uPYN4U4tM2T+zlLWE2uZ9UHWB05UFVwVmsb4pX5SEMqT7QWgcmhvr7VpL/btXeW
tdAYhNbC5B5Z74GyJ0/ZEqv6AeR/V8ip92IRFUn9zjWLywgrXbaMbsHLHfuaB8m2
8121Ta5TIJLbgrS++m9Ubbkg0VeilodEogEMoFdg4hYeVWBQKzpaWbdw7r2BD1MA
dkJVO1EFIMSxZ4wHVIcDpzO20KlZycYGKlNP/Mh8llC6hv/vpuL5msRIQjoguUuP
JQRZlxoP8KaLozLfmWiSU70Neza49asJQ5hI36kzejX7+389iREBFAlQQWHWqfyw
xbTMiN4/9KJ4RoiLd00WncjNZoqu0kN63kfQ474IsHp1bB5uJZZ4y+MS8Bm+OKpm
x5VA3MwZCPwpdBN6Sg2DDji9+P8PeoXoYFZ4eIyipuiVH4on8Y1MBPoHg7TnxAYR
wPP0YBT+jSZazjKPeRehxd0qo0kWupKlWmnAzNFLMTlGpt/m9de83goSpxNRbtrm
c7eIeM7Cl6POkDGiiPpdb27Oa4tntCCTatGniyDGpa2VYowsf2f++XkJYQRcfcH5
t2IiHyu/1KAUjwUSxM526J7ygabOJNEI5Q34zScw1cnQJvXe1lCNxGv4PvfOdtH6
H4zz22tYXsqbx0DHmxwvCLcyTlONeXAvb1rAIek9rH7g6I+AUuvaNgLUfIzuTFSn
kGGylEiM5+HZorQ3eOAQwMr9IA7iUAO6Z4CDJ2Dkdv+iYdw2IxtP2B877TvTIATB
IN7dAkccvC0BLMxSQRmcpc3/AZ6PmEdfDIv0NaIyTxVWPa28ytUOSsD5UfhJc1UK
yfIV9OnREu8+YhqXywPaWoKZCGuu7otP0nVqBXR9M5YbU1FNwmmKZ2Ul9mUNM3XI
jRVA8phdg+VfA6BpkxyWiXXo3KXVCzpa1JI3f5hK1ELDe9zFPCQ7sh/iwtfSKcuB
aKmJ4AdpjN3/Uo4L7RIMYr4MdUQYj2jn3Rpw50UX9Y2BZv4S5Kr25xgwHyj8RZqa
TiCOEYqF67Qq07sBpZ29x98VZItremtZLzgWXQNItOJUcUi7LOYZnFjaxHDJldm6
hJJuOg1kGchCnRSTzZhxtxRwnGOrEHWIfL2MYCV+YnoiuIVcqbZMktJUCqMt0ZUZ
9ulbqbpq36bu+/K2ljWg+YGRaFkCngu8uGR/wYMAzOywYM/kzEpHM3v6Z94BOtoQ
OS6LS1MY8i6uRlBbcblR7BAI10iCJXRAzzGLrtCoUASJKRnSsudfRA1IijzrB5lP
bVaJjtz01jbj2BMuFmOqN/7Z/1B262EkpP1M635kQI1LFc64SVhBaEh9XnhSV99B
hWUmLIlG64quLz1z90heT3wroa99oGP7EjAclmZdayFyVvAvkY426fgmoRce9+7V
8nPtGlwUzTVkRBbFDxPpYR7cIs0tpUZYWNswiNrtTH1CRcr8dyo1/Q7j5JDAfG8k
9GlPMAvvoCB+jIZtme6/eMepd3125fbHqycOtBKjroU/WygOntsdfY2CdbOqgan0
7IKCWddzrHwfbUAiwymqfagVQcEQMKJ+HdFr8jeMaEjfR1u4VkN9tUEmzZpDyQnE
1q/T8mkLn1ANA8UKvcvEHV8527CHdJCPTgCi87eD/PFsxENWaL1w2M4kW7dSMPPw
JDoQWkl+MnGIKup81A+AnWZixrwIHZFrVNS4A7sugeJPQ6eII3IEOiPYPeyO4JS/
AX81mpRtoPQW/rUHl+gPRdMVG66Sc3f4P5oTmO4TrIljC9qWf6F/0UlPYkarfe4O
YksnuFjOMxpDqbueAzLzMaNpgFDgZvBbzAJCU3BpcIHkIkI/h8WbOK5+aI1NM6m3
bpL6+ursOdOo6dikPRZ+TuYp/v04PeujF5JqlhCi/7+K5Sp/AJZ2UpBxkeYWXjCX
P0IU3krH7f8f6fzWNYNCrdXFS4DnlKi3ei0UjvYREMWipDwdAW6e1oKfJHg6W4GF
5Go7bWQA8iGzmf6sX648ZxyR7qiGo0B3voj91meWKfhoVrpFADLwCqi/y1YsY68J
4TQt9bHM2fOG/FX3LlyjnsUzB12JffnxR9tOTcdpEv4eQKaVLE9HrZFfQfD3Ehhp
XP8akHnsP560wnkD15f6Z+DXzJKmgL2YDHwOzZ0AoacEmrBmyxG4grV1OBceZjiG
qeAR36lulMVrR782q5ZEZKLhN7w6v5Srao2c5EnTn5IY+Mdy6/XB4isL0Y7gRCs4
WD9nUaktAqySRipnYE9htS+V0hRIiLOYM073A+ebLPi71LE9EcOs9bHWbiJw3Mnd
NrlNGCbys/i3YEP6rJdsuRAM+4WRkqEKaNl3Gsya7jQgvxjH7yvGvgfd7j9I1q0a
cRyF+bwmO62UasJnK7d+bbHaxSCB4ycqkvur4KUJ9shffllyCd8zJ0kbqe7VLZdq
VqBTPA4BAuDags3ZCoNH/jNl14KsdXG+iQgwuQeJM5f9Lp6YmYp49gY7VnmdZ2/U
Dtrw1KdHqhatLE7cHMPCpsgkRsIaAKNC9IN6gxBT3/FVCQvYm1o1jX9AU0N3Hg07
CffxKLDQdTW+BHmcWlg5kfrUbN5fweQ2K7eE1t0Y0/HD+yaCM4A9lDsAZb7D0r/n
WKpZiQ34kTLLZzGjKVaY7NUGqvbJHgGFfmpuxrgUc9Hflt07GiKwCVTypxz58vd+
cI/F13LgLqjeuIkzhDqfXE7JG6a+ScPXOXTf3TDc3dlLdGwwTgr2FWKs0+sKrLqo
KjpfdBd/gJkax8D91UhEJBJQPYUzt0GpDQhK0WWIqJjvia118LNpzbJR+/lPyPWd
mCrsEzfBmvJfJj3ajRhX0baFgkkl3ddwdohw99Xuw6ltnKSMhd8NsGgClUzBhYXd
UfuuphTAb643XCfqGP8xWnaY+8VvDDlN7Bvlp/yAGhgfyOKY+hMmo4taR0IWfFT4
FH5g+ZJwvoQWuWvAierYxXpatBPoJmXpyGTO1q3hTzqx4+oYyJBV38hKpLhmJ+hQ
1RRkpm4ZcJsyAQU9BrnkoEL2+7QT8D9UQ+yU878EyxFQhBaW42c748Kb0zD2RO5w
AfqRo2dDAlRJxGNcE5Nbf6R9TsS9W/hrYOUD21//iTPSBpXaLzbxsRvTO7shZmGP
1OFqeb8bsQdqAk7Ti08Yy9GW4qzM8AytyO577A9yw1Z+cAfU84PwxNqLLEDRh+AR
vFuoAELgrzXw/TP9RATwf6CF8mnKOqMt8Buv1YyAZ91GhXrWcliEhmWbKOAFp1v2
Qb6V54FEvVENmVyzgA4JU3c2WYxFagKHtfmICxd0qUOyDduXAeHYdp3ucB9Dryo9
soO8RoWqGpVWBXGr+YusnGFfxP5/MYFerxeqW9lOzR2SJz4rniqeyy1gJ6E/uQSB
7vome2f+w42tpIqeq7et5R5UF4VJEUuCVMbYogfG614ZLNCsc8A+Y0Zv30yXvZ4i
9U8P3RCloF0jTJqgxPVYnNazL0BBOZWry/mO9uaT6iXMSggEhv7SFRawjSOdqe1c
WszPaYANl0xe2BQHCrtxW2qij9qWlKOwW1PT79tYZvG3xNzM56jm6T/1ApHdtw/I
8Mzb3sULB6pYMTfaSB9KC3+Gb9v53To0rAN6eKyB8vRLyXUlpg9jtrADvZnuHpMh
RFtFuD6q9VKoi13iS51y0UvvGUERSJb9kGmSx0T0hk/vudDHGmXTbjNzk0dL+m90
kqTsXNE64T+XLk4KN6utLfAUUSy+AhRFULpokzfz2/joNdzchQvk6ZFrapBKmIDS
mDvCAMa/cCpY78ryJls+52+iZvm6dxbzu4Iwx4e6NGVomyHyjvJsiz5w5fIaZk00
++Nl90vwd7lXehtnOR1hgsA06B/4rjuXf9QE3GFjSJmf0/Si97QVYwKM34TO9zgP
f3fIJe7EiTOX0uLGt6lTJXWmfdq1ToArwp0zpZ2Edjh9WFqen0FaUgtsNPYinhTm
xemIcQ/aE3c55EcFA3MezGcvXAT+9wqtz2f5OwuNHGrJ5uvNuK0x7lQe9b1YtC/g
kZZT3Zjk84fIgH7o4kr3U1I/KzFYAlQGNxL/qifa2fRATPGvP9Pnvwqh6s+/zwwy
JeO+TyyACSXp0XIvI5ykONCTwWFnpIXhItB61Vw8PP/+btNZzk3iyPda5e4h+0g2
M16N5MJuuvo7HCJ788v3uSAk/xyGSRtiSWB+6fmUM1IusKTm2vxsT6Rno2ULSPCQ
P3GWxtxaROY5Fcw+1afbtY1E3T1f8FIsmhlxrtLNsYys441zMTRP5m4cZARI/pJ+
fw4dUhy8bN2joJ6WOBbgvTeqWZhFuF+2pFzrhQg8OOASw1YiK0tmgw2nHuTwED00
plj6ZitacSFmboR1yB0lwp+Jh6RhQEvyQvOsNGLZd7ozLFriJ55OccBpI6BqJm+R
znkmYd0/GO/bL3KH43U8CIsvh7e8OaNJ7+GiPZ/eaasVZx5boepjoKb3yLXRUmG2
aoAhCj/0EsyTSOISTojjFYqJD0kEK6llqb2lUO0UEpQ5+QXK8B8K3LIhfHF88ADM
yUC3MHCMST0Xtuqzk1uP0ty/XXdZoNezK1xc0/09E4EoFQK7bO+BtPU216+3HrL8
YmgLWwITI13+pYYzajoS3Ijs2BKpDcqHHzhz4Ujo+PhSI6uP9bBE0OU2I3BU7UJf
Tj86hvOHxtuRa2bevyF+LSBnJg/1FeWBieV4WLpjesRqZqtoXpuku0IHZqHBV1px
kutyVLtZcck4hRNxhlE9xOEPwcXEss9kr37DqdvwdoZG7bNpCReDhk3XnnHchQx2
vRdiuTSdMN/ghCrbwny3zBEUJiiK618NoFKdd4b5zMAMd9JqmYRnZAV9gKUUraBp
Y9ywVCsFNqZUkYnrM0RWrRpE8g74p3ifX/sZEMkSR/b2eHkR4bxgzVFeyOLlg6fN
qXfPwo8yZbmMEBRYaCSF82xZVb48DlpH6b/nRsUTQ3C/D+mnqtgdJJgRhU2IiGu2
a0KbpyFxpVpwCSATeMF3DpDhiujY4Xov7I1oZrLc8sNmJIVdKvcrDKsBk2JotD90
wScdA0OEdN+l6+Ai0jNBEl40Kjs+zys3+94r524w56bhz1oZOdD8BWaoylK7TUea
TNXlk2FJn56sRHp3vz1YzMRf6pnaGZ4MJkug6QoeqECMAQQj8LCnWs+yUz9ZBKEY
WMzFdKz1p9IiNpqT8/UJD2TbznXmSaErKeABz+/R6LqBAAO8FpvEHhPCZlKIorIu
7DmUIMIJz9BIxi+4h5XGFekTu83x8s5njn/zZz5rGlVgYQAybA0t9Toc/Df4wjyV
vUl1cbKu0MvPutaMy/Vh+d2yHiQo3X6hePu2Hm0CZ0evqNyo5WqEW5QHruj9tq7f
iXa2Bbiehox9Pk5Dfc75zvq5CLM2BTCqlkOsXkHyGN0puognU5kp16+mvolQZvix
sR6SZhQQPsRTnsW5oO9050nhJbQ7IsvUDPx59wm6VeBAS1c0fcWQZoMwtDyQMXeo
HINrWYE8EDB7A1b+9JFD4zIURzUIIbui0JIDltDuGYKrYbEdx+GMxTiTs0po/m11
w7yP0Dr6yTDzRRUQlStkpFfngB86b0AZgWJFBn759namssEfHp1cGqEoJ/hL2eow
jEKY9xlF7SLLKfmAVhTM9tsdvjbnPOESVRkTFoxO9xzN3gxKFJTVzZ6nJ3m0SHuI
dQuG+MZJn0IZXZGN9nrfEq5oZqh7HyyBaH+tb5DBaI/UpmZyv0fsmVocXxEmzP6j
PVVvNbjHI+lu1VL8vFXtn7BQyKP8yAbPkZHDTXl02OgwkTDlCD99cdEemydWyzUy
qoxF+BKHA3ulRmo3EucKmLQbMCa3zQNCgdW6rfhVS2pVRNCc3MqYzZyevAhZ9SEe
xYeYfp8JGnmcMS6growPpnx8Rc3vNO6Z9Fb7J5/mG5w5nY3clEEqmjSAIhUw6iPh
aTRHNNfOvsbFKSomqC2dY32tWKNwboXGUwUUEGARiGp/L2r7keWNPtlrC2u2+3B4
PIwb45D7vNq/RntGz/e6In10oCmi+bn6QhabBYSjWkEE03GH+GD2wqg4me9GKCvf
hy+dNkabZ/6FsizJIlABbT10fs20Wubeco2ETE2150WfxHCWhXRoTOInM9kWBBLO
EfcIqSvSuT/zMwGNZ+rhkPTn7oJsts0Eym+KZ5bQCps9gjRS6J4aN+x8jEdXBrlo
YYd+YCvJa1/eT+YkyGLv98E39o2TuZUJGJA8HkBW5lkHQajy8tdgrtyNKHTruz+8
ohMirRYUbIHgroWiIOonIFQKSisKlT1uhrGADiQ6meeX9e7y6CtmNxQRGVWbkKnG
rO3wOoWFom7mQZThS6jNPwzjHaML2BNT2aZZz2OWB0Q+Oyc2n0vysFR8+d542dZ0
1LMs28waxgAgn2tH69AJ3h5N6h1QehtzCkvXXro4HgGQZNtxxAoR0abIZsy8HYj4
4dxnn4SgavTGFDmuhA3mVvrx1ZVbpBbiYhxeu8FwbhY0oWSIUCeUSMMPnBq5cAsj
UdRvnRFYf7Wj6uHmiXaHFNKFjCCJHu3nt7kI6btrwincTddrvaqZl1modkw/gNQG
E8Ne773Dfj4o3LP5iTfvfIx+A3riS9sUyf81ExL4hRHLuqWGuysqeOAXZPkED9ov
GUYRC8BIa8wnJ4/BhC5Ld7hz1IU+Kbp/6OdSBeSGGftULK5ETyM3YrB4mf0ugXxA
wEprB6hmhFhxd0MKdfHee76UUSeqAo8q9UnfKn6c9F4WinEQLnvHjF1bQcUDNEaO
YDlg5/tUazHzvItgESFnLqkBpGUoKk7PtSMKaukxf+qVBEPqt+cJsczsNdgzQRoZ
ZF0Nk2GgKgtGPJB/JHRM1NpN0vcM6/zWhdXjvur1QcofAlsBjE9UuLaYvXaAe1pL
87WaLJKScxK4woOS2GPNZlm/5YApr1UCrv2XGYq3BE3RQNLriHQ/ZAuK7H9UdhA+
s/634WsXpjPqk17zSganEj3fVBwgFg98542RvZ09qAOdC99C3qqUPrUfvFrW1MSy
77aRo/HbhWu+6A1anHfaiJClaF7UUua6EiOn4XAlNCKPiurufHo9PDXGmCOiL9T3
X3cbPDudcNze6P2NYOOoClcNI5rG3iM2JXIiG9O68RbKuxQi/zG0uFDOVNeWZoJj
VjY9GZ+EgzC4fEwbDeX+MpnrX6cwEGna5ZskCiDxZ4G1IrrDGAkZKrDdDK7HZLNy
VqvXBZJLQNA3ONOBcWsdKYP/W7YlDYhtyJHikGDEM5LAj9orq7ifTWUVnZF4/aKX
7OC4/NKimza2LQDpwf6k71H8aHTDuwaZPsMD2l7QABU/wGdJq2CG+cGMAxEBANxb
spniOZqbdQGSEVyGXWUnHl0ND7jTg/esZpdiH6O0RmEpOeTwLfmdmiU4858hgOUc
PUWRLrbDp+qKBmQeWOjjj+ukep1mxBvODNe/eYHxjbOLx4kF1Lpc+5xONxS9vqAO
xL5HDH0Sjb+u0hkOaqMjqJjyCyacrHIv1uQFpOZEKt0apOj9viNy+JDuPj3Uw3CC
BpfZrDiVH8Ig9+YyHDDEzPvSZM+UqVUumfDT42ToS2ynfncYmsqHdWDM5ZqiXESQ
yq/heNpSA18FbzdBYQaBWVCz5VryCFSW2fcnusK1sQaloHtr3FBi36Mqwq0mh3Wd
ylsXnZBIWPMtltNpFpap61d+T6as41ybYyp3XzeRqAoAKfRV7H+HHHZA54UM4Uuf
XwB1L9ogCO3hW42abfheCauuv4BX2kXMsZ4BJH81p7NUBnCQSTNxrz0R4Koz+bLl
wrd0ya37beft+devFVlglPr3GoRmwV6ZetBtagbHk6nISVzBEjiZKw9/Vke8PIpx
8sMYRnM6y3VUTQwKIsq1s3V1nuOJF45NUe5OtHzdbblcTj7u7VA1++yc+dncimnk
48Zg06GW/JvWVrsU+d6vV4xTUx88Rp/g6i8a7KeduvmMpIKWyhfmheZ/fnuiDmR8
n74nq2S1A8Pd1Av3XVBVfbpZdipL/6FF5WvRwWwCLoUuuupg4jq4NEZmxj/TLcWM
AsHyRjbDFg8xD6eGDYR1J09Oy2uJP9ulBDtIdpQy37IKu5Se9Qd26nR7D1ySf3ec
zCxMo8TifvIHJ8AFoHyQLfvZznRV//qq37C+kv7zip03coI8fnO8rIdp9vYDFH5w
+EbQRlupSwdbCOmVsTUZop1hgymrQspgKZEwVMMY7LAyqfgYq9D9JfFoDmnw6Y9v
pNooQcx5cWQLZEu+cEg5Kb2vSJAYdRlwnL4AorHMkIPJL3MGBLI0tf/mJEFbuOIy
5qwsLioNfz2QkyUdqrP3dg1tQF6z7QoMe63gb+3FCMx4TWAA/Q5F1J7O/1TcTVB4
zlwG0xMV5hCyq2Ii4sEsOto0pon6eNB1gP8+/0TJhm30sU97/wYyLOl5uaDV9ZUf
GhGEdrGFMIuTebpSGdLut9XDlrATrb2POSP85aUVgoLe+yVIi2sx1OwE7up0vjSV
d56ERYAGWe5AxXQ+H0kC4O/hZMN+YsXlCeOsvEIeksNW63Q6wpJ4t1M4KE6AhUs+
EFA0CdQZ30xZ+S525sjWAJtDLSasxqHYq0hF1WLRkZ0N6fTYx3YD14Ie66A7KnMK
Ohlp3KkOoKeRAN0+dvkK62JZgyCcUG+65o//GPfBOpZUH/E1bDweQDpfllT83DLA
pHVyqkEtYNrxPs2Wgye2i5oNDWBG3bpQMK3sYJs2otqqmdIecf9Nvvni7dLZyQQg
PQHEpGvI6CI/bHP4ygK9A0YWVVAufIVjboD2P+r5A3N0lWQoXl2HaYBzpoEThcNf
5YVFJa7BGsuy26CiQkFJGU0xHG27YDq2m7jEYwCPCmBEUHa9pymPMFgs4IVpyWqW
i0kYuZ/r57d0Rmm2xqjzwxrH9qDwLaWvNSuGDFsM60xj7KDRtpVEasKM8DNYvzxs
kNoynufGY7xm7iu9n55Z8SppLe7qntO2POZryEqCpULin3cwrvtNZgN3Wd6zTe65
1aVcZU7vM/w6h7T9GfIY1tvNpJuUudXiCpPnRw16IYSSlXH9hrnw80vqhxm67/GM
oWi1TA3khG4DZfhVTLV9KCwpNE8AtGTuNI+Ws9wF3pi/qJk0DluGy3QNbH/spIDR
W4VY0AI/xdbGBdmQO4l/c4fUuXY+e9SE2kz0PkdqLQdgyix/55YEVN1CNzLSKyl2
MkYdN22Vmht0qdzaff/LWc8qqnIWrU/TDhQ5mJobshTKwAsIINDJ5PBE64xCCSNz
UQlG47JaCUcsJBCThYBjCtFW9yCVYtVqpCDg0ub5M64Twm79g93sY6dCuXE3QlIJ
EzVdRXVHMMXTJnKTJuoNRA2G+55tuZzO8rfdl9NzrVab3ILFLo++vXi9VlObmPqc
z+r16RXxXGKpBYm/IN/AvjyfdU9loWBKevPzEiW7xh9AbxBWr6tqXwktB9LX+j6U
cnFOXtRnphXofHdvvOwYxSZiEOheNpyBb8FVMFH8oPBZdEmGbB3r3UTCSFv+xLHq
RicN/3n9rZJct6L9TSk8PMpx89vVT5VLewpNfXcT1p0wpp5O/CswnIZdUnsqqHSL
J64ZkxvKvT1/EThgA/O1PF1+662UYEGfzKcuicTHvA3PLSLJBXWtpmTFc0jta+To
rtL2E7R+0/Xkv4jtw88IDCK3TOawxh/hLkUyvuCB/cc4cpvToTzFlsCgC1dBR7/+
qxLE4jPnwc6upDR7x4nBtumdOpmsfKaBpxTSqkyqC/BD6k2TSqTna444t1jefbfw
gZDTJgQafFBJjR2X0zEzFptJjRKjgz9NOepseBC9Rroi52+rJ5YArSHQtkXpU8zJ
SXWw5uuWErt53JuvAdRdH4UEf9I/S1nfP42PUIoQgDn3tSATB4typhVj0engkmWM
FNi0g8fht4hJwoejvJ4ZRh4THBhx2WBVV6F8M2GxWTZ2tz4MK9uJ3egJKIEKde6N
GoWRfaosMB61xuRZeZBwCpFJGMyCIH5V9Vk82MZt+TYh5hMIKvlMqW6MW8AVkaw4
9aF6HcfBrZY0+HRpPPgPFD2wsh1rKDpajeQA1grwZMlRNmzS259mlGReS4SWoI8S
jFlAgRGjLuLZpwoUgAIw/mYLvswwV0Wu1jAcfiORLdvNSpBqosx4+WwyotwHmNRg
tRkMH/PsvE5ntdqsiVYbfU8pUNwNvVlTDqbVPJtYdUSrBQkElFfi19P7260+ySbu
kURJqLiqa6/L0elbgW81AMFuS0bYvZipPxoo1DqtW8ZLGkSMyBgKfqm6Y6MbRB5l
0FzWhl5JnttAE0XfGVPMKyWM9tJbRLXaOtUtD/uRAfhV8xCq5sq9NhH32n58lH50
Z4OCop66EAO5si4Rqd9zettyoh1mbBV2l6JjZ6FCzc1rze3MYxvHW7OL+CM6+ckg
61u/w2FQVpv4FYQwc1p73Wo5DqjX1+Vmos7igJNqZTxpX0/cK9M0hI0wfIpHWl6C
oSUaiuy6ZQurqpVfYug7of9ElTACnwzbgq7o8DBG8iriZpgIvO8TOe2Ggs9NlnaU
A2w7zyWS35quDaIqAERUid8GuF19geWGXcXewIGtiRcO2ZXSnNZyov5ydSRlWl8I
mIWoTowBCILgKBMQMhqKZnfUac7OlE+PZtHU0gqTrO5D1rOZKeKuRkpEbyZl8SYx
nY3qxJhpfG1OCsxSc0KAw/1AfVG2BbX06IfV3lUIcB9ih7f6ngDsKv/m4LHdUvy9
nC+s00I/F4SvjH/XGIyg6hsfFwR7RGqpUFkPTvyIHUKxyp06Mg113KqABWPlEgrK
+T2buxRpxfUfZPjjvY+GgpYCDOki6IrLtWq0U8fd/tkGfqqVOckTOyjFjpjxPp+I
bMB64Ei4UFj8vP8LWPsako48feKU56jGxBmsGdYDhEhsSj02yz3cc1DoCUXSP87v
EyXsR4Q/FFMmhD7CT+kJKo1/xXFzT36xLNg1EGEU605QjsMQkL9PVkVnHUaxd0dT
tSS4bVObtPLLlIXRngn80oneoeVljpVY/XY1fuBUcD+zGl0MvjFQX8k6TPA6Mjfp
RvT+9oTi7TmbywxxmsRpexBUeTt7WLOs5E3sxXpB2w9m4qyExQXPxa2Yqyd9qupC
PbCQSG+JqNtLOMqGXgCod5SdeV8JRpLX2q6GJbtsL6U48E/087jVuIOYBH0R6gKj
ggUbh4HC4O6X5yh98gRvlrg2z00MAZaqI5xXuIK8VqmytXByWYjBJZgCpNffzXjW
XRnH62hOjnyrq+8BPfsiP9nCcjIfUSLPnMaD8s9TXrn/hRLasbrEXpy/1dQMRgIP
2vo7IvFZH8hIbBRDPQmR9zEEctGfLiqRZpZvmd3tR8KrqqLnpeJa17faUduvPZo7
xEvYl2/cJgXHXeHFkv3w2FpLlKPXLSuS3O/gXApgAsCwGJl1jiShVLfr5qMXzSpS
+n9asgURLNz6K7Gu/QQVm/IdCZSX+UoGQFYzvUqalX52Go5sP9l7BXgSsyPROPFF
MifdyGPgZzQWSIdPsV2I2JXrfbMkvnvnVLZ06KgM84A3D2B0rgnQR/eDrgi86HEf
kh4KUBuh67t8Cw1nzlCt3v0pgIxMqgBfQn1ypHma1i2LTba15W71h0fZkbsa4Wyc
PQl5NIdv9MI1na31H0c/6aYnPto5urrQRFrn8+ZNTBupv3G+43qDhOKZsrhZluGk
SsGRgujRIwotLGV8/ujIncsG1rLgCSHMUnzHzNLECFUdSc8Slor+tiecAyypDz4o
Res8PLMfgFK7PqDmaZTHloiY8sumJN9h/ZaYNSZvgyLTKm4Bsz8KN9QxCW8HLQOy
S8vtfNdrLswTDT4Y2f9qOWDGPYpaqjUlV3W2qf3Ax/FyXnigQtwT53VEv4BWhmzZ
sEkcczFuKO95tVrzTQyzXesuikkp1Bx3cdNgDlimMvZLcfl8kJgTTTV4h6vJL1Ih
N66WogrZU967fR+4KO3KVZI3r0dQOcNLBs6oYNt5d5NhJapwkeoxX4vCf+mgWCdB
E+n29UzYqsCV+dwcybjgCg/kPxrXYlyY9eQ4qHo6JDmhvY4Aac9HCXzVGTUKeFGT
LtbPihG+ap0Cf3574FdoSYe/4aKrqgOoQTn07kJJVsQcN0276JCutQJScp/+DGCh
wHNgIXhJBBqiofPekcUuX9AAmdNjzwCthFF5QzDMuYWH4wz5xlL+PbaYuUJ7Hwe5
AeFhtiuT22tQJlDbw8EYzmbLSTkljo8ApVl0jSI6UGyFwCdD37S9iTbi14ag9uO1
DyOiyDVYHfKurPh9h+kOJx16Y+MgQlL4ss1OXn1i1xODlCj55bBD74pE3kPMcwWU
0l8BZ3lpqtYz+8CE9BFM2Hwavs6BPrUPh0NCPLIsdErudvOyCHqW3vai9YX6bul1
FdR4SHyyBgkjpWehYJLdniHnThDONq23snIPvXiQQGSW1CAvND9eoPWrxyZzfWKj
v5biN28NU+14kOrFKxXZvencqwFPQ6pFXvVeGMMrbiBSsmrywLatR1TGIDldXGRE
XtD7QxmhzCVcOnkG28vog69JLkavXft1ek0Z4WB2LXD+eZo4VySuXbK4Ge0npvMa
ajcYCBcCA7FFetOIHKKLJDUSuI33pMOaK0gVTiHxHmDDjGPvJNlnt8z9mzgOC/ox
647ywTQdAA+bIBOgaOs5ivwbTNwQfMDQsybE5J/WZnJRZ9EmQNvZm2UVDhccz0yL
rTI4ws+EUonmsV4x4qckaGFcnrbJRUcbtp7EL+37F8dw8rg63xilihSGkdQ3Yudz
0ZklASXRbQqnZuCBMi/ivJSUb0TEABzYlJF/ZrTH6aPxz7VWSo+S4SK9gQDri6DX
jRaKn2EXPh5iXtBkPJKkqhSIn3Fr9dAhzBTxmZS8IDFpm9xKmu80Ungi0Y5xhJv0
nzvmqxF6TvhP6KxeSEZT7unf9fCDBowYfncOEXnesxxitKUkkCjt2fZjuYPQYCeo
sd5y+O+vSQDEWovRt760TKcCiZcELA+4qVvyLUccdiBzziOmCtA30cDZiKE7rpsZ
tbn56u+idP/12Z4tjZvB15EmPnSQyBH+IN5ZX1ZXDlajV9CHZsx+wWVjqFQ1smJP
E4RZ0CgkHvl2dWTiWqVtilDvlLpQTq09w/zSKXLbzkcEtcIbYNcjxcrmq56Vozmh
hT1cqS2gAi2Wt2kuh4uY2KaKS6l8qAUuKyS/PAErw07vI4nWmtMY6NYemJY0b9Ck
ISJF+RJTTngBgaDRf6EAs+o4lww3o98G0wRoCLmD3ebBlV+t0j6d3rw7xcm2Jb0V
lwSYkGD9/jP2w0dBuFHeGjw/fOdI8a/ok7n09ZvXYzN4iYH8UelFTi+5oqK/4vbe
FB0NhYvVUzefgCZBndkS0BjQVvVoxT5Kvj7awYHLIYa8i4+F6Gg94fnt0QLSdoOy
yXmY1ASqEs1ItRnTNDoQHVczTiDkVekr0TA9jgSOlI3tZr0e2S2xuKPS1enblPoc
AepxzOJeOOTxWLpYdsWkAOCpig7C9uNZF/wCxBpLvY+TyzxVd3A+PLKPHm+Y3LJ1
md4dmv6ve39GajitsRusg0Otk7RfrW4q974yYSYJjUJMm4rJYk8Ogo6717mlB/Zs
yXgeBmyfoFizpV886V9vZ1daKH3yPu17bARokcYNO/WZYQeRd3D55ExvnNe96tnU
0LN5PKyj7OBbXnO2609vXayGoPKwMDv8WvNeKcFrWHFNNdR4YbVlqnpDQw9kxVFZ
RtpfbVOZOy1S9t+3OmVZOziOT7OMU5Rpz++3ym6KPu84lYU7RG8uD4qVHXTWXjSQ
FFT9tRPzu9SeTD8Djk9/oWl6A8+C1+zNfWiIzLM5fVCD0qqpC1H3WWyZFb5WZYYc
51Hb35iHOzlWeWRdHeGSNkyt9eyDl5cRsVCwej84RQs/m5QN18yKkNQwbpI+D99S
1qnuP2/qka5Ya8IxlEuq0XWTFwnpJH3dKURCN5drOZHngXOeZB8gQmtE5droVRrO
4RHnwOKj9AlmFrbst63+8EIJyCyNDNZDlZtCDZgCmPeSLj07+kAmpYrJiPdR7yYL
C5D3PB1qDDaGk9jgEZ2ZQt0RTFaQV2i+JEY+a/WEOPxGtve6jGMk/R8/EnYPcJOT
2+gmjnLkPlecZRUli4Gwqc8sc5TFr5OhEgZrjJWmARS9RtgyumnBOMn1LP8WIOEw
j8jRgLJNk0zu9/JuNuIUEwk9yV1g+hoExVLvjfQDe/5IP3aGQrcUhMkicJisXrFi
cqUraqRXs77k26uFN0itgxI+VgAd6mFoJwDdjj8Rgwnbq4cZC9T2BX3vv46WhuXS
/QjxbR61KQMIFlwRABiIBlaNaQtxrVN45onApLES/d9PsO4+NzPoJaiQ4TlPZvuf
niiXoLg7ACOGGf+tguBgLo2s7JUu6chR5H2X0x2y9YkqK874JjLRWd/zzJgtQTM/
rae4s6xC2i85n4Fmhr3LirBj8F2tFFvgg7CmRTnWfFRRhIapnEHXsu4X9wpwVSJH
f4x3gcLAY7jIG2UXpYL+KQNo0V08Zq5jr3UoNB+WhJYELPtziqy5PE3IFv7AYbjk
XuvXR060QbNJonR733NEIJ+WGSSUToLqfhJqweUZjEALPMgdaIB+s93pnKLJVbpJ
+w9R9s8LuSEWGTgPvmfZv2wddfhnFSFhwhscBbniUVcC9jfqnMzVdcOiLC8kMXNC
EPl6lJ164vi0MhnayJUYYIK0uX9pEtjfNhbujfi2mmgwmcYeAaxUlQD136fEKZrw
M5b2oIXUCl2dpGaBwNRR3LmNCGJ/WCD+rxim4wHW7cHaFzBg1BAodLWUpR66uakl
cWFwZDnUWeMQiZIOSZXgkb2FJhxEpfhKhDOkWq1mMs7SVaWDv9ojncvNST5dVuR1
/v7KR8xLeydURM9MzDIiTjh9wLB8AP2Fh38tTA8AqUL48CqIzMF8Nuk/jh9S50u2
X5NLS6wLgQoFtSTwO/04XiSIXsv9nE9UZQpVLCcIUqEefAu9nn+Pe/EJ667pvK5Q
Y3fAAj6YtQvxoQdk+9dX75O8Y3aIVy95gFb0ijSQhwXT+MVUh1NaRLnAiHNNvcy+
prco5oNmuP8P6so22bzAZwovKzjlDQByxTPe2JXMrnM1Yy7apfjarv771sABebq9
6Ye6gFg6WmaaUhycFMK2UbJD7+nhF+DHbNdlNZbn6eMmrI1sS9cpq6MzYP7siJmU
wJNLTyB8gH/2w/AVwGqQyiKeryaj3KOtURWmJ7UqqkLEdIoWZIycCaB5sTMTdtm3
A3gAwUS0HyCNASWjDtJ9VCNctpG7kl9ssju33I5Kd59oagASkpM9vWeWEuhmlrhm
0Dj5vILJZFDrJNYHluuZbkPxzo1XxExScnxY/DveHdmXdR1kzW2clt4nlzMng7BZ
vK6YA7/tc0CwECD7rqiWrjr0lcKJfnsmOj12Tpb8ZyDjpzW2F5I5128/Rdl91Zxi
QCjfadgKU2W3BKjibaC7um/V/VB1S2Hg6nCeA8F9DBzxiN6S3y5mfObbrimTZXiv
ZDWnJNcta1O0Moop9l2A6PUZKV9Xn4W0d1FPkdwsk+GtMc8OlGTWfIQEFx1+0J2p
luDFuzgdK+9xNVNmCMjJ78jFMBU7vnPHwxmpwzIJ4YNfh/svetQcp8ddn5/R2zOG
dtUdgK4xib2bQIjmnDH9Sqf7KSVFxX9y+W2/wiYxNPhjf9xLiUvLVl9qipiJuV5t
yl5fbvTHjzTh3q23bb4+HQ7Xm49IQ5/xH6u/GSdq/P5QGVwl2avmluFuH0Vj+MOv
tAu0pY1DF+K4q9OASf16BjrRLDmhlyBOS5WMuE/hZZmAgYdN9xsDz4KAA72gfAqr
G85sBVIJ32H+8bvf6wGDgLXhq8l3Ryb69mM7qVdVsi1mU6qSAdQupKFIgaf0IEjD
9/sXNCLXC6rpw3Z2qMpyBVAOUCSQHqcCCrWxsVyZEZYcoPZ3lhegNMxIt+zTGfW0
Fz8MJdeiPL9mnCegB2Kq6Z7ypC6asim/B+vCukaeHa7R1iFqHtkLoP5dhuBMKiN+
APC96oMsMjfgxrEawNAIBxhInMdf9dyXgeK9E/hvC1uDlSs6Ijgtn/S0WZXCMEJE
VStAR/nOo8QDqDJfjkU/rnvl3o+hoLQr/syZIv0TnSCvInYeAj91DDqqeXN/GudE
RxJRPMfmfT6kob4qDmwCcVATSDkBNTjb+tWM7eGGCgH22gZIxGT/juKts3gcUc76
PgITZUVJvXWioxKXgFU2XRqXeMKDZER3KWpB5FrPSZ09KOiSAC/PR/gX/kmSky9J
rHhC8OAKevhoKDqyAkuo5R0uIU7Af0j7fAgWdxvb5cuT+QArTeXowXWLrY9l0tRA
Fwr+wdTtm7XtZRaTIeq6NxjVpwS9QT0YbQefPEn1uU1sacDVkVEeYBzfdjg9Y+Gb
YPJna4twStPIQ9Auy1J+Tzx79GkM6DFr+W2uu3VLjIFIWMPUKWJPOp1ZflZcCWdk
cysYZRBXQJ9+vcVU5jso0CgAfG/P/Ta79yvzPv48CiUyBv8zPrsliDxHI2sw0FHN
95PjQw3vYhiCX+uA3mvIrR/D6vIo7wP21jr+hE9e2bgPNGHlWLnSUNiNRIUNs5UK
7xQjO9CuO4fm80yDN4R7o+pbthMpzpDDHlP7OeZgfXbKm7TQu2PmjC4r+HlXPcKM
2Es6th7cmEjk9Tb2gThucpuolRIAq9lbjej5BAuToT+/oKM2c8xHTEUQyYgKtsxL
To1i4wuhGl89CrdidYAscdMYRMpbr1IAlnlW38NawaW4ncx7H9meRRb4qoGZdmut
bkaAhXnk5QCyEA/yfehimoh5cvSjGtSnRlNJml5DpPiYkvhvSEFQikz55x4mci4U
HgSFCjgvIktLbN7m6C8h0sKAOXv+Nwb8bj0zICnMCXPeJL0f9/+eHOFNAykgf07p
N2zS/MHkE6cU6VaPIxdzCdRTKuvygHX0TLl2KuY20ccQtfZEhhOdltoI1Vvv0v2P
Id4zEcJQIIPIWinFDIsOKjGEw8rutEI0PJfj45b8MH/vMm9NjwLqdBLEc/gWvC8g
P3OO2m2YEw8dmYVYV9RE61MTV4zzpl0KcZtjs+TecaE+hj+7inlaS48MFKFnDQfF
kkDLhxijvaQMvrmSS/5odv8WTLvDdz61bfcgekfsLm69MGFe+8u2PVTJP/skbXqu
0MHgFsxTMDa3olk3/HEpB6xVA6TdMnpwF+NOQDR1bOI4ORxqbkPmHDyry8rFgB7p
DZnK3eUwnsOks6J4hPru2A1Gdfg54Rm+vLKD8r5cjAogy/rCTavDR/YvOORifq22
pmZoueIsDLr/ua3kU32Z5jdAjGDS0LeabNND79qJsCEgZC+JwlPdw0Xm+3x/RquX
pxcqYb3RB7FtBZJ5IooNBt/o396S/ECBapYMnwtmMyqTKlPvqSEdCQSDC+HRMN2V
ZGg012yBFJKATKP1+bewmxTAmin1JPZi4Em2fbHpd3NaMAxRYJSuUsBDnV5aDeBW
kzDZ8nFcA/4tZg7AZEznORHozAsQBoHbXg/u96tH1q3c37aBAFMDEOThAucsEjDd
45uh/a8g9WhS9iuVTih6aThjQ3tMKoAofODWCk6ONJTefgNbrerDb8Z/H/F7kcHU
Jq624xnldNUvS5n2ztsX7XZt4onXqB72NmbJrjpr4LsabiNWde9ElU/bBty3hoqX
DaatpI+lkKRb6gdPJQj1/70vQb1WBtcqWVOxOk91WNiBdGo2aaE5M9+nbxH1RZOg
R3dGO1QETTyYzarXIIP6uuTOcPyI66WDwknBODDE0QuECftRSAJacuOlOS0aFj1d
5C5TrvNfymUqgrPAgPbScx3PT79j+Hn56BvYo4ZZq+Vh0EeY3pup8fT+Vybw1qT+
MxvBD9kyITaX0TuxVsbBG6hspv/LSGg2RSaH15H7qOI5G8S4IZ+9tcFCZhLvcCNR
EuBwWLqClx47ULt/dPdjM35UiKDe3CYXUFxYfMwqkdeS7bSR3t2jJNwsToRNLznW
lllGPkzhS1CcHudjZXc/4o/0Ld8DP3Ydo8zP1FUdt28IvAV3+oeuhQAMqan4Q9Np
vzbQYRsz+s8NuJYNnQOIByyxTHBFB00JTuaPMaT92V5JbBQL/gWxELasDeQ3xzNO
+XpyVFPxSUC9LPsmgfPTDSYZGJAymQSwZjrxYBBtnUVrdNYp63m8aSAnvX6wR0Qo
4GHpGkYy7Xh84c9/VeZkZ4uTBme8RISgsBxxZ2HspKrVCN4hYPrRBd3ggHVbFCOv
LAqvNI9mptvoP6p27qDFJonXgwrE+5o+phvFCt+sA2kUqep5Jjaq1avJ1FMuVJme
YDhdBVDXidXYqTIxlS3qza6h+hOaRu32aqVdCA+c+JpoDhtSKn/ACoYfWQ8Eqbj8
bTKxuNGZeM7viQ692IhZs64QxFrY/6ls6bmDxMworI6+DLZ689RljbUb3Z6AXuW1
qkDFM75G42w0BQJbX3/N5PiZcRQINhhe4NCtSly0HpZivbSNj8SLtevODROgKqEq
OmSrj5VSS2DgEv9WqwP0PG3PsLXY3AgZ0yxZAN8Z7V0dwCy5G5ui6JOkKbrnWX55
NTuSDs+/QNltfe/zJgEwUJfE+GnlUZmugm5F9bUj32JdSC64AU5EFHn5bnSfIW4R
1+BxmgE0hYyxjLCWbahNpJE5gcFrpLTD4X3bfsSoQxefev2wPxkXlvAkdmVh3/bu
2iRmDX0r95KQOfrmtvG2JOzN8KyP6aCnZosi/vpJ7xsm8veCx3b5Ru0N172j0cz6
KLGBe3o7IB/0lJC4XVCVkc6TAUmDike+N3SNZfA7MaaswBS0WT+ZGIa6TqVRoZPa
QedQs1Ho1vw+gO8+rFAQVJyaGkAp8KRN24RGWhGdut7BWy7YdpWNYUiYHY1K95/D
RKRDVr8dcAJrN36Lzog6d91P/PDTFEUi08rR8GrH0RsAHu5vRlQ0tdZnUQszdYtz
a+qvHQ6QwJ/g125W4HF64lsu6XmZjOnbBvJiOCnl8nTmQZLA+deCmDSjU4Rsnm5y
ykcP8Dxh5sySGaN8GNn5fy90Ni8sXE8FzlOpBvrZ/0xxP95/YvR9UdYgtPC5Bdox
UyOe7slHIyS6vFkJ5eLV2k4TXkx6ewe1gyt070IA+lSHVberIwq+NkMxVk45nQ53
p21pNz4oBckTRr23SgNDrZ1rDtqD8COr0/SqUCj9+gYgYG+YA9KgQ6tFa53i1oBo
8vC2LR53JwNSnRtBM3+ciwKmmq55r8k7ChsSHDnNtTyvmS8PlqZoFyzqiTpYoEil
PlwKttXFRFyV73DzCWnyW5Bs1TcmivXAJct3owheTzVQG0y8mWvOAAop7xq7hYl0
vbb+c2fe31rCMfA+7cZuw1ICvz/EFl164q/4tYnlrMLRGe4h0WrCukZUMwkCQLqA
MLgUgdSuQK/wQjIPe8iLCvrnHfFtOiYq2Xo9MAjCqGisD4jezsY619k/QVQiEotH
hJAmcvJxPkV56llXNojunYnMEoFYLJApfUTv358Ok6LYhz2XdKyzkitk6Jsgh0pt
VokrrE55NJvU6vJduKN70P364l0FGRSGK0i2qUaWKt/d3DiPNRZIaynpPHxe53xs
qQOIoIk8KRPKWn2dqMDiCvQ2e3CzQyMVR7L7BGJo9nLYu7VvIXUFPuPxXlNFb1nB
4S3DoK0UESYErKr8Avw3VWkhaM6QxXN1h9rvx6l9lPyZzq9K/7rIXygh/apxMINN
69/EQNuA6qnvLKNOrFEMULdT8EjQNe/A0fTTA2/1WTygSQGqt4+i01auy2HJ6GPg
cL3r1Vymaz5VvA48SBee1qeCLiAryWsTCdqkAVyEVUvfOzLu1ZuLpgd1FRd10OV+
/EnBNtmTrUe+BZ7G4nhYiz4JfxULBYMXr7Ai8Ay5eN6g5DD7pUQwXLskGR0U640z
dy7QBVD4/IsMD9A38W9URUOxaZi3M44fpOjita2YwnCA6ldpdtKgQ53n1XgJoXXa
0GcAX96t9rx++CXsasN/yAvx+sqQIXDUuh9/nlRFF2Zx8Ei2J971eQ9l1IRNDqBo
9d9OspvevHcHk85WV3FOaRR9yEWTd9tAMhr4QNmsG4mz70Gi/yA2Dm7rpX77qdWn
i/5DbkLbpe6Ja+P716k0JfBi41MOyThUD9dEZO8SpxcMKLIKFeMgazD9IRwI4APs
g045Q+4xW+ZsN9WfcYY1kwVQOc84E2hogY75hrygohVP17UIR6x1TbqONCmAGqvJ
2RQSQvtNbz2w7NBATA1r98fgpufxdy3x6km3xxCu1ZNOeDweazJGUTlBPWuTJb9Z
Oy/BYhEeQMNkE9hlFu8AiQh7N0Ng69MUFtEUBQPsXgC8RY31iBXW3PkqEfavjAcM
jvCXsn5SQKMWlD6YKzEn1CXXtCk6XawoVA/5q2JEdJZSgV1RynrHQkYVA0KN7BEx
fa1g3dp4V9dNKGMYW6cHcX1mI92e6HXftlvrDKbFjlmJTq/Lq7SXF4UNF2raKVyY
sqHuVuIm8n8wK12/snF/YS3X5YkwG7Mgkf+QMRxYDciXdUfWAFhF/HMnw06f2kVV
5OGc+8oPQ1zFAihoXLLzAwEi3elLbF3lc1ByWqsrkxCnsdDHOQykJCzsZPH9GOEt
JoIrXPBCy2SatP8bGOIQiGprOJmiQfIfLmOFl4yY/W1i7AYt/JRE8w6nX3OHVVc9
aqVYjbij3lipMObWAoY4ikN27i+lcqiQLtmRSy2WoLg1Vo6SiGPOotVD29WWx+yV
uwBthPkVTh3SjnsSXgSuzg+DcUnKMSCZ2KDXZxe8Sbe1yV4yCWzRJEhmEQ9Ph9eS
VEYW0LtoJ8luu7lI6x1fxFbPJ8Dfl3RfIDGafp+HWT2ZK40orXomdcmK8kVqXhtb
LjjbmB0LZcRpSnO/WPfauG+ZTn69leQsdgPm+UStGRhKmMNiBy8xcFHWhYE1ESj7
XdH9dYATqBeLIarUdyUeOipbi1tIM9PVAbSYsg3KD9vsy5tSbBFvXqjexYKTb9Dx
dQdaRIeyn609aTnYf1RtjwMiVTTZJ/Cy29BcGNOyRicCE0gfxX+EhPN7xaaPioOP
uC4SyMVLIrR6s7HZ0usG5p0fcxG0HsX9/AV+ikiPVMYfe/qo4KnTxsswhhfCRBLc
i7kwGkI8fffGx7hzvorab5Hn48+5aeBlx2EB+boJSJUKfAD5icAoPJhwIuZedBAE
WkxMu33wa5zJwW0kh3zpg62k50a4glCyF51eZPZAWvQvwvIuwqb9zph33yjQGb77
obgiCCw0L3JbGlpbQPyRUbvTemJrx+HSIwokMjBa4fAK9Bxur1Bt//csWKoRkB+D
36bdpw5DCms0jVmPINi2z/VyJYzl59k9C2lIFoxkFWwdLoJNbFN/U45zXANHJqPv
0HiMLyRTJUV+gMqTz0Rg6q/oMhhs1q/a8yiXsPxr2pWLYwINQdXGOXVNkSY/P8jW
M7E3sAR/H8HxrKl+gOAHYIs2FFKvEH9bDuPd9TCS/IZU/OTP6kpqWuU2JDOffvSG
sWnIcUxo8HDC1GF72CCYmReqj0rAJ6dTabJ4N4jSdLJea4YWTJ0CVWfJ72xMcPCb
o5JARA8Vp9uJuihG1cwau6mB8fg1cR8AEjqHZBMJEA7rQ44RImeXJshOXqYy7Ku+
oTTZlQvZhztIuWMn4rFc2On+uez1tWpWjpXthZeDKDX7IzVzRXegMPtLL/zMmFQk
wBJRVGsaRpuaIKks29YG9p9/YJAtTJ5V10Nz5VOdukB2Nu1gol/wxteNed2VOpRt
7YKLxoUDCT+gOm4192G5yPpLmXoSSqAGJTkNfGek3riiDaTk99CLm3S8WhqXB8TX
PDfX0PnxIFJ9iHJonnkvxmx58JTB/SEnrAOD6muHD5or0MGdaWLE1ylkN1Z8JmG0
D4WjX0uiyjV+Cw3VydmtU5+MmQghy2Mnb7Bq8SfzY83+phnSLIbGHpeP1vBmarQ0
1Rxm76pNYHsVrebyRdBqCA5MPx3swRFppIyJQ0uZGzSBcAXn9+8CxPvrAFV7c69t
s9iua7vOqFizm510g80k/6we+Ouck5Ued+R5/g4w3utw8xBFYZLhEpa4Gzrb161V
UQG0yX2k69E2ob4jOQXB1IzFIDkQMtZK8oRohxxZ2VlytYjBBRskeQTI6CQ8sMxT
Iq76kEmlLjH125/9Ksz2CLueYcMDu8Y1i84VseDe1tDsC10/XgYTJtryO9ejmMnB
AhaiQDk+wJ0NYqcBu7taInqkKtwK57LXI5UzKg6Jb1nKqYvA6ADfR8Jzb/pEhNdA
PPPfvja2IKbL/Rltrm3WFE5f9S/miZH0fcKdQ93lZc1ANdKigncG9Xq6scsLlfUd
fSa3/MDlr9BIgug3MM4DI8VUp69VgMwFF7BQMWKYFcVB4geBYibqybhIsiPZpHSp
dyQ1XJEd09lM/LqoYGvDFATAOcWpuHAJVXSpjl2447sZHIjySqcCILtG5KYSGe9Q
eVoJKSyCA5aAUTNnKtZIGxjJTey7ibAqFvR5UBlKPrr+tGMI5Lb2RWVtbFQ3qPby
nv9Sa57gWmtjrdim5xt8uO9oRFMrFnUQhH9JQGxS3OvSlhOIPUFM26zTQxlI181l
MuiFVbK9Cuj5XWxgHp800PDMkE/4aXSMbVb0VrlkozCOUEEszl7dukv6AiHje7/p
zISoDkA10bySB/JPpERUfuTeZ3SuUZ4dZfrxJK7w9YK6cq0jyOL10haK6WkCUCYr
gDqDWJ6ZDIHYHB2xGyqm0CjzZm7BTEenzpam3bd7r462u1T6CX0FgUsGFWjks20H
18d7my/aSLwco+aWE6z5OJ3dKFPo2cSoRcKUdU3lk1/sVOSslWVAvKic7SlugzpY
h4RitB4bsBTmXSM7IgeVaLnVClbpJccrEE8kIErn9gShwDkZWPmkzFnYktEYgcMY
M8tMMTPQYVh2Mx7g+xs2MjwixxI3yKCOwk8vGNed6oyf++k+iBQHPPaOGrHG6Hhm
soCUbFLNGyTzJLdzJRZ4hGisoSIyEiycvTOlf/aSWZ6rfJeEhcZDAQ5Ii3GcHg9S
UN6e+bex4WfXWQwmUPFa2WZvRjRNgO306q9iWlNmvHi9VxDZnPFh115S+JTPc4TI
5IFMiEdnHjvGXdzK+J5M0BpPIheh4TFoaW7fGvl4Tvf1p3Ub3LOVyP/IA0t/Fego
GaOxxd+RSgaU3zanONAUFQb4aosgNDWBzcC/zjJnMGAKmbDIjF/Ump7sQnv0jGH1
aqcRYRpfqcXz4l8nF7XHOkxLdf0wakU6M2HDe/xCP0tA7dTiqi5oWMJFCw/sAv0j
sXRU/lrVSv49QBG4ee1C4E8WPFY+aoOuKgEw+Qt0ar3IebjHrBRBoeweQJnMr7iQ
GX1zgHf0pdlcZGJ1QnHQBwbRFXf+L1JVJpE7/7MbfveCSjkn4xYvxsabjJZtJ2GM
mwGv6FeGYyqjhj7ySFUKbG9edmybaNhfc4DAQh58DF9S/1zNTTHxKN8tFXQcmyPO
axp6BUbN/UoIymNVYdjIIIw0klbGpTa+nfa2wXiBfrF9NkU1oYPR7OJfh8PQlbER
ECf64O5CbTp6ctm0w0H1A5rTNa3IuqgFPDR/hf1CygIYdsEr/ZIOBC4jzLc46HZK
JYamZ5f2JUWULv6IvcC7//dBDy0FynaAEpXoWrpXFIiCcVZ2JGV7TO4Elm/GABNI
+d59sGK0kt+3ZQeNkrgNuowHQQlLyNE4riqoupH8nQ5GGm7gHLhfgHPgdHj47o35
FutXC7zyl8zQZmBdjywLpW7oVVGGkc4hNm7hMgUNKItWqzGzWMHzJBZm2yvcN9L4
Rs3gxwRl/b2lw8VG8tTUCAZ9SHGwJHeeK5284Lm/4ml3XdCaHCqDvQUxewXi1ADv
fvpTItdxvbBlXuvWBF4lqQpmGqfh5qFXmTbO6yA0K/FR/JRz0B4JzrI9KVulViC2
Cwp0H3hjvmREavCl4Xz/z5bPRKq98tn7Db9jL6bLjd1Kkw7u0BFHbzb7FLQ2tILa
hGmXn3WcHi0Go9bbMHwIIWvV5PZHAzSrr+oW67/Q7ul4jJyeYE6XLEutqlHepwy9
BNSdWXXPvFRkzH8kaE9U5Yeoaz1WV+EnKejUVsdi5iNIJOVkjdCRHVue3PT02Bzr
Pbc/V0flE0oa7zDZVtj2B4OydE1skTm7Ze7FFGDnT4ViUCEvCfwVh0OEFvS8gyid
DIAEO0lz1t4MsYXCTvtM54kUgfj3ZpTqzoLJSUurMoL5IxRivJBQsHnTBQUhJGs2
IUKwWMcoNRK8o0yujQvLa4zXra714UMXrA4HKdp8FpLDe7r3+OofjozWvB6rICsB
yXyxCvmh/wFA1kJ/mHJp4Vp0n7WgX0GjXgRn3TPqeEv+KR4LfYAHxCEr00pKcGy+
xx+52AIcF9pyEflcUaSaxqSMWHkImz2L9fHiQSrQDskpuvjCDyCxFmidgWyDrHFw
Cm03kzEnv1jVfHKHTnVEGujmbYmCVE2L0ONpsVivVd5n9qW/dWJc54Ye1SYl847V
FOq57Y5YHieBCRpB+W2jERd2BWx7lSe0ygllW2WRlJvMdHE79IsUeQ9zT6ATKGYF
myiM6IJgC/0kKTlMTlNnI/pHzoCuZNjDohT96snvjhQbHH6VV0c/ZFL7v5pQoswH
hY3HHzFVPE+x5I8Y/7CEKUOgY+rqrjyHc8owBWX8hr5OSgoG7htfhmajMamiCzXe
lgGOa2kQUnEkCKi2FND/NdXCZYvS/CSspl95o/qJBYP08bYT3+CXB3QYo1gLKMd4
V5AfYY1lrl3dMKuskOKcVHnjkTdX9wKl0S+P0reGBhqGQUBCrgqnFGMvl/gpgy25
QjPVH6J4aNS+nGt4MJZajwSGSa5/9jcEf2xzWppnMcnMu0T1g7CAffJEQxl5P+3N
F66CJYV7FCWJcvV3r6ptPkvPvtVOgpn1Jnv8Zq5GUA7Ah+8hLBN+hDjPx9kWC21p
RJKtEv/9n+c89TVY3jcwKtVWieu6DmrVYPsKM60E6Ds45ndqM7weia6p0fEBZ7/D
wjIvVkszF/+BOcjjLuz/92JvIKWmbVhQRMYPhwejaj2wRCONyqLAemYtRPLV8L/1
dJfYIVYyiwMy7WPurDNynhzWhXNY9evM0llU15fQnSnsz5730uJc12euuF8HpS9l
dEqTnsjjV4e2oKAUGuXDBV3oIOwhxEynhZncturat6RtGwtNJJEcX2i2QvibiSYr
Mos0c06b+0RvG4oF2LRv29rBF7mlmfK8VdPtwLs1akzZyhglnieWNB4Ejg+e8mom
syEKRQL04u+AIeGN11gcPKaYIt6qUriMAMiMdGZc9iymIionmLaEkVxjt18PZnj6
yeeYraK0/5dQw2EDlIoqxpgTLxcb470IPuEwg5rBJtQWUb5RMOkTrz7DdZ3j9C2b
hZgb2RhFnjX567kxG4khDoqYmyQJGSCjubrKJ/gntxjbUrqCjhwxs8ncizRNqPEy
1IfOZTSdur8edzOnpZD59Cx+dJAZ3AgwwY36O7tX3WG9Mm3cE75wJ2ApCJOV3AkC
sJ9c4Kv7tjSwkCD9diIlyHYNAyuqLsKPGpCGpePwjV6wDdN/FwVSCxk+Nfc1aG7V
tkm87DeFbCiDjPfe20vyogoWheEAY/u722dAeQA1oW0KbR/eUxyiqkelGG2qb7RM
qneDJdZpcjzQoaYKc4UiSxWvxomP1CnyRg+JNYxvpV30f7SCbpYfI7dv9LROY8FN
KZueV1l3B7QyVCc1/2fasBpzN/14WgJKM9T3/YphQy46GQkLkGyM65X07lgjTebr
in88O+ZLpxBVPlcIemQCdiKVlWBfydDbPLcmt12/TB3eNCEkwSysHtLyVI2Y1agY
MMttSag0VIN6aWtDQAavylUQzZxgoQt4TyKt8+PsVYcJ2hgolyC2eUed02sxbV8N
YoxgqIiObbc7uf84sCrRhP5aGCXl/qenpzEuuI6QeX5Bv8tu6X7yRbjbsBrkaYQ/
FYGvq9Z3pzzxBa+fZ2AHAx7iKn+gYn8xtDuvhw8LoaXpVb7ArkrF80EYSxfUVW1I
efYsfR+axdcnHWKw9u2cDl9Fz1blKpa5V0LGx3OrKnhb2XAFKm7hry+QyDfWlsHo
GYZUvOhKzG7ygstHGmrj7tXpHZzfCdyEqpPIM+2T8p5zg1BHTaT6tO+tmrxkgCTR
vCVRWtfvXXpOkVP0XgJxAIVXs5GJ6p21SuI9kZ6VVxE9L5ZUiwDSWCj6sIgl9n5d
T3smK39RlIb3+girYrIBSueYgeTjD2Jg9w9796cjHh4AT1egCclJPixCdh9u0DLX
xkEysSuRxExVdh+umUjuNlCoLFB9fT4cnIxkRuXYONgmv/EEyoM173hoNMkTbEH+
rMpMDsKJA4qbyYYolSTIyjFdwPEyxVZ5721+4NOpcyR/f/6haS0NtISGsW3j0vW0
rFtOGZw1dbLIHwk3TzHs7hRfo1RWfzsqCL5XVCSQuhp1LcgTyWsL4APBdKZttPaV
ixjlsKVkNZNpSjPec2JlZGEXZtZZBmbtJK+hLMy01ssiwFUvlWhEYmxrt+dbb8yG
ZFU1w9f4jRnClz0DrTNPL1EODYU74xZLeRXi2Zq9RM8b7Xg8YrvQunhn4YG7de8c
a9kjcX37Ag8q8TUVh35xs/sh76vwsac2a8P+oUaJvWhFU/IJYzBahvgCT+UfRhBa
DD3AQJbyEEe3h02YcfuCjqXkVvHiJLHtkG1O549nR4HKERwJL4aVDxk0ceuN3zwW
eC0I3XmxssvylJCn5GQDrkej+gVKeyxzhd0ybo+FbvSzmkbHvh3+RGwHirgw6fRt
KdJh09Z3YWIbg2aUyVgGSBTIHY2lGTTZT3LE2zfDyDMZpwQJeOrmsKHUIROux6uC
oSZIVfqWRiW8ln8gx+rBTYOr0GXtVxcsDcRCd1eQCxoiOvigvBdaAaxlork2vfZ+
ecROv4L3DAfvWBTSmYZo2C+hZIlijkXcrzlAPREVl5yENwPwwMJqY4DSrNLPfnNp
qQL0axpVuMAO3N9cwLsmZ7w1CWW6VZRxstGplT3phNCgMBgPVYV5xRIS2LJm/eoI
Zo/UoXYdMj2Na88np1b/JTOkVaMsOvxgA4XIhua4K71e+QqcOJDfiJJUuOmv021u
Big+OBgwXbiYjsFeMxI5HEtmxLHaO0X6Ac7xIgKJA2caeTt/4DOLcguaiw2zamNR
nK47J8fpsSQuGA5IUqnpSKcIX9CI5gyN+L/i+oXYe+oA9ZNGZqV7M2JgjaQG8iPh
GDyIFwE/mIXflqkbF8CPg6gTu5mVZEbu4EFVL2VX/Q485XV318j3V3328UKihgGt
60UjjEvJck4gLnQ1VuFBjk6xuFr4E5VEyBFvV8zwlsxLAs6zd/L+w+RnrhyoMBOZ
GxyvLbTKNDiy26z+ipA9UPjqiYMwDOcHEB0AJVxVlMEe0EP8EGB31/XW2c2b92y0
tsCZGyG+A0mMQ/YA88zYb3bF0adS2CJ6Je15+EJfMmRZ+uir+1pMeXxxuv10dt26
AE6/rlhHx6wrEbV+Q01f05Rf29xrqmCy9aMY9RunUOUX3pC+NEvg4NrQtFfyb98U
CRTP0V2I3uwYl/g+J8Asg5rq20T7wlJDn6H7AsLyWN9icUyXbIwGUDUINXhFQLS6
LTYEHB2l0OExb7CLtswFHayNstUJxrw8AgYFbe88kIKI5kRhdqohNxW5jIBqzBRL
YmUtGGcpXUN1zrhglKEt2qVQYFBd/wxP6HfAJ0YvK0ObF3ZpjpgBQ25sJARGwVlz
JEJsZShCULl+gaZVsIhOEjDToTp1Zq7dCfZgWfDJQi8jjCdePYA7UEFOVBeAZFUh
JbDwlq9+nmseB7nSCxR8ZiYFm9cXJfmkc2dXPj9/oOhdJFRhDmv4wKI38FavKLkZ
6TvF0Y7cuIT2TSfAgLVDCKscMCa8Hk/xJyKNupLnWGEsFX93db47KkQHqpH35lfh
rxmCITNSKjczlprwR0f4VH0jSWoOBUVC+ndTm8L0gpZTvCydyq+PsWqk+lQXy+ek
T5JTSx/Lgn2yorCV0pG/pkC+dHQXzP/ye3o+BHZszQTvZyUdrj6WkA7EgnVyaXvP
OQtwjSfUjKRmu7GhOHT6ytR7dW55CYNNzGotsS6QA3Ly1qfsdqgpJWzD0PBhQQBN
mHl7fbRk57scRPj33wCdHorB5d4hTxO7K+HK60wCbSXsR1MsSNSxqcy2o4YEjcvx
zGtqSmBDUT2q+4r78ymxzR/U+/X80qk+CkWwGryY06qnqrmWZMQlQ2hYGo1gBFXi
NfoJMwX5Ux+drKjTWi9d7gDg+jxzOsaODmDrRiBC9MoU36AgPTfWr2eldQ7kgINX
1pEB6mckR3EoPig5A7Yna+aq9b7ekcvycWSp7BHP2ONJGPNErWPX2d8XaKzq1A11
oPbogyqBKhOT2YaJXIRjVJR8mCcuT9rW2pPlcFdV37dslJPy2IZegTZr9R6oBWI1
71LnyFbh4H0+JOnssR+pbR8g2R+vL+2aH7s3iW45OpH3aAY7LRxSA4RfVp2S+3HI
Pc0tueLw6y4F6iDIPv6ATEjn6xPblrpI9YngXm/CGk39sUWkIP6qc2ekHpsvI/Vg
piVgOEPYIJXbrtQJen+8R5EwxS/Jgn+y76vgHHvs4KNdgc4zG/lnYyLd8Mc/V5JO
BsR2KOa3y3n+/+r7e/Gj2BLZRsh7OUxXHWkDmOjNGN+ysTzScLQhD9M9Oy1r7y6z
F0+qB2QMkf1pHrUhTWhZOhGUKn13yRPAm/okSMg7S4qsKEMe23AQIfwjk/2X6yQh
B0jQsJ2nERWK/Crk56w7YEclS0L6Yp8U5Ph40NE+19Y8hxHVaU2Qyc6hsByAVgg7
1qa51EPy9lPgqsOuVCwYQsvg1wcZlg2fpfXq7sqphH6GFopqTGMVI5iAgI4oiprX
J7bIyA9KGmQhrl5phNQSPve7sk9swKHwZbSfZaYsP3ifYYbj8Nba9mBJb6XP0d5w
B0Sa5aXMIqfdW7gHJ6veH/7XxEF6soNxkkfooK1z7iRAb+ijmL59gh+I9bdyOrsM
i/J/2ammMUcVOPEOAAi8aoisJHcELkOLIb6qSzeWR/02gc+xUcfX57Tu2umBzk7/
0vB8lZ7ioK5QyYnlc0reupKlQCHOFDZ2Hgqbv62IR5lFWBdZh1Z8cyXmN5BmeDsL
GtvE7Pl92v//8Im3L9MartYifH39j11RSWau0+n+m1nsOYZoyYGABFCNFA0Gxr8q
dmTj4zV46m0ddin2mXUAcJWdps3/BEEpOS1RjRrhu+dVsfgABfzTTbNA9fEURSYD
cLg6UdHIj7RqAdQRnh4m+oymK7R9w5WVOhvCZNQkI3XBz+2fojXu0koWQVmWCdYa
ulUasASOi8c5WW/CK/R0RBgqHLYWEg+CXREek8Yf9Dz+q4Vp9oGCXcMSnx+Vi/0V
ZvP9zBOTcHqKwTtHdj2RGTb8ug+zEnjjnu82PsTHnyogDhm7oBhRmZdT/CgDnvka
fCeYQHNfVb6AYKynWAjKLmW/dt//PdCNue22DGM/5EBAuWhxM78rd5Cpox4mUyDd
fWR25VJYhHQIOKs8W5KMOoBMF8l2YEyBsOZDaJPATA61Oz8dqj3Gtf0ZJYtyVqdR
Oclx2VdsGO5DEGAegzBk0uSOeaD+MOoreioUlsbuHSaHkEQ1FZm+Uvv5puBN+YxQ
HLGpF1q0ugc1ZC5hTI3II2F9w8mpjmo5FLBYDXECQ0QdER0gZ9tlaYN1mz6/1U8Y
vtT/j0u8PQ5sP8p+7uknIFo2uPYAcggLTgM6ybpJYZ0Xmfb+C/ABrWeKWZl53a0D
KQBCbcFa9Aq/enFVGwqnLPZ11Q9BwHZTj4SLYVO+t8lvxXb/fQ2RdyNJiCrWLlul
2e1F8SF9W2Kb9S5z/nhTPFsGYoobMvBvvHh3yt522aiDOE36qKvPwjKffOVnAj2o
t+Lqp3HIGw0lgp1PWdFzxjZOh91E/GH1tlf1cLJEvLArNUfUlY9OZlOOGpCjOZDw
VU2zfBVhUgzTUUvBcYUBPFDGPuk2u5+O39A/u4aKeu8eelOuEwiZtakSxvautQSo
w60Fn2qrzT7K7sW2u1mWVgxVfPPh7u/OKdeEniyLlzhr+j1eRfKnUvwojsT31WSP
gGjcz2RWei1zcFi1V7KLGdZmfftQH4qeOmw2EhODCOIzlbmqJ+kOM8trLZNvLR0p
7ZU0Pfck2Nb/QdjWTPlqUNxeA0IERGWtYchzDP8ZFtQ6YrS0PgDuZAp2+mG4CmHZ
yIdrKVMtBDsXlkiw3E4nqGft2D1K98ChXG2/K6Kec0eLuBeZDcko1V9ieZcO+exr
byivoNIU5VLgZLaqS+RV2L437arcAnZMfchXuCAphBP0bgtUhGnmUiRsWepGrArM
r0m+OfFt8pOcB51E9QRLauH89RPX3J5HCrhPgmeXkh5gXcnF/JO81V6DSzWv/2y7
7Vu4+BpmWnt2PHwFM0zIOcNnj/CS16NEJqSdEBum3deaJ8vjBzBvYVNLd9s4Cz2f
Ed0gbVeRs1Rb/Clna+s3T6wa5SKhKEXXJvNg0Gue9jtf2oBg195oM8QqLU9dw94h
MdajuI0FC2B2S2w/nTPrwXx2IVMTILv97u/G5+g9z9tkKRvgm9bK4awy9RykQM3o
F4Ac8cakRu42os5DFzFTZEqQZ1izFvqPLIxv/Wk77Z1qH4zyhGD9GqDKuH+iM5mA
uzBnSJl4Pz6xOAITl3WHUnwfcKH3AE/SmUV95we8Y8eFSqfrBz+OOgfeqaC9u61n
NtC4peEaIiMwg5rAcc2p0OJUbx8ZykPeX/HafU4i63kL1YQ1fZorLl9b/pfRMrYm
ShIfJ2AEC2ZwMnaiq6NOUBx5hXSrGMIa7eWVDh9qYFMD2+xD34M+rOg0Sb/rbToQ
NKoXCnxmSRG8rUu+MZfzg6RxpQvdxndROMDgsysmsjg9/eUlPIKZ7tWVAqiA+w+x
9OmR+eOlAl9t/zChuwMv2GwabRIn11bMoqU9S7rls2NmvwmEINioZqsy4eRptSRG
97EKxBfK/UENwwumAOreHavr7K+dXxI5c3f32Gj7u0cR3IABNZ5dV7HlqdRK9dx4
saEGDwyC7sO94QWtrbEdC/+cbRb2kFCYVjCtLXC6QZ8P2cC1Y2GmRJhkM5TySLv8
UVkPocswZ8PI2u+GG1aj9WiEZcvUlF5Rn0xFfDO5dhXm08bFA63zW+6sWLmFOUaJ
D/1go0rzCz+MrbI7BxpAKQWG/CDdE+E1mMkxMucl70XiVsMvAfUul8r9DAnSbnw5
e//CrKEy8jB7500izZsK8tFo6cGXy3JpTG2b4MfQBWx+DCD0nM7c7kTJ/q6e93tA
PGUQT76lSGVNH13bJteSo0Nzsi5IgUoXErQwGzGyQ1WHUr9jsP0Xb3E+7ORrYANy
Y+xRzNN8n5slrxX7gbML6Gy6mLpsjoV5ohquL7Grwvtd8jaE7s30LgESXZ7IOzA7
AMdDdWucMq8iNFiWrXKl7cfGjZxKiESYPJYjtb5vorObhKS8vgugRKQ81rDp/URl
MSJIlMs3VeamZ3fRPlo3vbl+CBSBPnlBdN1f4gI83hc/oIqYeDat1D4UrUvuw18a
RgffPyIdLRdALXJF+sm0lC908mN/5asGby9+Q8tAq0GLoLry6+z7e3LrwLG58j8/
Hg+Hx4xrWOP0vwv/rijGud5xkeWn0JOdH9OveYAx81YoTXO/eCFJ4O5vu/5Y5x5Q
72V2QLPP4KBkuU7jf8ZS3V8cFyD046VY1zpTlZ7B/nmRUKSHkI8EBE7J61e8l05G
q8LB9t/eKmi8BJNaI+6Wvy9L6DuNFjUZpXAgRL47zl5UmH/ZzkjxjuRk4jtCWbc/
GMMKZw2wjbFMVZkqtfIPbb2iE6jH20pjc8FMylX0ipovssbn/VwjDeRMYoE/L/vy
DRoxjBWVqVTu841PM2iCu/BNA1+Ow8YppAKVeIiEtRhV27tlhdoOM1o9vIKPoVAK
Idt5h0uFRbh75QCG1sYDRi5s6hUs2PasecIWEestu3X83baaR0HZVONgusIJu/oq
tHuJeBKJLtu8tKgNcptLfEbuVwBRyplrD2TW7p4Xp4a4wmS3vhUIoOXxyAFL3Vdw
CItey7ilmbH4ev0BpyD+0NMrT0H7Vx0vMj/ZUUSP5rmEO5JHLdQ99LfrJ01eap/+
/F5PR8L+wo/xCvjEnu1zqrqybPTzOvo2xkfSpH6uSaA8eT9LqRhxDP4fnUWPpWZ0
b/JNhtuefW3Gxshw1EtpXhQ1Y4P8W3xOFN/d3yx3EKOYCLCb7T/wrIXBq+uvxNYr
hL4SVq1vxHNNwn3QCmYyhsgXOO7QNBxO1hBpM/S8Wy2R0zUKOp4OBXZ3tlzc7OFG
gD9KGmG9x5pAD9PEYVfixtvmbV3JL6H4uor/I0RDfUIRuHcyVkECsIzFDdujvchf
wyCB95dS1z6rx4tIaT5TdmaMKPMF6rBMJ1pq0Nvm1CujjX13ROssiCDNNappe0U1
9jOwztctjDRjK1loNkdWWVOulAMv2cW1Bq3NwiJyhztMbtYP0IYMYBZ/o7umCn0o
L9S3ct+BST3gX4p+1mu03zWIXgCkBnrjALjc1VPgDbleNGORoLUJnsVxPPGvH3fD
4UTe+BT+dMCFiqX2JpVZjZ3bz6MVi2q5dSN6Mvey7jNT0z1rksYS04MpUB21Zrea
svU1VGxHzN1dHiuu5aPSdsERbE1+ITkesZsYPLIjxEpciCl4pWTiGETuT+RfT6ns
U5BwlJRdXAMb6vJuUHQni8G8fdBQdMEYgeIOnBdi4hBWrKyDWE/gyIODxUEFIbZZ
ITMLByQe2dRatqC09yAxuu317CbNH/YxcuJKExagdcvvQq1CiGx3EP87GPK3NlzY
iIVSdqEUapztgeCPlczL2sUZ9H12U9bzcdf49U5sEjK2+3oOtDuQWAGR4zo7Xuzb
4lp7HdwxxUT7aAWuejbfslwj7F2sBGaS7SBWkwk8H6K7qCbNvwOPWTdRE9OwevoX
LkTkMgvvg+81eC+6wG+m5L+D67TfiHtX2tqPnCsg68zwrXBoeLDHgVGNVSb6kaFL
vwLcDpTNomHRdsbXx6DQGYUGAfzwBF1IAlbo3OPWB1yO3fasGtM3oUeMiSu2Qixo
eRGnLCnoQHARejMT1damsfT8y6PB0krJVn6SPZYavliS8WcqA8ZnZgQSRJSqxc+K
3J/RqgPGibXdhbLL5XW6oISyZSCzHt8RdoTC6boyBsdIzRgSou7goClmyC0yHTaQ
cRHRwRmjRII3FdUCrafv4Q8QZf8W2NDQjz+xZY8i/e/02xXbh2E1ln6fm9JNQE4T
F3/or5/gQD/nFWFvUP1yYGGeguKbm73QUIUFGEr6MUr+f3HISxxhw/Bd3PcqAZlM
qwE+IgGAT4yqdcJZSJSudNlSMlJtP2s5nWE5gU2DxdI8V1ipKyoi8Xwtc0OPoNyd
DXlTgZYiR2M7e9C/FeDwHQMFt6Um5bEB8hrMbvUXYn43OABuXMJ9shlWWhcnENpr
y6vvCmH7uEGiG8VAsOtu5YGw5GGvzbjlOj2VjtgEiBip+xDl17YRYlM7+f3pcIZ/
8VnJiErKp3rlXNjC7b44YJ7QZ6GAL8J+xsroTTxsQJgjiz05YWQD8LlFX1SO1IDJ
nxWaYfLQdGRX31Ytu3OdVJpLF8CfCn/etwf1SowKSiu6/JuNpwYRkytl3DT+82Fi
88RePkfOtNz7bBp0hMVs3Qe8EfOpW0VQJu7MB5g35I+ySrUAyidV//wtF4QAt8R5
hJgswp6OjsmG455pBtAls/lHq3jy4jlnWaJP5JIwRBJoDp8YpKK95LWypHjBbkMm
lOiiznUw/4qJDqSYp1pzK7LIyI6HyMeRNvLlhXcuXxzGOvX0a6zJBk/dF+FIItmh
YB83vfL/+HIDKbBpZ0dGCrXtEKuoftIjGdfY62VVjCzAM+uWjr9MzRLeOLeaEMLX
WWYJ/rRjEziD6Zd1dbOfrtw/2SIUUhuESJcl0VbMNy72c2ByjuAIKHr2Hu0EXZ8d
+T8k0bPSi3PTXgzs1rJUOxuccAWA+ZIzykQKcIh7No8+REmq8oSJZZ7xGhn9IZhr
a4kOD+AiQJeP4g2hMornYxV78IvFQZLKda8YCsTICW9ETgb07qk4ODjuADIbDiDj
mLqAWLtNjwqVZdeIZA9V/YhMy8kDfa6gQWXiyQhUu3zMLUVToU8T/q9vnvduisi7
Dfwzwehp9HO2MsY4UU1zCIvBM65gADF1eg08zU29X92iH2P8iQxgSAteU7jcjZxr
zfK8MH0tlpJqKIa/lSyisAuQa8muUAmgrarm/Uo1NgNNOgNcNoL7dJpVpAvvJYk9
ICRYHzXXNKmYjre6V1ZTLhFeQKSFo5uuY5mFDaBfiANoAvldmMG/588wI8egPcIE
7vq0ameH3ly80Og6a5RmsBJCr0OdGgRebWNKOTfFdFnPxIyWg6jYSJp+cSR3W7RD
wbjXMGQBYISxJmXHoaezzAgTlsIWEvA/6vT9r2Nxs8msVtaLDZ0cw20ejyDGhJcI
1MFH44uFftRBGT4TrEsh68S+vqzFivIR/Kpbypv4lNjH5cR5bWVtyMz540p6SE4x
Nir6HaNUpgSaROrGaLV0xS2qNSCrqcuEX50U9Q+fhC7F0ZMXmzFe+OwJPU2/v0v5
8WzjZtUy1eGuerOGTjL3Vh7xrmvprxl0zk7HQA9baDVH3+DanQbsKpPW/+EpicHB
PGcL9lig1yPRCG4e9XrMBQR37idf8A/mpsYzG08Nysg7X6PTFcRY56RRfo4MgMPZ
vGCsjJPQtQlxZm8RvgT/vdqmaP8399X/vU8c4h3aeOTy1LCmvdLFWpRMKENxH1ic
WNsC5EO2jYGrwjVMKlrdWOUrcqzC6njA7614K6t/ay3ueF2uUFBA5xohOKa5t7X1
5ujcYmquA7p6kQaZzK6k5KnzchfbmsdU4IpzqcPWtNwzhg6jlgR0GbsQziQVLJrs
w607+vJuTUssv1h5yg9pyFk1jTmhOszNcRjf7c5WeRJBD+LhNtFOxClQGEf6HMIe
qJgIV+nW7PV2TutFG9t2wZgTc2nClWsPsGLdCS1rNhjRbnSamXrfSnF6j9NJctPe
wK1lNVR4lauKqxEC+FJdB8PLhGXRzogZGHVutQEwmhZmGruQKMjHWJtd5/pTbkFr
apCCANAUDyOIx1vdcX5BqH3zxmySf8GayLMJqXt8UCygVdwZNuHkGDHb7/TwLi70
LIUlPkfv2SrQAbBAPB55DcOIrOO+XRnY1p/Mako7XxhZFDNYiG+O7Whih63/hEAw
KKGfOTkqJu0OhKel2Yk/1ccuPvUYCRPZRMNO6/OVOSdaWBX9j7PGWd7U7ek8YN/c
zkPvUHEmdKQscunu89CMVU4LndYgs48KDrgIfcEKP7brlDmSpLkqmHu86yFPZlVH
N0I/wUys5RgPvPiNto25RbzVLgNUs+qU87KmcoxOK8i6CrePZ8zvGFqGCHduK3Rk
VEU/rkaLw1opmjrcQWOX2vtQl1lPavoufnpV4hLvzVqdXgvTjIYBR00FMWBZDCKy
pshtpbsATYjnlg2CfUl9VtapG5cl07WrrI6kzcfikyRU1/Mfotz2+fUGFpwRVvzY
/itgdbvUwjgd+2wAcit1aVG13KrOymVs6h5C4gwap7WcrCCZX8kJQw/XheyLzQow
SntKExthemJceVJ8x1d17lv56NMytXf+WQVyexRyTeWvkHTuUheWqsVx7mr3GtA2
emrrPm0ECt5t60m9PjY9i/QjOYWcqUmu/6jKdlupyFfNG1bNSEe87aPDjRRkE68/
Er56J6N31nQy+dAJHRRKTiu5880sv1nB3aYOudlpZtWiwaRibDPXi4z7F0QzOr4z
dX4bgrYiSUk+yf0m/K2joTOeiTw6Hm8HrCxcQxc87u9p+YCbXaim6vCcSjPZzpIj
GWDN/vgnt7/e3JNk1Vb8sGfUc/pIfqpe0iUWGsGZW7GBZyfcQmV5RrgBBjC1nq5O
XDmd+rtnFlTnyHypQdaBwr1raVB42sw+HEWGdPppcqvIDmvDkJ+mLsEEdwdLTu6g
2Et+FvjHwWdzqh88jZ7cenUFxBaVbXEVfjFn9Q/5AYdbOi1jwcltgUWtZL5vxzMY
nU+Tbk1reL/27gq7OcyYybJp82dmhjOz6a+WSsFA/Z68uemkSJQDgtBWVMmda1fE
PaYcWa/NTablrLe0dNjFTejezmT0MgzAHLtsgSmZFkKnu/qoDd9lNxS4q99LlAZA
lAdBLdi1UsrsQ8VhrDNHgtDDyOdAuGuNJnCfZ5vG26bbWd2MxEDm4J0N6LtqhZd7
5XVeQLekw5U77tUdRFG62d74ky2C84b8JgXSvow2/XoSuCcOncDf5dqUUQNkczfx
ANbLDplHE6HJDl+s5TK4AhDIfmP7A05wF8/dRcWrT8+rk6KM1wVUIyNlXUa3pbyM
3BIg0scLS6HAw6VgDQVH15B9zn1cU/S3WU29wvLDg6SBL8xsyfKskGtZ/aVpurbS
dzyo95eoqF3ITAcbHDCOLbj1Ci+VFd5Rlwtfmq1HLAh5EsxDVGqyLxI45piixFf0
F8uOu+vNWBqGdrRTq3mvVzHqeI/AWFhXEWtjgLAHSNn7ytHHj2qFTG6PuSXQCMcv
eCnvpe0YK8T7Cyoy6flJochBgF2C/DkoBtKvyEif3iTrw5GUpd3yH3xw0hrBnrf2
B7GR1bR3uwSVOl0NdWi405O684KyROxjUTFCwBok45otUcFZfGKgv0E34pHWKm8W
sQPvYXyQIGc6+zf1XNvUpbTnDwlsvR50OgfRDaPLdIImkBNAGinirfe8l0kmevOm
iXx7/MO8/3AgcJOwBC6iboO4nCnIsbGidHxYwudjAtY7INeyz5mP6da3dYeM0nR5
9adxFv64erUWFQVYkD9kswt4Mo16JRcekLpEYhj0Rsoc6Px1k25EDa7OQiFVzZvd
MrxVB5qZZXn3iD1A61BiSMTAFeNXAsMwueyTQmWFtXNmgDiPILsXSR7kTwDWKuhV
jZyCch3AmrFDV5lI7Cvyxbii81Y74QSDHGLhlD6SOiX3bFU5AWeYCKh5WQJBPGKe
c/Z6O9kRk7MUFrNJ3HLMi0whPjvc16FYqURnw/yK+mQU1/RDGvbOgqgFah0XgOJC
Jv+LCP2RcsDXXUb7jXaq7DkPyXkGeXJTbaP5idAgGdwIXv5vzk4ruaoIIzEd6gul
AgBhU057guCBbQJIUvSEDNlHtNoIKfYvOvW6vAWPrPLmDEqfY4wrnjlbgiZznsG8
Bq6iPGOpwlzSmXJHtMPIsf7ko+rt6YeCk6I/T477SOKRLfiYoUmIIQuFKye1Nyb6
WT7HApe+UR+TZ9ZUOfSQq1LGEQiAlRPxBEDBLgjxlgdcyTUmmLV2G4eixKj9h5Ia
lhk1mKeHT8Q04ttNRdBQNuPaOpZjZ2Vb8TaQ1/OTGA0Lx4eCH9VNETSgkvmDBk8N
5v5ocZF4+F2n1BtUA13ELQ==
`protect END_PROTECTED
