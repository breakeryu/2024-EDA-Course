`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uz1IfYkY+IOhNb3mqDfQT/Tq27s8F3vwjhmn5sDFpOah21NHsDZTJEHC4Ik4bU6e
TbkQArvfG7Azs6FVbOASOYv6o3G34aO/q+hq2mHWZpgQmjomiNuBYqoDZGkB7GCU
b+WkLPqg1d9iNKSFX1fsmlOcAGaDUppjyBbImfj3h3nEVYk+YLdIvrClFD3ouhq4
TmXvfyZ7GWJBzB3qAbOgYt51cBOIqkCgGVMFmsDV73qG4KnSt0X8MgXmV19TYwct
bjLUlQWMaDwskLpZsiGShfPHVpO+sMgmSc5Hlp22fWe1nA0R1ps0DTUv2yVjy0bW
qwS4sKUwP/hBsxsnp5vi47f8x2cWfVGzetZ4hE0zrvmO6WSO+OX7QGqColBK2ptw
L/YxNt2jnC5l8izejS96SLG6e3/df/X8VA1CFVlnmyehoocpdYsAWF/yDN/OO2oC
ZxgqjYTRdN9QRUBMzUIMy7uTQZSaYcxmAfNRvsNdbYGB3NbiTnfr+YkzDBSpxN2C
4TzUHbhgV017wHGbylDqovEhQotT6zDqoHzltcqUEYpSrAlbKSIBjGtrlZl4SmEn
m8BDqS5yxDY8TCSa++08vp5rwWT2r2a/5rgYwwRGH5aQPXntTN1KSBaYBc60NQiY
qfHnP8SNn6bZq/hHwNL7T9ZWvsQ0lIHS+GREOcIx0y1D67+kQhKO80hoo/t56SJw
zm8DCuNupiY6IwAF2MZJ7u0GSIhL/wdj0gY4W9HKcP+vCT25atsiKt9Lnxmad5NP
bot2dfhAOLSqRPUTwurQIzngpwLyF/SBBUh5tL/GX8iSXQH6+cH58Lp0wpz6p319
Qt5Ba5VD4rvoQONsRxLAAMTW2EQobx6PXcv9uoiUoVE3zlVPQFB0BurhKZg6KCkA
OMyEf8yyvwAOPYbpj/RtEClvscNZVpLpM/yuAf4EgNq2fhLFMWrxYKnzPPNk5bnk
p5Is7dkLTgqAgjOwW+0wpe1t90yRw53zaVA0I3RgLYuRi7DJaw5d21+MYEEb8kNq
bgO/42NAKgALmG8lSwLn/aK0TdG4E7mUs2VV4fGWCzTU90mUinaO7iAB7HQDlfxa
LGab1Ze/onj/4dSXREXTMTkcISy+fVlnsB9CFT+m/8kYhZ1KhV67I96qQNDvF1bP
McWGJL9wWqPjqDduMWjk6J72qis8hOyE8qPnWVF3wkgBVyIcRgwQepDLrS6RICSd
QOHFqJMHRU6Ik9KUm83MG3F9B79yBPF6xX13eeMtCVAaJFI4pQve5HBYEe59UmvB
z1ZoCayo3bTUcINEvWKRO/K1VwGQ5aFy4D1KjF6wZVZmHWZWWX8aRsTN5DxiEGEG
LTjXZ68OkwzvlvpuEqF74HQsHuwztwI9c6wvkSgYv8D21gXdIHJV3VwIIS9vJwon
HUj1t33YG8YE0d08DSvRF1p+OYoqkRHgDHdXXDatvSh6MrT0R535EP9FPiJVDT93
fnDueYU9pM5rkH3lOxBOWhNedL6ikjB6VTRqWJMemBD+9ARD/WjZFNxirHuHlR5X
rUJ115fF1hDizIRfwlYp1vnBg9synVS81TenVFkmYMVKAeMWqY1JLT1CxJyvdryX
uqsYfSBmJyLnl4+lRAVEheJzeITxInPo2Xyhl6LISM8IpXZjsqeLvccaXrVaki0d
mqUW59Q6Di/vpZKTmf1POPQh08BbrZhfvX5QIRXV0s8ykCZ69kx31iMU0iYj7DMx
xrWLFqAOHUjqgIof7LS+aJ/UFfVTS4ovEMgvYKRECPUEi0lm2T+uBtS67+uAh3MV
PljdgJknHlr1VDGA4aW+95v6Tu/nBd4W7PEee8IaaLQgrZq3lCPw9DKlloS+SShY
FbTTaCIv5lBMJlVAWP9ndhA80VfypBrB7X1xfYamqx6Li8faEBIENNrGMq0JrQoY
FpvBBRZbg/XVSKADfic8drH3AFrh8LXdM/h1s2ppjNgHAC+jf3idmdFNJ+NpItjx
3ruvx560Vvf+2KZDH3FVUKw0elqNt17gvTCdT7LmkW2WXiRz+LMCavnHK/Rx6gYk
0vnGAmXNEZrkSwdDQgqBbRmGQ/EymYGsl6TznWvYNdo5dhZPGHsXPUKspoyHxb0Y
4MEG3Q/HNGylLi4EAA9GAP/KDpRZnMx9vY1URsTBU75lU7N5LoQSt16ccZ+807eH
fA91sRaLvtEFlpwHqqUyI4ieU7vwckcZQSw7Jqd7+xM3W+CSsgIlHK3S7FjWn957
Mp+bqfr+BHWtWJAhn5r8QdbeJkG2eO4sb/ziN5tvd4GboGkB/BXA6rxOioBzokq3
y+IJtmEizSdQaQzH5qtsC+nRtbzTOx+V3hQuDgDUa/eDvKHZNyEp/i21JzllZDDb
5NV6hHFLLT8tM2tGu+PFQM2BfdS1XFz+/PD3Q8onHbpO7xSogZpxKgcYr7+jC3Tr
NLVFvObqCHlQKV+TCZcnFPuHbSohb8YfkNG/clBYylDiMSgMP+jp38vpsAdRGDvx
cydCN2eJvlh6I5ofOvQ1XHq8rEZzb5nU62b0EVJxP1aZnj/CFF++p5g5JpCnRxI8
GdTBdo/jQ0gPC8KsbJQqJ6jO3IYso5vXV2j/NB6iRdWtkLjgwGz4IYiNhHXY88Ja
uYahJW2NVRiZ2LZ6knTC9hEpVmazKHkijWPYF6CFtjmmO1vcp+ci8k4/jWvsscQJ
OJ3Ycubwtui6CZRYR0NhRtXEcEpESsFu65oB5MiUH/ezy0gEXkM6tD8xocJftflE
25SGAsxE7Rb6HkVFOIk/pJfK3LjrOi9qASDzjhaic8UoXBvivnsZVcNTDOA9LO9u
P+emafm3t2u3MvK4/InWCI+2n9Wimz38Q52jCyOVjV4nQuTqj/4MGgAKAWhAyS40
DS9mXZWBuhKzIokMWBSO5040MVSUkORXgZC+vjfmV6lm3DjQfCUwsNlEEjKmMEFF
VTiA2Ief1lXBzkQcJv0bqanWZlYInrt/GelP9a3VEGLh4AfJf3Pr/EsAX4miOtdx
RfDGgngi4OwBwAG4hqPPJ5IB9cQvG7AOOnhcXpXSDnpYdspj7MR9BXFSMwKMpulN
+izIEW6x/VSrNmd6Urt0wKtzsPdXuwNkDpkgFiRFkbUGenrdyx4U3MKsD4TfrR9K
YKjgjiFmL+swW0XJ2O6nt8DFU9ra9CiyQqukbyViA3r2szyAVlnctj2HeNo/eZkR
I3WsOuG2KQ3iqVsLZsKjxlOSX2S31kyyC4/N7NDHMUV4mRRpJ52whSgO2rWMrQFl
Z6MJQ55DOlBhPAq+bWc/eB+oVZmc7AnxSps99VcrtT1ehQsXDZDBNFgPbyLWihhz
sUYVzeOm87OMrpyq9Yf5dd50sjBu0hjbcgvHpEVEbntZUvqT8e8yCId1kl/wWp+H
MWCqmMU4lTNZmGrK4DTwvHOwYk6m/4Ql41vN/OZnoJATNu7AMTfnuaIdIV+BAQrZ
AoMhgqCdnOuqJeZP2a3yQcXSN9V9XSv2CB3tQYoMSy44WHjSC3edMuCp0iTFOe/J
AP8bzjyXZR46NGnPWvCy/epUFXxu5/1U3Kw+tJuP92cMbK3wu9s/PHqpU+IYfSoJ
h60PInELXcA+2yuHKVShMLaIZA2CbYv84SzmZlKah9spreRExSbnfO7oCQJey2tu
Gul3LRrYRzdbK6bMWXyvZJNZW7TNYFWgQ0DgyA4DlOKIgLH6vVcXI+nJubUxa3KE
TWuXuNEr6yVP0fw5ARHr2zE5d8r5dQVLebm4WE+h1wxnQIzmWLgFxYMEXLBncAQ8
T1bvr8lbr5F4ytJMmhd9Gbp3Q1cVnB3hSVfrEyTTon9bkXN2pcJoe3CW4bJm3xaZ
1ErAE3U5JidVvpS3tFGK3FokEsE90nRzSBQbWENnxcup0TRaoWkM+wH4JPbJKLR+
FxAZvyGowkqkjKmdEubzULS8KQk9NHM+YZeqjGUbLwOe99XsxS0P5RnhIghzDWLR
8UUrQidxUo5UVfcYMwnQgtUOsZdzg7l7UZPGXWxPEDx+smaArswd90XmpyKeaJGQ
nVu6YAlZnj9yl9xQw2KU/uAHqTn9zCzFb4/BhjFCtC0VVijGK6KGiQOvISZSfbL9
wz5pnNNsJTv6NK61MiTlrRuk9yu7T55pNtRGu45V8/1RJZ4mkT3l2AlYbrWJq+y2
GFG3WNPEPEP0Qe/CoIFpa/v7XnVANTQpIW9uDhVtJfJP/C2bZbQoalnHCj1Lmt4e
ojDQeohwyqWS1KiiJYT7GSdI5/B6U7MHE/0wj1Erec1OaWMvuNk0NkolTgekuzfJ
b3xesVQKIq9lvtpUtDX9WEjHO0HOELE8/O2RTVIyPzDg6AjwkJ7uCSQSqoFCnbXa
xzYX5E+Ul9veEa5If1oIW9PYOvLw92034q5AdObvXYHohUx4hdqF2saEjyaCVC1F
6o/cjug+S9Rx6huNm1zr8b8cBDYHoAbcnzYEfHC6KRjSuuU3DAVEF7+snjk0KQgi
VRneOQbZHizY7Q+/14SnxCAsVs3LU3QShemz2jMoE7gilZQxio5ey4ZSwAr4VnPO
ugovtH/RKMbj4V3mtGvdyh7RmlYBOVKwwrwjhnN+v9K25wuTMlZKNSJF15DDDL//
g8lGWtzYRh0KJKD6K+W8vvSfRo1n8o0lBeipQx6AvLtodYOPvu6EW+pAYclxCn2x
blHgwMvJUyiFSmAY/HbH/2ONFpdkVzXnXTeeXH7CiWg+uSqCWo2agwXP/pQGZWwO
1DvwAUHEOYguBTNxe0XJ8rHSgknB7BGaeDwUuMMVepAU1KEgbqBlBsvOqe2DL+av
AuUuKAyI4aSS+UkGZg5jqJ0AMqWzsiYB304k1gpFTWZNkgPPZt2OQsLJsqtrvQWJ
kuKxn/tbOuF2+mQoeVFaMln5svwMu9hDhwlmfeJNH3ErkUZhZj9j2iVdvxnPHi4W
q/g3wZc8V3WKS06prOe0NvP7wbzZ6yLoWWyuauBhJfLrup/2qJ9YM3NXy5r1XiR5
GvbN3WpFtHTdlJrtRfuOEd1gY7CmVIwaEh7cM+DJms/FBF7ZTryUuSJ0nar3wAir
CuFBE6Aabgv84VP3SAf4jtSSFYi4JhMOj/vDdoNKwK79QN1UpKqttd/XixLh2x6L
vKKIeslv9uCIqNsJtHH50e0g7/aSijrkfgk6iRJwEd5K0TD+RYOK37iuyH2ZWXaI
TMzthyePKwDaI+HwS8SdjvG5XIdGQ+sfYaX3iMlljvF5xPoprpxOPVtaMODHnmbV
dhY/66htVyNw2qg7dTbf1Jipt7ENMXGCklTnmcBdD9FB/YNj4NLqocHgGk72XzdZ
HJObs6lPIWmFyNJcLqWCbORNrb9F7jJVN2W05d81xVvdIrFpZZSTXq5fum99eR4Y
YiGLlvtvmY5Mufl9txCZag28uAM4o93igAgQzYtNvAtISXqEI6Db4LL1uMZXHCRQ
1ZWuMmgQR1irmXpscXEZun5HGbGBLdiLotDoLz/Dl5upntGWBiCVL0iJPUEN9dIe
zdkE3VmTUXebRBH72bcXMjD+I/T7djbHsXYdfVLSP5p+o5rTpOo2EsbYdqDyN+ym
9t/6scozVCLuIcvPnGGh2dThvDSgiUrPkXcdOl8V/W6zqFcCrJ2wKLiDdS2ebia7
f+453NsCqSinOxvOTl9rl9Wi8JQYJELjF8kjy9N0v8IP/OxS49EcpbewZyIJ9gTx
L6ynVZNSv6EKMNEnurs7tZFv31AxXEjAhbeg5NJT9ywD6ouznYs3ih+rWWfoKnsx
3qw989AD5Osy4jALFQ2FpVj6GfbuSdjbyJjnnPVLj6VYZpWU3jGYg7SQ7yq9Ssdf
v/6F1d0w5DvQ9euAeDWVQJoUFEHfys6axU3gK89JIyYr0ABEr0TtmrmLv2sSr59L
aykf9Cf8A/uzdrmeNlm88I1fPQBw+/CQVd/Jv3bAYOCN65vD/HcIxNejmbT5siUZ
s/+QHG3CDz7wAGUFByv/h5o30X9saV0Vsx48sfxkTp+AzwMA4AiLYW5H4IWFbKPM
R7PQ6ABLmVJTnlif3KJjpt7cFnCunBUGIaRBozghilMD7NaT1OcXykSpwk8+T1Cz
hzMeQFXL41ZebazSDOI6M6sk6b9efmQ+2hMJcZYKQWPXFMJX8cjUhw6PUAepqH+8
dUsqKl5XuzdwGqGIX7DYdL3VT9JuS+EW++EQJxY/3tkqK44bY7juqLqbEo7lgaaq
2lkMRykT+ntQq820omtqCeBGTlPSI98JznUJdDV4OyVhNL9TukS+5nyOdv49y8fl
hOQZPRyYDj0L9oAHVE4mZ3CSQkxC6GBegNo5VC0my0drSkDj/SoHg9PzmqMPTexL
cz5iv9LUHUXuJrTMl5dv/q+WRRA5XA6KJ0gcgrewYiGIHe8AfQE88l0w1OOe/IQL
J3XChlc37Z/PvAXUW+83S5CGYp0n8fRYzTfsnZo4UyyKNDQWrQEW1D8UB+dJH1dn
w2xR8IpVDxunQ/Ip+z5FxvUgTgP1I/j2O6dcDYC48ZwiMKAqB0wpTkcnUu9k1g7Q
WUDN74FEer4V2gzL1vGpiTSGeZff4XrFDQeoltj2aJuF9arXrhD4DF6VDMvSgW/Q
JUgDfsiowliNaklLzSp/bL19k4rTzocwZhfstkgpmVcvjE1btbFcrd+z8gMqUndd
KnaEL7WfNCI3DJVnLWDbc+//MgCE/FNS2j8jEY1DztD0v0rpPQuv4mAjfe3C0uxo
iPN+gU8wD+q86m5e706IL4My0Abz29HIkxBQrEslLVAsU+TMm/eh4OWiQltucqY8
7N0Xe2Jo8ltW66pg9NsZ5k/7OOcix5wD4fXIPIybax7QioaLQe27AqL+qIkExECr
fWHXA/e0j9J+H2FdWqTxT5+vGVgZ5BCzHIBgIvuY0kLfmRLBLlbsXZZg1C2hsCmP
ioEmC07NydWU+mybAXUR36iPgJ+cNyBKWpY/z1XnV9o6ppmjh6ZTQERITOy1DvVl
q8EC7O4gvByH4MoJVw8hfUdBg4vxEPLz17zrbxqEg3LdzsWPMo0GZE4fVN4HKmIP
e+4bROwVKqIot/vwyXQRNF1Wc5EaBXATnlAvF76rQNgrXsxWsKZXrh2YZKQmOmK3
TlTcujjnefa6mMb4ekWbRl8UDS4IWgIXXj8TeB7gstEdYr9InrlpbFKH0PbEcCGI
FFGjV57eC0QrLLm65TOBVQajT8g0VSPgW9SFJYZGFiM+Z0unwQ18LgHzVoVkbIT0
zbNLCoZ5hZ+kJuJolqSRGMo/r/c77VND10JOXSUXkGF0Bu+fDMtrgbz/WroGAS7S
Q8zh2eoEn8sXrf5hV/iM9kQlMRR4tKH+5Uo2NTvSCfkoq1n7SIgtfnon8AWq98M2
3eCuetL+SZhUjDBL49TsKAJDXM0jFOEP/55wY7upZkTYVj0MTCpKX+fN4T46foKN
pALTX51TvGPQzL3y4gSyEuHbqt3ZObbTlrVaPEKthDlW/k1g+qav17pDDC94CZ3c
zUrqBP9u/VfXhO+Wujts5GvenXy3/hohfCvAwdqlVLaa4HStVyY3rAGtet5SLwaX
iCc9FQ5V8GEq6ExS3sb8GP6ZIVxQEHlnqWkBTMIgGTumdUduj0o0npBja22Xx3Hy
GTCrw5M5/y3vOuZMVMKYNGhNFS66/Rmb6zNWkkT5yWTITXjOhJfqUZy/aj93AqQS
zvhd2v8QNEvIAI24PX6+cLj/Rya6agr2Bgb/GSoH3l8fm9kD5AZBz62IzAi/ykxB
kr5/SrRO2K4JepLdbFbDpmaCOfwzO8+WBngcEEJ/IRnALiNqoSVaZAkOHsJx3jyn
FDzxkvEGbH8JAsMdMb7VBf9DkfFOG5D9q+OzjgkpgUMD1oQPDm/Z+1X7RMue2QGR
2c2amNEFhdsVcImhF9f1Amnzn4aMaK8ewl66Na1Tt4/QzZ7KNuv4UDhhspVrdZmj
kNnY/hiKBdMhiWRQX8gKUaE9ZnGjFXS09LQtEc9mb90m8NkgmC3ZM/0TT1KLHSVx
l3VKfq51KnKhhjoqtvldd7F8Zeh8j36VM3nswidgle3t1MEHNCXe9Bx7RIHt4tDo
jnJWVH4f8lFWr+K/AkJRP3w7QytLbk3nX2Ep4tfyqDgQ2jAX9Hg/9OQ9tbEhJcY7
YrfT3Tiz5WM+Gc3XXHbBCx44MBa9MDatW9+Q0nIqJe92D1rrcQO/qq15qYxbqErb
m1B/4T/NP/Kmv4ncLlUB5pGc9VhKE+Ja7bPJq7Pn6fHWY4ESTKO8MCNdMN72pZLm
pasFKUtByLjnAQfw7D+Fio14a7k2jIAhOCZ8njlnIQzBObR87bicx7ozJijeA7ES
TJH+lOYW7SMdWup4tZtQ2581W7yjF9wcxW9boPUZl7ypJCFlQ4V28P9zRLrpcorU
6zPhdNacQ6jq46usd4PobY0yDFBpETMxE6Ny8tBd2CSgdJYloLE4HqlicbmM78+4
RugMrlz8yta9ouJEScLJahzqOkzi3qP6tKwj5wsbte+C9e4gfhtS7kRuBKRYGzNL
ZMLRiNMCCnJB3XLbuFyIHFI3DkArtepQckyx9GOy9HkHDsiDpArKb/v3DNEyyKbZ
TAgvl27yD2storp5xURgNCpFTHiKG5tw27+uXAR+KX3Odl2F5xbpQ+OuxC1nlUzD
CAssQqOAw1I+3r5q2qFUm4VY9KoZn3V2G04Jl84B7i9LZU+Pm6OZEYSr/qcQ6z8p
raoDM3YIiJ4pYN7/3uYFaqyivJMQfJ1T+3tS4fKUXJru/fanYOAeYdDtcEWfRvEF
eOajQ0XeACocdXGWa6pN4D0+oQpnyq36x/zjvxWrs8fTOhNa/a4upNPdJi+AP2MR
yiSYur+056B2qpXxYB3Yw5P4NhbXdZH1K4Q+Jar8FFLno6Jwtt/vUJ4bYeEb5vc7
/6Iv8YUUy/2gYm/Hm2l9Qm32Lu23B1RncpN084ocaHNkfWWEnuIA/uSyks09sEzi
WTQgjAJbIwXU3HVegV0mdePDo7OrA5sXVCqixVdC9KmH5RFDki5m5MbEH86vcO6J
lE4Ol1iylCZm3RiHPEc0i2FMOuyX+0I+lsI2W2stiI2BBKUdkEoWHCjVCm0TE851
+q5tsPfXJbM/1aXZ6jT7DGIqvSGfXoF2q9yM3mUG4tUeX46KpYrpmzeq9Kd24nbB
iCC7FVjAo88IhhQP9VYNMLvwpo0Kk6cDf02cKHoTtb0wiZfUt8ejST4HIQ1q20i6
ZYCF1EECSKMSX3G6ybxFNEFs20BJwnHzFOUFNzW0Ylw2P6hZnPkT7KtLgY1m45vS
MB7upEUDsl/Ji3RNNlwUMN+p96mjm2xGET+LUfmjGYQrMmswnrO+DngohD/uNA4d
SrfmpZBBXaquYvZtvQAdbADAo8+DhibhzwsQw1n233fs26uCF8LJVBdY2GO3t3/z
LUwQ7Zorqj/KTsRR1qwM9gfGt/ktFXBg8aX9NmZGsPa70QAOpSGpzzv0/wQIwjMs
TGlIko5bJBpUK4GQLQfZbdKGgPQLzaiwHYrq1swvzVXwFx3QJUOZsjP0DgF5jYdB
CptgXWWrxbvu994glROAVuKbVfjF1F8n5b40mW8VM3XSfmtZksDCJjAFC0jFvVK0
9uRsySCfaaUKFL5OvlHk3ovG8vmpajd4KEAJ4laRraKM1TV8De+FQFlRxu3QTLJ8
vPWVIdLAc8YznOqu83e04ttslIjNhDwrSaFjTuDdUz4/90pS+9jXHugtDRyMoRXs
TJ7v/T5tKk74340jiFezFf0ySLYPdZ0ERyqRTzl6hOa1hbhC3m/vUFCHMzkW/+HF
e+V5uJPj94FNbLC4WyidFQ0bx08Gr/ZVi09fPXketLtcPzx+VhzwmLdak+HBBp9P
b1jbmEVeB94p6DyBlkYaAh9BCWu5Pef7WPiBczMvlaQeEa4xkwBYRmGg0aOpFVfj
DsUGIweeWJy8Ohz6qxkTVdR+hUEBTpu4J3v5rAJFJmnGbNGxZtAHZEZ8MCAP0/4A
mnzVwtOKv/Ym1R45Xy15lw6Lmht0LBsUTjSz8wzg/zoIlM20juG8o+ltmaiE+2ZG
G5cTc+YSiW8TMRabE4T6+UUEWa9N1CfVsUgnQjJ9ZphtJH6G1sijJHkXo7Z4KfVv
w+16hNAJBlOpjcKUKCqnjBzTkV/D+NgzHc3M0tz4ck9a8bEVWJGREO7tKSan0CR3
X3RHg7/gdixbReWQVbzgmjPcs1BljR0949CyyEgjTyMKI3UXVFADNFRP6ZEVKcZo
1Ahq2Wofa9lSgz/vXdz21Rk+y6+bWfER15ZZw0FH/LskGeoMZL56AA2Zqt2i6EfQ
5mDJkUvC+Yy4peHiLZRuOvmXXqJ7ovfdEzC0Fe4NQgtYjCo29mE4wyr5J32NMnaT
BKX4J6SrWaSTqUEa+ahEIUX0RDBO0moQO6vjUjo0WRYcxTEyClyc1ndEfBTUgcw2
3VMvl/fKsSI5nbshae+Forj8QzUJtfZNEjQOzlzlSz2e1xnaiqrbMYDpJGABlh4D
khVZI7mX/bW3cqoNsx3M6sOIBi1iw0ZPCx3wdQEqYJlF2MwtTph8lbLt59lRUKjs
1yH1GR+HRTRpc94rGff/KS5zWseQqpf5B/IQzyeg//50Fxf8X15Oc2P4pqcnGY7z
JsneSZw6LopSldmtR0U99Onn//of8LGZ62DQdqALPVh9Z2mnJHdktc6xPZxMC6Q9
E5X1Zl6yh0xBHCIz2/uIyxICX4cpSl9jSDxkzrijqzDt/8qKbtPdABRqRmi+lKEz
d5JeOBBrhg4hLpbWg7/1Tgble7OocjC5BOrbmZYsCno4KsHd8YYb7CfWDsdki71i
Y7l3GRcWZsf1CmUubxGbsUx8nUS+5JL+SE3jmD11fHqUzCm3cb4Y8IsmCshJJIkO
Wm3uDa3vYc6pLPiNf7TWmrRaEbwhbhLPdPkdsjXgo2U=
`protect END_PROTECTED
