`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Oh97Iue/JCwZbcE+FNZjsVK17FZM4EkrUDIGnOjIA6e34u9RxaPyzDaa80Qi3oP
+7xLnx/FHG+KK8R2iws7ITg3jNWL9yD3VkIHgmdDri3dnMNOriOfBklva9KaoI/A
Kq1s2qbqXSetf6HZYFYIkwqjDMj0QqE92K5CY7yRcc7VRqwOXe+Dx32WrYp3l40u
d+pFLUoK3kmqHKY/XbQ6jg8r/MCdx+wzOCYus9SaPvqfWzOTkrXvLtsAYHWCoAiW
LsUI7b797lE60beRXKIbRwSrIMWByCBKhgKajFIktDHNPwrlgjcYKt2lwfkkEPMS
aVdDV9tB62tQ7nta7DslmUjCEo/BcLCeMcVvjsvf+UIE+FHnwdKzP4z1ir96zBKf
9Rr3ozH+6blHLNw1VB95bNvi2xSkb6PX6Qtnrss8u7GcQQt+afutI0IKxNPsQyX9
nANP+s/leF6pgXkyMRvIYDO3kE00myEuW//Sp26xRxUYsE1Jk0U0FAga1OsR+veO
nedWzJOPXknNE6RlklDJssWsWSXh2WtiDInKCoh6DE2MEfAdkX2HnDfK+tblkcxR
vs613yuf0ldIGqwqhh2TIQecDNCIlmed08BTXAch/f8oePOf671PerUWAzBA20j1
A/UOe8o3M6CqBYtlbgX8AlQCNK+igsoRzXsbKoqW7KeZD6LlD/hTLAjFl7uzJ/kI
oDv/G7Cd2Z/GKP2dC61PIJUrAYijde9C5Gcun3AKUMG6QG6zjhsskGW1PAgaIboN
tW65Awz827dGWTH7924jdTKqQoux54I9QLc7N8ZBDDLzsMlo53QDVvTTfDCW3Ld6
rs+6AcSWAQiUsqITjWyR4zhTatr+3rEt198wrPIbFTO5mafqH/HAY5MLTWBjihOd
Haq2D83tRuJ+XjuYHBCYOIeeAxqd18SvQvlAM0q0a4n4iqjJZ8Xw8zkqw7xkT6KB
yebsXCO4Ck/kEhL8dKjGaggz2EPtI2zV6IXWhItZol7MME3vNPLT+orD5u94U19g
LIynDNclOolDJ9UulGPsCov+Da+APM5GiW+RWoqRoaZpN+e8ZBj9gSL36fOyXSRx
u19o87W+4SGbIzWmMvO5VRmv78EfLBF8y8KHJEsXjRf3tJ5h+gtTNWXAKOTKOBtC
SucmxTP8w8d00xkjA5HVUhGOmjw4sahB3Q5GXh6y5y1aJ3fJMcuGnXZRbjuo4Od8
ZREg5p9A9V7/K18paPLbBXExQVg0suIm1wvXgXhueIvqB/WofAh2+KMlSptjm5+i
oNBY5m5lCoOixj8AWfVWy4nmWnhZfrMsHgaNjXXp8UX4DYw6SW1K5TN73GOswCfo
9N6wQYZwTt//AhcP2T2AdAuOdRYYsL657OcqNE9s3DKQpc+PFhartnDv4kSTZQSB
VHnpcLhWpC1F4aO5CRWvHSTdoeJjAtk+OiKxuEAE9ry8VUbdg6EXG6AyvdeMf/Jr
LjIw1tQr4vPS7JBEc0zqLw2yeyzkKCqUH3KAfSMHkl/gMKNklRF9sq5ESX6lbYpg
bmDo4ISO8SjWqvA+8hPJ8BubNxHPqshKykutG5mQwKjwlXKIVjj68IA0q0oRGOS7
WRytsIxc4cGiSGPAQLsm36dIApkcPUnFiGs6zyIJE5Kx1Y09F3cBV5nmICgG9KWf
1J646lLDhNZ4nPzRD/ANJSOOJgTA+ZeAwfeyVafxH/Vhs4qUCxM6xO+1Ih5SZuX2
uzSmUhVb64B6Jrj+DU/y2G/URwNf4aQsTkhuMJMyLlH5VtP2H79s8WSOvngUP8oY
awslE+nMHbvx3aKbuRoLnmyjNCXPjtnR887jqYGjhK1oIb4VWZkEboSEdnZC2XkT
tzV/WgLx+fGYlj2BjQNus9pZ0MxjVEdkfk8sMDbygPvMDlVPVxOgXZ3PXbfRQsDj
yOqLQPMwSnHLqoAEJH4MYKpygXI6NVVW04bcncZSb2WN9fzMdrnkJnhlQSB85wOF
csC+kQxDJpy8h0go3rnGQK0q1cc4Z5GJeghH5BPYtf1382fAqJrMgrxqGYH2+QuG
/5yN2wYQ+nOYdbD17ZWFMy6HTnmSQSojkfdB3+q2MzvQ2DBGLkAajzxW8xysGpIk
hTzBdNeDDbZFGqlCY3kPxQDWTYSfelWGU5PJD6Afx2cZG61IRx9lMDElV8EaGOeh
E7uZgZFu6yZQjsG+g6ZYoMG63joXjMY9tIaBDmCZhoazfPF01wChlAJsaQ//smFA
XxUoIP0pnPbCH2B/tLP0V8THD9RKBnShGAK4Lwodtnlpu9Je80/zhBxAnCG38Ndj
/rcWRuWnw38ZmSozGJQekwqe8RVOc0VH7PeGFKdDamXmrE6PsUslNcyUEnY/+Gwj
XdIeO02uqCnCkh9X3Y6CO63YPFC9NQgc0PW/wj+kQ8Pt0AjIB0QQ+RW5CCbZHmU/
BqaXVV9C4riMjMkwNXK6IjQKIwBDSPRT3SdcbpPE0i5IiQv8RHrAIH88Fve7GorD
iJjtH5pg2j0LlBU/hd3Qdf9nn0+bdfcjGI0b/Evfhdf6nzKifQcB1YpDCbP0JruZ
vg+zYWDT4pDnkXjUBaLm1CGAIMQFH7/7gScAmCBXv+fvdOmKWrVI+7kJNyq3Ic12
7Rvlkp+U76ePaW6g5Vv9IjY77L9BH0nXwaIKBmKMo2Ib6Y8dCezZ/C4EzN9AsH7c
iKaZ/E4iajUNoq3QtiqoKwGsGuRSp3IgjgGtDrLgdRWPw5fa8/ilInUhlXfL9JMO
pTBoedWviSq/dlapbTVGxaBZ969ZA+pu3Xl/DZrLheqMh29OUgXro/iakRCKSLjI
+FqEdjcDxGsMZ/6LRHjTXgnV9VCIKa0tudhnc/h9PzAaZFjD9eP6ApF1vnVXnoHM
2q3tiBP7gG5VdtnWF/PqMHsMZ1LfoFtRBdTz4k/8b3XS8XpB4Usk3e0qJHIENoL+
rIz6rY5cGbG+YtIfUaG6ZDwldP+pw+fyWTkIIZsJRCh/IWgVVDb83t3r2+hrMY4S
eqEly9KXn4X6UrCDxDLroXL68jVKKXkm/2G3PEYNHhq+RhS7IHN9vHni5CwQ/9tf
t0vc/oyekjpRkqHE7P3WkNdp3HVqfooGBg4cJ4wlh5c0KPYmg4AAMAtsdt9k1Pmb
qoKKuh/ho4yNVuxiyRqsEnmyq/tXfcexJlh1bJ39XyUcLFZhGH79r2I/kTBSheJr
gldcbl95B29ybHb/NDi+b3ElFF50IwIWESkxo+95fRbGPPq+jnsmcH0p0GQ+grdY
ncwWMy4FzQs8xDQ43fgomFnRguscSSPiNb6k/GklRRpnq+8gpUEJJPIDp+gSFE4A
g8zFoXjNdaSR4FCBLcZx7LiaFtVL4Km3HfDRlH96Rz5ZfbCfbVhb6xr20NrA5AMe
L+o48ijVFCCw7vCLVZKxJ32Q41ret9uuNLKIYjkC4yMW4VyXf+ny1rBV2J3rcPjd
oP8q7BD3wQ9yyDZxT9o8Ys51UKFZYFvi5rUgEnPYiydIR5szQU87FTNMQ7gKGXEL
DKVbt3K4nJM/WJME8NdXTe4Gq1/d7mehk1yAYOOqBTYBz0n49P9hnSVnZUiK+ufd
AL894rm5dJ7plG+mE3znTTC87zRw4AtYMHKVkteJXvb2m0o0giQEDHMeyweOxMlO
Mm1axFz33pl2aE/Ct3/yQx/JOaQL12pzlEaGqdWNLn07FEpoMAp1elkBpHiQS7im
VB9RYjyKjWMWdktekDx80F+HfxteiPOu9He6HYFtNIKAr4kaPHgd0mHpfOMGmCd+
JMHgDxUYKVecCYh+RFOcwm/qvMp3rvEp0xjQW9vmSU3AMdTTUhIsVfFg80/VR3tp
9+9DiUSorSmMAGWgE+Ofu/+lJwa4bqBpOQdj8nFmx7hHwzpX3E09SKlAP6xS4Jwa
MBXCEuHHfEC7r9P1JOLmInsx11x+8FxWXP9AncK5pFg0ASx0jOFGzpjfX5aj9Ymc
JpM9cj1KGi+d9I7uzD0chDLE5OAgn9cpjLNViPUL4L7iOjkT2+0NiH70npoBENOn
KGy13m2nLtntOowF5/JoR3UQCJcN/8nErEOBse12oeuSeCBJivE94IDMfZGGp6Bq
jI5Rf0Q/UB77P56Xi+SuTCgwpEhrZiby/eKehQA35ShobLURO3w1TuG+iQkMqxft
eyy1DrHshbCe35fx9OSzojni4Fim8uqw7vWyOY7ceXfZFx+r40yAfHZEm5hPby3/
y6MRq3GAzeQaxOAmvrS2FZa23yhs5mN+3bMe7JCSCsXQvEv+8DpTVgTOLOUUjiOs
bfHlKKkUMIame4Brpv02sDWIz7nf+4XVfCSz+ur8BwEXSDOesDmUCeGwCen0JP0j
no1nP0LwAR9BB07wCHGB7NlHIAz7jGrGScDupgitC+iVXM2OVBJ8bhy/MQHyVLnr
DNbbiYD0H4dK7CV9iCtWFIS3MR303oD5bLG/0Fci9jO5O+3Acv2RWFWgT/ylVrHo
y33Pswhgo9GJhS3Y+mAoPv1Jeu/Q/Fw1stvMAvtGyFWBJmkBG/Cctl+Kx1nAoOkR
bSdco7D8IfYUOLCWytGne6Q5n0KBVOMXcUFb9cDp8CELnJAKLwRXNjN2ozljThdF
C1zSwDux/cM1OMm94u0zbTekJIubT9wp2Da0uZaIlEW4L+LHdJzMm3x2shn/ps0E
01fA+kSHwz8+Q66zZ5HM2o1MCpjJMq7/RmTwRL+U8Ijfx6YgzIuBYIyf/2xqYYYh
pxXHOSGmxwmWxE66EILhkiUXuO4dlOvnn2jfLKK/MgagUtr/Q4EsKwsiwLKCWnWI
YiP5AkNWyNDbS00KiXX+Fh0hZXthHDTOnpEWWSUBqMBkz2d/mKD5U+Lt2L7JuGTJ
dVrGPaeeKWhjjFkASWBWOu7Vudjf6or8fu0HZRqH+JDpw4m6JQk6oUm7Rjr9Fy3J
GqKm2zO88vO9Iol6SMh7REdtrPE7LP8ZI9l3RjSClltRYQhjIKiseuERZ+jKU4Zo
mlgLohCQjDeAnWpZEsjEXdIql6qtHX9PDrbYvJI1TH7kSc4f6A99ENQmi39eAlWV
y6RwcuyRUvZpLnqpvdnHatjTniHYOUBQFzrSoajF8vvZw2AJCl06c0neSn+TrhCy
QnRq1+xzDgYgvDBQ3ueRhl5+aZONgHf1d6W9Z+aLWaWZ0n68PrznMHWQfjTujeLp
Auta4yVH5Bn47vMXTaI0QzViNFsSaGAcjmSZRNiwfrVG2rUaaRUdbuqESqFd5tj3
pTkkNFkKb+Oe6CFTE1XNY/Z+xiuEAEQJqh3hAY/6/H5HFJW99WZkNP6t1QgMEpzd
Kv9XgrKHMbkanAf8dXvTUKg0eIPLLHP3Pk5AfxiwveEg4EF/njkPT0rXmP9IeC/6
dsNL0khlNBOpK1sx53rNselUtaQ50gdCi2xgUWNIdcpPgdutTBHFW/lh3QDDAFGu
xscasNfUVx36X+kJxeuAH+RIexVGfV0kDyP/rjtji+4xQXNMT6G8apnplmRWp13k
KmVdgJ50kGBbI8taLj0xIAwcFzwSr0uYkRe06zkW4CXAZRHsyM1rAMtfw47/3hmm
qJEmcnlkRQ2X743iEoVlnWC5a8VX3N3nvKxoTMz6RCHuA/ueWbBzJAEnLjXSU74B
raF2g5sxzELbb43+TavO5xXa3a6AQqLNDSKR4XIQ4waooN4WFsavFXX27OL60r10
B5u6Xg286YurpyoQaTW8m2TxvSh19rhmNCiwojAuds5vYpph8JAqxu1UogpoQggW
yNN1f3hNhqhsSv/9Hd23S1XtTCvaMd3T89UhcvBBsyqPuVi/hpcoRq0IUiD6G1mo
6AG8tm4Txbg1EnW4EnNhhpbnIBfYvCNZrVU6baDNJkOGpxcy3ddl9ByhGYJgMcBH
007nBZXa60x6UeZ7UwMM8N/qT+JNyM2JTN6oQa29X5Mbmm4rq4omgrFIORY6kKTD
1fqspp/Wwqw1gtd9RKB5MExzLM/pPS0YRCoKwR0LC7kCoZkOv3otUekA86eNSTOY
bjTY5Kk4xXO6U+MvCnwbfo9H7eHT+PXYxcQsPsslyvdC9Ar+7EkQv+PiAQV/izyu
6C5pJH62Tn8bQGDIntDc6WCordiJaejY6EUMoYNzaHjxeN+AmRM8Z0ojinjJE8Ba
QurA8ZXPR0+n20E38JpsgCClc7qgIfURK/7ScK86WKBLYt0fZ9IX8BldVHhX8REI
TUqJ4Y/MFezgWVXshk4SOozemSj4fauWc+Xp7VSIb4yIzmXda4y1q72Iqr6Wu73o
2Qt/CORepsy3oXLpRYXwlkDIugDbzUDlwT+PE4d9J3XHJPBxidKFnwavakF4z3PJ
HNH/EjHmpFwQeEHonRTTcaUbJog6gVmXOeyj8OaaLUW72K7kznl+3lmBWBnL9LCE
ZKpSqDt0wTG4AHXQK5u8FkPQm4pwICeywHm30XJLDcFaPnIqTxyd0o35ZCMgrIhX
tANHPF5dA8HZsERVDlJpSa5mDcJybailNIycEGgTOJ5moXGNxuH7weCDMlbK//N9
AK/8tdLDBj2nlU7o2LTFAxomjbcnHYrOgusnIjCEMei9V3MaQcWVQy4cAGI6NPIt
qmbB2K6QAYocXI+CtZyXCpNJbpT3T+BCHvXkk0kWxBKhbQG6ekdcRL2iiQ1ehzz3
USVz8Qw0E2JuW0e5t/xoWpr6z0KVCpZrNg0mx4wXgiz94DmmhD2XjLG7VeCa2pGq
m9akqrEX4p/SzrQvRqbBQggE4VHvqcTxLvYDHwwNCJg4gLuLgBtdyFufxpIfnRUZ
PIkODeqmbWSgxFIyOXxOg+Lnl8n5PqcH5ycHPF7IumUsE+EyxZRUvmZ6z7EY0te0
gKhxZZLCfOtjgeOZ1ZFEbk0Zw1+rnxCnuPWqdWV2//ABEcuqFOGUA4u66K0+ly1k
K2/IJNZltrGtgU5lAWQvbKy65OCtqQOLCVsMdza65SdB+zIHRY4bTkkUNZA0y17a
xUrzJtHAjmz+ukRuq5D3D6IM8d3WFGAnDhLtf8+69g30ckZiSvNG9CQMF42T/sxH
PD8jZNRBIvr7HEvNy9OSzKlaxD+gG96hUXv1kv2qVpQSQc06dtLyVLRr4SPGvkFX
1nkjcrnfqest1dA8r/Hnnz1h2ZYm4sxlbRjM7meoJyJo6DhjbFlKxio66pRYigmL
RYzQntV8kOpmiI/pZUUq7ljXnVQ3pB0XFv2Sl9/UFLvV7SFZt3XIF9lFDvQDbp9k
8iYW+yDEAsCV1l8fNyQ4dpEeiLy6ZcqfIXeMrPNgky/W++AeECSPMT5H4j8X/k8A
X8gzxl8qa12hXQne3lHmGiQp9tmHyHcPfl6j0dx9UgnfvAAqEMcTThns1+miXKwE
iudcrlNOaTyu3+2Il9rihtATQMyMhnXUAEjteqXqXmUzRcz54txHjhCa7hLNxCuR
o/Y5e0F6cPDD4rvWhXxUhhPp/mrnnn3oRZ5SwRQEPk2laINhM6IUQ7KxSPd/5CsR
oFwNE39SenQsb0X1nyeQlhsg3w7n7CG46hrluWGYnM8e4LiNOjDlk9RnfWAGavjF
54TMP3NCn4UPcB59bczxr7yV0aqHyd9piulAPuOZmj0UTwKP73jWxJAmyTMshRP8
wJW2PCajDB29SKOumdsbSNNZeWrhbTOdAW9/4pqa1dU6P3NnQJiN8/DmIjDEfS4v
2yAy6F6WGmZD4g3LPII/sMy337MVRTbIEfOz0A8Ew2lcXMtk427RKcYO7OoxRaj2
4PW3GSIXzr4CezmT0qLEHzZf7/cw9FENA5PU8/QfW/JF0Zks036T3fHi/CzuE+mW
Rvlb+lmFTLOEnLMhQjUzMEhe6JtFJ6sqj+sPeSTxihN2TdMovmAZoKCD1FLIFBwM
Wbp914RW+lKTmy1AEYXA37hHYHsCbSLQ4DhBXs8tlgbqE0YnW2Ljb1nrzVJGa/1m
SfuefnpyTfwYcem2ac1oyplVJkGs9cc2Uwuvgdl/o+QKpgUtvFRM7jVWXJ3KM91Y
eW29tVp+jzJFRhvqpw16Tl4Ne9BKP89ap1W5ikR1myfqKxuzONzvmNVGO5IposbY
7FgmO2eYBLFDVpE/hR27c9gh7fh+Yw1nzbJaYhwvgUjAZoZgHsqo/L4zxGPvg0jh
F24gieQAdTnD59GfTu4Bg6GKAND6ke6RaLUspv8lz/sUqos7glb2eCBwKhz05kfN
OcJ9IbgFo3e67K5m7SK2zfuKN4Czl4gnUIBA/CjnCuV/xb5tUkxU5OTLNLCbkHt2
rg+AQh0ccSONgA7Q1BtqxYdKLUeItXuDiZh8eyZD4Pau4WRIFoVOTllxoLpt6r5W
h33hB3YAe8inynSQVUADqllkg7oXLq+okpLZFOoaqlWkftfCcJlw0dB7y743A37X
sI5B5n4Q08hTqz39cETmRSiDc+erR02A8NjT8Z8b5zCnNb6c/uFGblKRE1DaU9XC
5lyACjKTuFfRrucAfyrntNVwEnJDai+VVE/sHrqpMgSwPdoOxNPVwnfxb1OT3xYX
IZUm9PQLbLXj2z+NXp8IaPun31kRQ4mCcg45jaT5RNWK8uNPV/cqGIg5xtDfIrpj
WbSPG/J65roawHvABd85yW7g8eO2apxQTwt2SS3k+mu6060iUDAI2r80BDTVb52r
QOarak4K71vUz6O8CFnsRIWYtTIE9YvMaPPxg8CaWhcxiqSYWObyoMWjZXFgIx0j
09i+BddLB7QNbilei7qVxMeQbzwtr0uJm4ZkD23pEk/HJWiDOnZJEppG5Ycnzvtp
6eQX3G8l2uiy04GFKYJvwSD3iSV7RvPsyYh9mSGHYwGcvoIKDEa4YLC1+RYOdrzC
psciOSTD0hJCmo05AL+Dw6jLuIc9Ok5ejA+eM2oWFgD9mEFMLT8D04Int+KUthh5
Y13pOttePjbiGgWlrZhXDxxnxKBG9Ou6S5JjpoIBrQk6cTMSBxICtjQfHfhd1T/Z
shWT9YonYSvB2F4JOxD9N/C7UfifxU1+NzqqqQfZtlA8llKjmeSQGZwGOfNcDl+S
/nHrH1U//HiYXgVFVm0u5yRqQ1fKiKHHUzGeyLokfgwNJxwr9UYVUNMe6gLl1kOG
AFPgN0anZojI87iCCTXHZKfoxxHOvQvAtPaLyyPX26F1cVsDNjeYKwMU63Wisygb
ppDmRTmBqvFgxHtcwCk/EEiMGSY111HRISUaaopEhgsXdpYJudNlK3S/UmjbVWlE
0j85LZmcu/SGNDqfrn7x0Snq1Z/Bqk7Xy2n0iEJod3tTANwKUkoyPoCU7eeTt2hk
JlrWeKB8KdrM3gy59G8ylZA6asE1K7DAXq5HrfEpDMtrHFaIZx95ohpmWBHgam5w
FzQ/qYhIcAcefOPL8WrKub2cusTUpWFGlwQOX4H338ZB4TKUX3BShD2pkXNPMO8L
KNqN6BrJEXUJO480DgvkInBZKGGGknF2+Ds2RFndhrRkbngqG93HOQOTzn8BCI1F
WWILyaL7ovJ8tkQntmdfOGRH14kI3aPA6gn50Ydg/2ngG9JaubHYAcfRN05j1jjk
C/fNbC5F9NMpXFBc7X3D+qeObuBNetSrw190M21tDEOgORsNE99zbB3xvrLOtwai
w/0cYy0TLvWw8hfHWny5NVRuuhjsY8xCEm6sfH/WaOQ8sO8Zn0LAXXT2/+VRenJ/
1Z5zvfT/ewkOVd+nfQpvcl98eiQhcZAOg/W525KzOw9o+r0weNjTWY5e+FRJamK+
cFnwvyQaLK2TwDAn54Xmoau8K9kyHhnbzhPmoCJ2v8zaYYbP78JqjBjVz9dN8NO3
1AHObCQU+QnCv2Y52AqdD7a37N5HIoeVq1sm9GYr+1xgE1bdfrDFC9lOucfM2UsY
IEsyCByus+a1vTU4UogJ3KmMnOu4b4wcATTII8j26Oe70uHQ3ITbCcd2wiJ8E/mJ
VuuWcZbjy8ar78TWXQhJeyKoKM8T6UkHoQ/hJ0dB/hnpkNfj05AH7pn8cNGge0SM
K3eYtF6xuSZ0JL900LvHA8nNZ+cch0Np6ZOHVd8ly1hik1CUtgxqSIooRIklGQmd
69Ha+hLltbkmNY++ndlx/vq827khsLowp60c91ioBLwbpZK7R6m0nCZKhXprZLMp
GUUd66/hpiDCSUODgfpBiRGPOvuvSubjG5LlEjEDPpUU+47Ty0+iOuMAYL25qIZ1
Iw5GSL0QkjnFCWXqInziW+jYE7QENLxmtbIUn/+uFS9rjLXHLfcBE5JMXQDU/dns
UxpbFnSYQbq+BoG/RpNJdSOUnyxcFs54RGxCv1QdHXc4c3TqcrFcfN3N2jc30wZN
bx44XgvObu0QheEcma274pclezJscm3t0QyeoZ0GySV7hpmw65zGSxlv+C7Dz7XJ
1KTo3WtrssnhObwUun9LO/aoeQkpbD4Yt4USLwFjbtvb0+teqFlA3+yddU8WjBFZ
m8luAjgNiwiW/hiHH80A6AM3htfEQVhZ6s2NubLo92LaSoCtnuXzdKVhkP9C8WIh
mBkl8zOOBghmaRqBi/fgryX1U+ME1PkcPxoYowqS5YesRqqj0bFMIrCdc+fKG1Zl
YEYdK6Wfq65ijLGhY0muRkh8jV1hJ2EzcqvOZ3nyPsOmCPaUTcJ/FgFP8NDkLwxK
lG8S1c4oNMUzzAR2wgHVJCSKcZXoWCHtbCSH+9UMLC2eLVa+GjEyYmooXQ5ZSu6T
Ygt7/lNTIMp7SS8bfFvJBIX06Eqv25LhtpAD+fZoPd92KRfAeMfFQRt8SW05DgVj
3TNkLR6DeOrGCp5FRxotbyxW88iRVPXm8YKICRIo4nD6ciei+5tG1zvPx0b2X6mL
M3hmFk38ohUQw/zETXrTVXzZqNE9xUCx3pRo6NIozLwqXN1WI9yD/gS/hzoT+SpD
rGBPPhy2efzs7L1YreDUILROH/0ZDGIw2GUST/vaMJTx9XfM2FS4yIjUUFI+MQEm
cIiTzttCQOUbMl05KkAlFTy/Kcav7Pl+ahzG5ZNv/96PoV3mxIRl5bjIxXK9Aqra
ZuvSnW2z90vHokpXTbY9OWGSv+Kwegd3jLw1uUgfpZauG9OAg8VTumIUBpApjLNr
aZ2R3DL69xOFpu61wQUpX3KY0txLWjJsKcCy0A+mcKNHPkYYhf1RUzmwp84IHG1s
qoJSB3ZJaQKivKgiF6cafsfuQ+ulLjg0X9cepgjaRovTv7lKUQSgO3xjcoMbQnwg
IRwN777qfTh/FOboWPkLHs3ilznM6a0JgZwcGo1//4nebypPcyvjJyrjC2TeW4gd
qzUk6+1xTan3jFPfRrNT/gfF+7tDTFD+zFdnRhB408QW3yRxXLp94uSwoacOdy7H
RFMXIUtyhXOEqu2/R7WvXP4doeOCy8pDYKePe0F9+LqJnhyA0x/xjbmVn+wn5dr7
ITIUHIp70AwhoksZERLZZIw16kuvOp/FG+4wkg+1iYKpmt91IuXrE/Zx9sfDL7Qj
crewFVubYMuTlxxSOoDzGnLSvb6M9mAtzXINbqDGm9cVB4w8Rw9JCCulJzo6jS8c
WhaO6HbPimm+9aKK6RO5/p4jnrfJgX0Kcrg7vvDx5WoZNfYzrryMqqyl+GALxB25
unIddfTDi3LrY7WZjh3/X4jfWeEnJ+DRmyAM6rfyWV5symloHkkSVQ34AzI7LvT3
UmL77a4D7AzGwxzyiMOtL6ta6uOvUVNT9B7rfVXwi7UkOxjWAaPpNot98x2sbiXr
ygchzvYzjyewDwuSiHBFPU67szR2E2kaRBi0XnmkpDR5TUqRqRCCBXo8E0hEEDQy
CRn4yD86OyG584ODfgrFgjW2IyKrrNGQRvz8ssXQuMKXiZ3f3UJUi1suqnR45Se+
EfWanYI/4Un14WQPgGezhS/da1Tj7iUUO+LM7HdbSnISSmgUqQNewfArVetCs6pn
l+vTa+k9Twx5YFZ/Xpd9XeP3a1boCrQRasvXXVbjPD/vViS6Y0oORrfOIP88AiwW
iaBNz51Gl4mYyoJkF6OuORmBKyxxvMWym81BKoIzlhzoieHSSIoNVVM9l2SHmPYf
Dy1JCBKn0cRwh4VbI8bZwcAogObGvb/tN4touOJzlR5fnytM1Acw51JklkSwfHmJ
EIDL6SsfyDKHX+eIEFuOh+FKzNlqJr+/yBnpdTHC6vbeZPmsh5Nc9FqcCNbBjUzZ
2FZYjVt5n3rdUu/fO5LWAlkiPMztQY+FGKiJ/P9PPvXadprzBc7oa+6yp7seGn4L
coLPSHkDtymzW9roonbgNO5XWTJ5tP+1YDo3YF8rk2ULeCqXu4c946AIAF6Hn7eD
2bKRVQysns+wE74cdhzKr73eYgbSS20bFBdVoHZO5e02dR2lY3egj/6cE96nC5C6
TRtCbg7qykQARFb+2XEqjfrOxjJ+NuhvE9q7qzGpNIVHvPHpvwtdPhrFDRLOajP0
g+CZSweWODSAx4PTAJOpr9gTmYnLHQ4xzbvlRoQ6u/MKJlv58RsFI1eObDzRJjNH
UJSdvlTUKpc+HShE5v1Bk1tldTyXbO8Z9ZKgBGXC6HLblXQm4jCseP6Qyjt9lrHF
lTWktK4YXBy5o3m8gsVLkocqoIDJI6OY/Va5iPlgI7AnIwh0Uaw2svfM5NPZbVoc
WFRKqajI6QrZT0AhaIREcXH1w11pN6KhlipSf/7sDYqMIHE2JGXzABlWdO5pERPd
TDnr1oa4X3OHTMSDCf/YgOzT8S3YcpWu/sMp/fjKwBvVB3CPB/hKkBhHfS1HlAcg
43YuYC75+R3p9F4g2u0ubfciCzPjp2+EckYiNDITqZ07PsTl6+OAFROyXybdOYHC
eGfy6TdbGYDGgge5X1d3rDZxuwUYcHF2bWsr/uINe4Dth7gqnMuZwIiknZhSGvKG
X+xszDn8s9fMfUxeWU8Q7KZLUtkwWklzPxJz4RqygpOE+QKFEIygBekl8WbmiWhI
jPAGIvheIzLJe4979HxqluQzO8lPJ1Ubl8O1lHYuIiiZhXvm7Wqg5zt+qD+c6NlF
7hlO38HX10lgxgR68r/60Joxs0tNZx8WRRktJjA30uHk7P43GfVA1gJt8oPSHhvM
Gyax0X07uVsTjSy/8rgwEzg+ji7dpBdIEIM7xka2psLH7UUg2VaGGUEJSSid4pjE
2wXIpom3Mk2tsaT8VasGP98JIwI59nrx2TybIqBNItzcq2c9RTWCQj9IJ4SoqOG2
Crh3E4JkgzKvQLyY4R2Y40GhIFLAB71OKLqDYXwkkVbo+g9xYTbCUtepckMd0FNr
Z46VK6gbnCNSfNVOdgHYMy3WAMCk1kxftxqlsEQD18n3dE0eoxrzE5PD8A4fdmyr
LEdz0LqqSZ7cPEkdtuNfHwwELbu0iV1rFQq+5TrNi0r69dcQx2kzMUzedLP1Qslg
7LX5dWbEVOT9MQ/1/g3pbmvYMi0SRMJMz6OrnzRn+VoyDp69vwHSSXUh3w5Ljtv/
y+Zps1z1qhYXAK+dBsaPrg2mAIK+Zqs8tRCHVVpURK3+XQ1yQY7+wtKKFeIcfwAr
RaJ0K+yloa6+k9oIup3m6Fl6DF3ktThRzlOUt57oC3DntpvckCx6gKQQEgs632Yi
R58lLQRmRg9IS2BFzTqvGqHZzN5UsY8MbwE+qUQtCMMMcsnPDM9MwWWw32nBUqsp
/Lcs77uIQB98AQdWytap2/ijxi4vcxZP05DYHlbj4XTQVQ8+VxaXjdl0ovfPzL+X
iPgYvQsAJqFYyJMdl30FSZhJ+fC2/8k0psJwN8b7lT2Zo7FWicYyBIbvreD31JPo
cl7OsGkTFvVj2Olad1al11LWfEoejNRXPnJkR3dDhdP2bnACBIfELDfkAHjf8deL
9qHa+xgUCimjbzKpbGFj9TxrAf6esIRe4PVgdx9dKSEEMwaqlUN7S/CznD95ol37
FWyV1STMLfpDPtRnhDpV/Wmjo+kV/jjCctQPIiSyb7kI21R7eijtD/MORvDXDAPV
Th4d/uk1uTahtveSm187c+CdPPtcbrVOVydEp0xaHg5NZCyQunv3ANDHW72wUnBi
XllLe+iFcm0YK+Otha/rzZpPc9Spr9uQ0SHuJEn9K6ZU5pMTvkSEbJ3cVEJodciX
vkFQ2uM5O8HWLPZ4eDBX7+JDlPpC+voqK2k9EWwAsZCP/TzepLP0tjdfV4FGIz9n
3NdFz3X8lcLKVzXBphYhtlE3uu7GOKonpi7+aIE8WmNP70Mi+EDgj1lXRxUgRxwk
eorcM/G0VPDQIjy8Hsuohm6mtAAy4LSTHSnp9a0I0dVJA1S9+ikSdqOPnWCWoX2Y
wDbpmxy7W2jrO6bURDPiO5uRmSE+zBQ93jpwS1LXDvCsTo4C5n1syDgamSH0kEz0
hb0n8xD6hXFNtMOlgrS7LQm7Emd2RZ6Pu9PTR89rYxF4czeOG67vzDgcWuhXAh0+
A4QUIq85ByFBOZHmND4Dka9VlhgTIjo7ZkuJ8SDtofm0X3yCshGRpceFWO4wzr/2
bXLkgt4Aq5gBWfqX2csT4cEm++EVLc83FHwokUtXMQGSIslqjwP2n+OzdA/wayQ6
VbNcThEiseL7CPpv8uOVpiYYPFz2WRh+ApSqlX+UII4TfIN+npgv0Kdeogv7P9lh
ETYrOGHHC/wnuRCjtJzHTy69Ly+0X5qtvpbREuSHUHIcw6jJQ6bE7VX0SSEVfyxf
woC+fZ55E5sTnxqNInEwAkoDkD3V1i1TAs3vEq9a98ba7gp+YSF5vXVSVNSMBizR
FXuSuWOLrUB1Rj5uC7B25MxO/9NDNXL2d1blEeItX6bS21lOl+Co0NcE5AJNYvyK
sWjXpoyqOWT29NAa23nzAT8urA/dA69mvtTgswNn2NnmUTzWjm+oL4U/n/Msnk4V
07pSA/oyAJ6K0VYWu2TNlZ4ALEQyDty8MoI9P/slVD10tPm6Tz0AVFd+vNd5nljm
RSDzj15TVWVuG/QJ/Q1FMuigYk9NagO21aUDsSJXxVoBsQ1HlSKgK6/wRJYlwhBN
/Mt4nWzqhlY9JexatsULg50j2AAOy9t/iNsgZlFM11S+Mh3rIPfzV4MJ6pRDbG1C
8d/kH081Dqom+19LgTew4Xz2zNguH1MfsAYUuu4Xx6MDKHi0GzVahPxNkqX7urN9
Qumgj4NA6rH6h0y1rH+zq49VASAd30XA8Lqx0+fRELkJumTcyTL2y0wO4h7zVLBd
nX4rr6vahCenSWx4nJ/TqHRaet+SGFw+jKu6Nx7wXTqkpdF3h+vM3QdKw1VzENWl
JExnaurm2+iwUCHG6PwL2vPJ+hCF2Q4v2Ft/apRPp1LYL/410vfKnN1QYo6rZwjf
JoyXS8YKZHa8S9EWDsvUPxDlEB/O2j0NeQWp6VRvdfYDsqNS30VHG5MbEo/YzIam
CA2l2XqyQ3hBaqlK47TDmGrU1ejAl8P6Jp+/5Vmk68H+k0IKzkbXHm2aVRWcWpND
nkPVARr4Xoe6KmBZxOMmcbRpv/C4ejnrbhjlBhLuU3O6sQ2wthF7nINX+ZmItzg8
DhaLtbXcqfod8InTbDVq9rkrFYh2le8OHGqm3nm8u+XGgxJ/o/9GDruJ1ZiVti8g
qljKjeEAcpjTwGsLG2lLgoBQ8DyKeoNvZK+nQjlZmHx66vp9rIq8pX7pfGsanEvk
Jub0p867PFFJVEMNKEA6Nb9vjuIjqyiHK/UCY39Ngn5n7CKaqrwdVu+In08WvWoj
ROb1ibBvaw8QDj6iYsIrkqHaMIbtNmrqV08yPDDnGLI92KTu+7kXljc5gDqDf5UU
L6sfwoU+NRJNLjaIGBTLRSQJFog4qoX/c/NFEOywGtFOlwP7ER6AXNMHmgzmrZxC
WgMuMJcmfwe/Gkx0PDO7DeEre+ei3kKj31/nCxP2QqufQCqT/OMzQAf8lmXSe998
DkJwSE/z1URBlW5v0lSDRAHmJ01TP/IAdirPz9yFKbwGgn12VMFQS22nnYOUW3MI
nHeLfiZp9IKQrmjacm1dSB1GQVOR2fyFGTKQqn5al35EjHy4EKpbizuuLFKR/wBx
ISpmpKg1FQL5mzDGbPp8O1bT+kWjg5YSebCQC45MxovsQ69cGbPifhXJ9uNIRcjx
SPtEtkJ8lCPvrgJ0OqrbXuFKEcmelr8O4oZqYA0NNaUReAfieHtH64BL1oYSMhOk
3s4NkdK5nn7+3Q7f+yqJMLv3Pr9H1dh1uI6YKeUIcMEL1WAB8faQFLoCnjZexfyW
d6iHtngGAzw5SjnlFKHpBFX8XETKZbtzSbpNpMacymLYJtov1VEU4S+okxLSgSz+
JXqCicaXbIfJwXaWk1btgnPwgJZtNGdit5SehJclXyeNr7WS+67qhNv3h+DN8YA5
iBCtQCtxJfvZozTcqu4rB5y9IyMV9tPYvRlt00+dcn7e78DQEBFEZUnj5qcdW/Jb
kP7E7+1P82FfUA/yIM6PEFHzb5Ty6yShMes7NEz/SVHb5JGge0+Joxn3V+CUaVSv
xUuEj9D3B1NOEbty407o4xa/maBvEBYkW6nf9TiVjWQb4V4pXqHT4Y5wuljqmB1v
bxdxP+u7KJcteYGKz+iyBJpa1Ypxi/SUc5XnoAkmqQP5CY5JPFyv3GAVOu+eOhzP
1bytNC58DfBwKL/pGvopOvJNZTmpqUNO0hotNgcFEq7Y6j//2ZhPRhs2kBSOyT8A
3lyNVojA/zaU61iiqAAzDmxoMaNkXXqeaDdJfYDymkfBl5OCxYnVNw5NZEg9qe+P
vxHUfSsyxSaFTeruIDNVWbe/lCYyIArjAUwRCTa9iopiJwvI3J900p1Wetiwl6OO
KP0pPSRASJOJyQajOLXLmJNSaTq+cMoz/YSw6/h4sgYvCTnjYHNZG34pHSbsDelb
UeqIINP4o++GZCDEH1kvhB6z8SNK6Ty3kVvvm4QvEcgr+oPO4cxlzowfXhQET4LC
niIhjd+9t16N3BxCgF8XzNKIl3+h8Ds2UzD9unHVJPzJff7xBwH+coE+37zPZ/wk
eF0ccC8FpD3tzzYe3yW9RbqCrKyuBu4RmL81ITkceVQvvZwGHMTO9vUs4oAOUvND
bAcg8dVcaszFi4XtvvaQoLml9DjYz+vCTLmO2wIoi3Zj+fhz3oa8cUV0GWlg4aOy
uZvaGmZLBJP4LIM3/OQrqNeH+aZ5UU0/jxjUVCSr8KCDr2IG+3kcx84WrRrQN3xh
yikzfDYgMB+MV28+OmOkWVjT41VObU8hiTaonvKjZhAKQtlqT6r6i2bmX9O0VT7E
SE/FF+S+WNOZrYPl7FV6KMBEax/i8InPE9venpJC+0yKtvkU69VizCV1cmWsAXdQ
dBxaYyyZHOfkTcilAeRElvoGdMpirr8MKCEm6gvUdteipWdf0mz1+58IhDsyQhnl
B5hbLOldpBXBDWopyj3sm0/WXIaTv7dK3NdU68wjje6vuFJI/mbH+qwNLCmhRq9r
kggxvWcCTpNGlionE1IOAj+JziJuFIDzeDdZbJGBXNjI82zaDrsV2fd4S+jfISeD
6feQpVHZ9+Q/z9JGoBAdljknfieo96/vwOLrJLxIZ7Dol3epnK2TUyY6xq5MBmmx
KnLNnR2iqvjMu6RGaSqe7SLA7QoObbFIEyZTeEFt5fWel7alOksNUJL0vonGw9NC
zn23g4lkKDMt8FWhD1gXHjCkjw5TTz0Oe0vvsfO4/57jotO8LZdRJsYwXTr7sjYW
X6I/n9UdV4Df/Evg32ImIiO1M5bSXGa7Qk/Dy9n89gW3/ZGIdXC+Xjw3kf3eAOhQ
i72eOBslsYNmUFE8czdUd/5hm819epHB9ngXYnSfYc8SpFWB99zkAdM8a5DLpMoI
yZVFzonqfjXj7JZkVn1Sld1J7aG5SCLH4DbGdeHaQ9BN0IcX4YbpblSThS9NBp8m
O31+EYc/ETaaE9FgkfZcx4aLB3HhVKVcXh08A6svrcQEUOkFUnvEiq3bKC3P5L3d
wuxoC9zZIgAjPESHI9MEfJ0uaLLDM4+0G8cGgVYE/DcHePoUv8rgZcs1OsSwa80A
7umHwpGLjC9d91qpSPWjrtC99W1ZguVZuOyP+67mrQHtlMMAOTaZ5wSOJepcD2k8
+oeq9W5dPxc440jTofFHorYlzCYm0i3dIn/LTCU9m10jqS70I1mcwkeXP3f42zH1
iLB0mCnoov6q8l3ofbz7l/iZJYrVyFk0S+1fzCH44LgbclwZcTzXZuuKQHTy+myG
r4wxnhEfwWmGLaAbMM0YZmzEeiVz2MlPI1+DYh4xjTwDdPYOeJmd0cMyYTJ/SnnS
pe8Ummk5jhp2vOwGFNvxswXTIHVNS+KMmrzJwNFog+uTPTyEc1BUBUIsAAa+sTBB
JmpD69ULL/lU+3r0ZfyJBUQdSVf+ZEP7YgZ/WLFHeYdSfmz+mQJVkdkClOTyTxX1
Sr3Gf2YKUgb+vkZG1ZBtXQwr9zKeumNdGBGXCp57Oy9tAmIxW7t+UGpSPkhJVlk+
00OBlUBrnNCJzEg3vUWLtjMNWluG8D4Uzf4TdgwZlylf554hZhWVAcnwmy/W2BLX
/jQLRgVmj9NGqC7f+TQn8EyYsntK5Vqzk8F9gOl8OvrPs5UyubBrt+2c+wU3uXMA
/jMsTU7jfRNlywLyquLZJgrgpqI1lAlcSUARKlCEWnN9kET7+pNcDxEwWuikRwSw
I29npaSGkk9a+rlflbXYgAqI74hlS6TqVcBip9Ypq0U3phbe8JAhLOIDz0jxxaoC
3Oi4bGKZfKduerpJAOSZSq5Z5HKX+JnjV7koykgqETCdHXleEN07BgIH9VRmLgYM
Zz/uDkD5x473R6h1VI38yWf94fPTXMzy16HIsZ78tIFv/Gtrz71S8pZRc+HiL56g
gmDRi3lyR3n/0eECGRIPnCJiD0dQCTVyrr08CYYuIXNC0lxTr7z3ZR3Pz67U4X/8
+1r5z3DcyplIEWq3QAsYOVMfQOlm+Od1xCzh65O4vHavFIL5XNwuTjNdSRp2qCK1
4wmJP+GdH6yQWsU80mLGmKiUdOGi9/rXW3RGSDlz+u0yzABePk3S1txKvJqtgUNI
EJk0ILcCKlCnTB9Yz7kyRArK6rj8VOVrQXmY85vqZFeKrPTnHSeavfQO8VviDRNc
st1wEuevmNgBwn20Lg/HTeCZQB3Ie5zSdQrPmpDCD9u742RfhB/ek8S6f5AzeZO9
o6OUK0wbml4ED3ocXSU7hJom9up5Zn0hnZdNfD6zi6OJ3wEZWawosWGeayKqP4C2
aeTAlbC4v8aMhgUyiD/8KJSas2EZo3938w9+gcc3jGHY9bMzuyj5UzKC11HV8Gzz
2LYQY9f3r9X1GsRgxVX2RsrJnvdVlDSGYPcdbgYpJiOQAupLiadJRWtyrAR88d0B
nrYYRZxbliLNyF2UcTlf/cdYAw7e5xRt02Vn6Z1m4Zm1NGj0AEeIZWbSWvuOb+U6
mXrv8sK84Z+M2xVPqOMOA0ENYl8B8Ne5vhq4D6fCzI/TYqT6B7wiszT4ShGQyz7m
RVJrmriW1jSFd5GRIb5/mtf0Fmk5kUHjJbw2Qv5E2cwuzmVZwuBtf1lqaTyJI2D+
SqPgHDvaYjMeCUoMs0EY+PVTcbueQ6x0Q0Qwkd3ELeZbsIQeZnj0bUyfoBGGcW5T
OrNkh5cZRIUcjBdyjVYaR34GDbCIEsGheErSUYJ4oQ4Iq/s/It5RmQDXWfbOGACJ
ZW0QXYmiXhosU16eaSfbJy1pZPzFU7rBX9iXvR5BpK9L8S/jB+MpBOFrsN4wvx/k
QlrV6vBbz71esWYglpgfwSKXQaWGPAfBo8OO6+J7dN5GGjAB0ncN9u1zaZWLbLxn
pR3DRBtn5XZ07vhLAcU7RCGLgxkMRBuakoX1t9WLZavQcaOzWUtWvqqva+eYlb6s
sbUared/oCvPnp01VERZZ49PoH9+c/XAyed83X/a246RWx8NGqday+fLuvzcSWgv
p8jWhQQCwQorbztqX94mMlZZGNiOjOioGkJudfExnt6WzRxcS90N2f/u/weEehKA
aAZRsNc0HEaO1G3WTfgaxNRW3x9ZgFHJNS1XHQkHZjspNk4zQgCgFheJEXJ8Eyhf
OHs9xOXwxTD2CE+lmhU2w8emcQogEP6KZSJh9cIzLnaXjQ6CDMkAQzzS02kSlgXN
MEqSQfFg2GO0k/a832ieQV+xne8DE5g7DxPQ+9KA7mljsaF4x31YWcJxm8wyLWhO
P2do16ZR1d0olpzpPrvn7X/MpF3EeA32GbpeDGuTdU/LpyCfha5D50Lqzu7+8RyW
QwdojK0kcNo+GOVwhVK798dBVoKvc1Xv9BbnpW2witNHPxyAoM5sxlGx8tdZPiOB
2adeoQcUL+WTIPnjcfzosTvRuedKOb4Gp0wMKgYG7QBftb2lMX6qqTx+JD84g6DQ
Cwi44q+YQPiyWhg90zrcWlFI19kL+SurFbsiHYZQQE/3IDoE9YksyV/vP/PwE/4O
BjDTtFKCGPqpBONnIHxS5DdpESRTbGgY3RCiY8JApcOxxZ5TO0MlgfklztOKuOKw
FE6lESf+n/kDDQU4JB3gH8jRqpaMM/w28wC7v3D+ToxtC4bol724pkoyQgSwgJku
ujuz5vBlr/dAzwl9S7fpUbAr91TdMVUto3uC21jqJIOaCWp/swQUxMjW8znFhvDX
P0QxH5E4sfpRr6cwfiAzssNGBIDvhF3tmNlXw958NOj9gc2e6+vCveilOO6Xr1v2
LxBdBHgS3QA36NXG2WNeRcl7v0nQCL5gXXqTOstrlOzSYRDD7x5va/kSEut5RD4H
WY2flGyAELQ/zIgmnLxgdS+JByUC1I9yMhTMDp++vbPbdF021SM/4FbZrUYMz1oN
RNIHq+Sgo4ce1HFK6Yc4zYBG0z+ckAArcnz3NMOkSz36afFltPmk46LSD/u5Svjw
nUJEHF/eufSHVh8HZRD+3nwLgjT1ONvvbck5INhRGL3+dME6h0LLMk6ut6Q98/Fj
M6OFXxoQ90AjfZ9b1FwMskYE8Y0x3vQRFQ3eD3I1nkKVMnF/rP+ueuJb7gC9hhEx
YQ5qSpzb2ATFT0fWBWTo49DclCsBGxPlV2+liBS/1B/i55MPuXhLSZqM2b7Ux6vw
PQ8tkuk4wmA3G3sOPphwlFADwROezdgAG72OeYJIh8sHwykSpNlLpjDJozNhT0hG
Aww3XiCCGzG5wzY0uwIzbGJND6zfofowiJeqtpiEI4Zfi+FtdcWvUGVWazplGrT1
MRfIQkyWXEK2ms6ZJ0rvbHsCj6gG8WSTgzylp2/DN7KEeKTQ75v/ZDIJbNL7/RDC
6FbEIlDNLqgCYkRWAkN3MhBN5T4Q5VyX7r/Xao5xW6n42GLkR5bi9/PMcM6prtgE
qAKJgPemtXhjLMwX5dVvIu9sLb1K6qvYODSB6uyANZ9T+9VTSDu3uc9TIgL1418T
/iq9B2020rphiggdfgWNP1AYiYGhsioOc6IxfEK+DHP9YLlmizdvVpFK2wGwJ2cW
iR3Sqpl5debTsJGqcklIyYKZi9x0gPxiwy56KjLHQNlDKEoqwMIwWzhVPxvTTPY+
fFsa81k2Qu2JTmqn5sVY8A58j+SOkTD9aOiZdUVFZ8fHI+nEuGsVHv4Ye/LjXG17
D2iePthItS9DOIPWO2pBjdNeyyDQKOGbKKhHtR/+2pobO1FcbXbI2t6Nx8cvNYDK
RA39DMOdoeB4pZOZeWjmsnXy9YKxg5pKDsnZ9jL6Euj7NeM0ZKLIRkKRPLRBcUiA
Ui4x6umZq02ZOBJl+qeIPi9Q6s68bijglFtFDHJPuKxFD3U9LJcaOBi9jBHqczoQ
jFe0FM9TZFqkWzZZtPl/85TgFmsk2gPd1hlAkFRtZ/usBWTWiqER9xqucE6tQZw6
NemGoW4y4u+Th4JY9vRggj9uGdtFimrB9Fxo/YQxESO3vUCpxqZx171LIvyxJiqJ
5ldrViqIPlfinHAaJLnp2HorC23cnQPOxC3Qjwjhin9YIpllfO4zdqK45WyNEbHv
nsoUb8XTagNfjI6iZT/dbPniJNSqCI0BmtsrghZjFd3E+7gS5c/K609lQk7oI4wM
ixKyaAcyNMs16C23aDG1UNKEI9D+MRPSiZDoxgnJbDF4l/1LrIy+pzSSbnZjnYEI
vCAzEL2yATbvGZDoOaOLGHVn0Wa+lkJNaIB49VEQe913c7iicaO0PTq6qK3czEZh
3+x1WsVm/JU6iSNAgmOmvUKSU2/Y2YIj6ADycGX7lEJ2z6IODmkvLzlE2JGXCXaV
t3BoPY+5j4VMz4jvYqI5NI4ZmtmErwqxDcnOwxI5uuSxegJtDgifuKnPZhVJfG5r
+XpzYZ6kM8XrdrSqktXaFuFwRVyu//iqEDnFGF/CRtAnb+cowAqr9hgDL/zMLOv+
QQp9oJtise1QgbLlbr61P9J8crGqWC8aByHGZPjizEI/Jwe1lg87bErRlDnfiTBA
cV7kdCUGmOUZwb5DWkaTUrFEKWKHqEL/6eP9xYtTynahEkBCbizVkIYYX2s4C7/2
S23io8VTw2UnCiPeREpqfzKNY9N4j85lPIJGkJcBiIBwJX51cOXXwWswjDE7af/V
C7OeMgWMr8r8YUvckQpttIxp1MaLl4Ku//A+QQwVmwKsYC1uTcZcoRgWTev1ueRV
E59u6u4FFq1p5vErLyV6cM31W5nrEZi60Azt/SF8c7v2ONVbkyaL9YgnCpgAj+IX
p3H05lYfUNKW/98m8Nht8kAjLBCRlrPar2e1q/lUKbHcHdaPyb0CpwevfNqUwvMb
6ipBgZG8GllofRQ94SJbpW9YuUCOK2nY77FbprzWlxSYkuqH1bnCeKphk9aQzWNx
8udYwptk9a1HaKGYY5dZv5AtRekFKXQ5tuVGdHMHzjmJBguN9wlKdC2BQw/i0nW0
5ms+44ElWfGO4JDzAbko4xTbeQwyqRs1pGwW0bO847kyxQiXLrCQlTPpUzk2rk1T
2ov7TTJaqiLHl0mrXGwB/ooSwnqwhjwBr29bhWf2UJ7I4j5P0I597idQGEoaE4dI
H+p+N5nUHeuX/nbV4Ls1iIY15+l/BZRgh14ZozjoCxUdc2FKKdYuheE4D9Owj9AK
UP5meZ7gwOqnswhJ7hIdRx1liPLn2XA4GHjgWOihMTMhS93eMHK6gucLrHVHOgkr
bfiP9JkvLQdCy0/hva+FWSpr9LprunaYnYnNLC6DBB4MNaHzAILl2OWgkx9p4RW4
g9vh6rQPgbFf4qApmFsLl3glMBB6GUidP2M0zvdP5LYwdmlT3jFHAnTar8yuNFtG
EWvHgI3+3CnvhXQqPacZAL37Ix85ZRjQqFnoQzdGunJIjLfNFmluQVVDxzrYR53t
kRT24uKN9vr+5bIwAhBT40pUPPAqK+fTUoYNdJSJe5tKf5hpw2Yjt8IpYlDTBozq
SZ1K+8Wi7VW1O/5tGhA01sLv6ILtv6OO4/HY6uZewzBpfOUPTvpjAt9w8gdlt9O5
CnBSmcyN57/Or6yaZtjDI3r8TLSwfvZoxDxDo9FjzvzYOoLXrHM08fLpkc1bhd4l
fmqRf95tTYybJpM+aJHsVVyxSKOCqPCCe75GIKf0dzcQyQbKlmQU7o+eb2HIiMf8
mvI7OA3ehSyYgH+GOYvlYVGGYoTVBMIudAj5TdRY2rA6YkwgJUYZpULdPMwHMBz9
TatHJ69poZFH8YQh0Y4Dq2DP/gDi3arxTUBXJuDfLI0r/pbfdzhguAuiJ4B6Q/7X
/R53dKht6OH8RET7VAGj7H0A+ZLaGJWpNn5xfreQEpcsWu/QVHaPyy7Caw7b00NU
cuZwAVO27GJPSPwirKmnxLfFSkN5Ffjmoi2N8UnGQ5JqTzssBIhb2loZKz/r9DEQ
v9OB0D6H459zvt/EMxIEBaJ7JLpSN4oeGNSMfcTTMmVsIum5bocJ6TAfU081FU1p
f5o6upT3AaY8zJWNpEgSKqxruqsn+PIo88+YfiW1NlY/cLIIKgIkp40bIapBVy5c
2rZzlgOHZyrXD8SbKVu5sWnkpgt2LnpGMUC7QAVBfj2QYEObNGgQT75Ax9Ne/GtB
ZVp+TJnkvPPkRqFLXYOqA4DHhSvrlVqfU+fkqD9Ar1ht1JHtPYqSsjbvdvRON8Xg
z/PzmFPiyxed+bhKjlvsn5R6XZGbyhgThYYmUX7A/zlGdmSd/QpFJ/68rlt8oW1k
CXuwOuyyQxGXQ6RuLPIdP0QAp/CNNYrPJaIy4D+AOnF0l5iFHCxEG8ZpOzDQLRn9
6V7xFOgSdKrZDR0u/4G+lGgTQQhpBgR4AFxqVilavlZytOslq0C04Wr9FEgj10FX
qiSvOQFEU4TXr1am53/2ZJbqoa/X3Tx26SibwIp1DT1ZNr8yiYra/dZfFF4Htd/X
20ZuWx9r5rWa0O0NTfssR/xe+rOQBlQZLozGevBfw+HmKvpq2+I3g1rC47vUkSrl
+We8UtCnredjeiyBionqWrnZbjWUUkYR2DpSEMXAw4ydTyAUbSxVZGHAp4xprYVw
+3zF4Yck0kZZgpGGss7FuvN5wKDmVc+80yx7wVwn2bkFENzIiYHeubHAnqnN4NeD
HMdtoHRn6oee2GWmefXYuBR29s4cXcR0iCS34EymCt53dMp7mr7l4k6NSLCD1gAX
dq7kNF2273Uk5lLFnl9KxShNhtJQ9jBEL6JMk8oaUjT9CiHN5vcmlazp2xnhBx9Y
XesOL2KPtnNnCrIWnwe8Z+hliq1JLa0HDmYPcsay+3xyk4+fHQehWnYltEMus4T1
ASPgE0AYsIX+q1TIdVDC7hZxZQCKCu/Tvm3ebVtJ6wa500KYrz4e3sz/OkXFakvF
z3Ma5AF6Zbky4nusgT4GZkExYweu09EM3dgPdybLdQoAvttfJxjThYYETk3hKcEY
ay2rOv3k664cejPT/QjRHIld7OhC+AvVJk+6UPUtJktl5Q+t0lX8wqVRGFrMdH4Q
xnLkN3U75oz7jW1ChJ7YSJdLkG4xGpdpI6E6Ur1XpvDW1Xbo2SXUk1G7pJMfWKvY
GoDFFPaR6C8d6RniBImNX7P+pVLy4wl5h5dd5BYk7HGZl3hdmmXIIsTVafF8Vm9c
bPYj4DPbQiteCwSnhvu6LJPNJK0bDR9L+MbN0zTFqRbYX2J2kVRXGWOAtBLnFl4i
C0Aa7vKW7DmKvv3ru7by0cyoi3FDC8T5g6MKPADSGhpdkWIm3GomyBL1Bp58zDpL
N316PYegvOhEi4leLNfrQsI1VBJ0O1iWmlCJlJbdo4EkVxVf6cVkWGDZjgGB3NTa
xj5AVGEIljzZ8gJzra8UNx2aVK77DP5o7X3UCdun9rd2//Fo8NX5n5COFmT0o/su
qkKOAPeQNKLOBnla9r9/Xh3dL5p3iXVTdpi4Gk4x5mNw3dhbHIT/NQX4424ijOd1
2XanCZHzYM3CKy68PBsWbwqnShFms14Moh372tGn3Vuinuu5c6opFB2DiPZdehyX
zT5B8WC6ZIUMwbM2IvKuYKlZhs8Q9RSKGYcyu83/J7vfTFr+YV44T2PKLxErN7qo
0GiLQZLzNGWQHmwofmrqTn/r0usakX25+JnipCCZJXzdGA/c2aapNvUnD671kso4
OvjbTm2/Ng0AbF19OzyRAMzN8+gMnlCIe0icJ3YwiZpOdJXLjRRSqkE59il+8yzQ
RPFH2yi4rumuidp4ychlrTLyD7JtrMHqMfsSyVOg16E5EBMsyWn1agZKsB3rnknx
d2eIlMbFFXXZIfIOdYFMelsSHjT1FrcNDETfXX7EFWWCcq0d3xn3Xr+pZQTwnh4q
0l17i9KFMMDMycJT5eiJXZ+pojxUwoVbB59c1tBhQEU7g8n9NH5p5Gd6NAXeY8YL
gS9EWIpmD7/SB2wvI9cmbsY0yg3oZsr7QeUSclZAvwIe+owVQSmbaV9vnVjSRThP
LoX1wj26X/QSuPVveZr0rr3UuCqcyFHgaWlqNw9b2bcRVsCuhViea96S1Ww+kUQd
tEq3Rr2C6yYuuTF9kpYnaKGLo/YRLic04arpR1zUJQEIwmY/px9D4RUkS4WQr77y
eCeYpxibqr54gztUkCEmtlmaWlrtZ1X4ecIbSyyNgppXvgUrF7S0Krx6hblQIYh6
UV3LfEpBiM1XWqM9KdRxaqBsVTGva0ESqy2EtjLz7OY6xMWNVeArXod3nsfF1Jmc
tBFUakb7bhtRCwaOXT7eqaL3+PU3OIF/TI6fWcUKgsVRLPumrVJGj+GxdOev9kT1
DNJdLXbmpa5YXV4R01qiqmmdXIE1rpqpcqDYXhaSBLnXDi5IKoQfKYwuTa2uU86k
WQQJN6lUpaolZ67+kElnNgkacirQtj3EG+sX+sPXsNjJwfaaBqZ0chMNtUjG4xAo
faVngyezbtuSdQFe/Y84zhRnA1dy0QVrtlAwiFcSL3hwkj2q4pnuPtqK6MRMetzr
acwCV5e2HOH4bvs4ScXFMucxamc5O3zIhhF4IKvsqvNnah8FMcQTdw0bD5/zWX/h
AaS3oj6YPGUv05h9igwR6INKgXNzoqegJksJWlOWhqUTnAwhEsXr2RCsBxFG6u8Y
SFuc7+zOFhiLaDDnOcRuOHg2SMRQbh+VUTVThCUGEIwUSaEVm9gkJYnLMgVW+lNx
AJagpkX1EQtGKUjqG+2dC62tNQZwgMVhxqZoaUpoB5gYsAJ7xrsFwklddW3RFN/a
IhBQo+iIWWMWnxzEHI7gxfRwRH2CvJRjUhzYb85q/NxxLhF83Q07wqgbHU1YvAmI
DyMrq4QhYCsz+sEPjbtP2g/cMA3nISI2o0Y4Il5vGGizj+0hOFreVp5o9h7OwmIK
moaaMseC9Z4SWLnk6PRQb/nQN875UtDViEHHLnlRl5DgO9mpO/uRLaQncNOyZFam
ZEzfFeaIkucgFiDvowbTgPr3hv10EXszQtaV0KtKNgDvhMgoQlSuEmKlmCWJEGSS
rx8DnJovsbF1IMm4o79EkkmqML7tv9/LrbPld6u5GGRc3A2vVV0qocr/ztrI50uP
yU5Bjjm1Ezo+4pbpFwjYFy5YJRxdrdp3vGZH+uvgEApnPN9ebfjbXaPW85pgFw2f
bO/40B3xft/YaF+qb/ilG31RqPRtzWVYakAGuVOHbdB9r1yoKPNPiY+KgOCb1Xfb
kisvEuxvSF+nRs6xD+QDMsSAbHZ5O7ptsoqwOA/R+BI1C7ZaD7vLK10qoAvMN5J9
tubeHb/32IRwsJUqVKUvgIjmyLElNJQT/Vwts5fcHOObr+JdrUvoXgrO5BWrvhbp
zA7fh+pxMXGnzXRNwSwNfTVgXSgv6xkbkG7qLs1VY8h7rsA7Gq2461AGD65mV4aT
j/J0QZF/PhsYlp+AyaNaPTnLxVBz3lKN9zckVs3SEF7yzKxa5CQfufT8fnsq11Ze
r16kklADah+cJld6Z2oMgsEI3Vp1l0WZs89IHiF3lyZZ5SwOIu2OnNbwRJN+4AUu
eyrD42g7QFPrf/x5dGlPMby9etTrAa2Lv4at2W4DkyMfd+deu3hdgw+e/4kjOpDU
alIlXi1MWFlNghIw33oteH8o8Jd9lTwty7Th1E9+eWhiiYxRPIZKWcuGiHsOgYkU
xgND6sQRbhyh9pGIr7sJgmrYMjxVB79v4DIVLotwwVmteb2GQighB/ngB/VP8Ol6
eKM+wm2TtSWf7sQ0lAOpInq0MHkEoudf+aWQ6yO7xtOV9B8qKl5510QlMihwSXn1
jCSZlP7skryLhpejCvXXd+K3ooNUbY2uhn4benZD1EPufWBf5UoFFaPe6N+a/PS4
vpE8hYSRCbfGEpg+5dzH1elXqX3qrMbmEENaKS0S9hM1Lb0ZjBlLnND1JajDYULV
Imo4H+lS3eIk7HZUYsLo6eMrn0QmKYDWsCUYz4u71dfmXbxymXeozJBe/kzVtZpj
tyk1a4nUz31dxO3jTjkCG2YcCZ+zGQltKu8Yax47UChTjkYu5KHktrA7j4CE3b4H
Riu8b9YQUph9a2fsejZDYwQMvZT27r7Jv9ewH8pNtyCqagmnqj9gAgRN3BgkN3j/
mHg1heTOsW/OGwORgAf/YgeHp0SiyXFdZriyC0FEmjk3FEuyTmli4hFiz8vdi2r/
offnXFYO/3pwTQ5Li65bZVkP/SVCBsr5qqu+n2EGG6V9f8NJaFGvc6yMJrP60vBR
leSeW/wUl8aH1z76SsK+ctjcy2LPnImrB7XiVsLPulsrpi8r3SvqDHcopGhGhff5
ztIMtldJVs8/BkDUW+DvQXQwIpSNBdhDHK+UObG07D31d7tDVPivXXbCWK2MvP3D
c/ndGI9ppIZpCD9rDdKM4RPnqAObceGAj+nsLNuQQN/PjLNabCr/Q9ZZK6pzz5ZQ
jLoMeyHAv/I3TwYsoW78V1Ffs9dR8d5umubfTNOGvQUSzVuGvGEQWcbQ1fjxtMXg
S9T/m6yDX8ti2Us6ADApnpd/woaL9tDB7cGKzKcO8t2j/RMwGJsVcNMVmpZdjy7t
vooLMqpaeLFm1fhc9/PlrVU4Gz48o5Q7xnE1vjoiwkD+w0UD8wbY+EVbtxzqDeWh
svsAVHkwJe/0xrchIF+7nP5B8rJWkuLHTikHNISYppViyGTeVpWjoxfIswVkXafE
79eqzg5bKpSHg0GZhA9O3vk8cYOq5nqZNqEX2uPrt+FUwVT0pFrbXaNZt7G6zfmC
1JZchsXeAWlNmR8W47gulSfBZ0I6fxZmoNV4qyzGsblSiQQIP8bV6zC6eOwwDnmb
J9N2cOaM47NJdVTydTqvxo+qyR5P+SSEt0DbH9GaScp7uDOmK5s6Ey4KP7h4kyhi
Ku54FefTWpHERRvk/TvAcdUBULj6ds51AIfrJ9Bx3z+488Kw7n+oDkLsCIEpdPAu
nBHUolFuGFMPpkYenBjTjkowam51BBtjhCAIvJ7tOxjIbtDXDiQNSzGJVkmy1DlO
I68iHRNjxFjYEyH5GFF65QxpCn7hYymlBifgKOF7jPP7UTcMhXpEifS1kL9WS8fO
wuZ0wHoCUS4ss5yp2E8D1VcUcPyHOdbNyT7WDVT11hs4iX008jEYuBxNjIGPtV9+
xAKs/sd5uEzgYkhVaGo98gQjKJiMaKQR3a2dF5zd/hpylg/e5M6tW38pix4b9OPf
RZLECYxcWYsGbAJ4I5EjM4IGRc4VvoxyziozBEs783S4xNLVtR0DLVoizD9EziUt
rrr+rZSRJLzjvOdl08Kk7hGgWUMMaNWBemqgqAvMqPdwCCteNqvYmVphoROohRYs
mtSHVxTIyXO18VRWX7ClyB1LU1zu4nzf6d9ahcJzO33XSLh5u/ApKQ1GXHo8R4RC
Bpnxsw58OYsm6+vFn89WnKr7c/mY3CewSy6f9kWBgTGaXfmI9MkiRmxy1fbwqTHe
I6lw2l0dJTJVPQDZpeM55w/oeasw7MAAzXRZy+6UfhIpf2EXEGihiYp2ZaBPAQTf
2+oDf7xw68CFSeJslxzQEPgfTVOyZ3ZVq9/w++llGjmeZa+3tQVq6lGW2N8//Vx8
CtXmbOHyph2L7rJd9dmKxGvQo3WShyHFvK9u7AMzJzE8mEFnaILvl5ZI6Hhdjsna
tVBJpsM+m4VCFgBc0IM6oCit+x6b8y891Rg7SII3gV1Tal2WDNrVSfbfR1LD3RCF
8zWkHZR2H7RITElg031W/eMxK4iB6IwrwFMI4jAv9se8kTRtVAex/+FrUW1ytyS8
Frt6X9sqQMDUeNehVkatnQAnpkJIHXvDdma2jPXhIQvNt12a9a61YGZXrZBN7vf/
YzY4hyXrdlR9GyxPd7EvRrEejuS2Q+sN3H//lCUY1Id10JZaw42604GrkMLOFNNw
NrhPjlrwmCyYb/Eay01Vnp6IlHEaBWfs9o0g7oStSr+kP1s/61ShWVf+nsdjMzsi
xr+8DGGbhr46GHDMU6TtuXItWPMXbZy2H5dkbYbX2YGTUn0j9+OVRB86hrFoifY0
GHvzi0Ik6P7mjL9NorWs/P+R8hEZsN71fAuT296x+ONFpLeq4+3AIdJWkI0o2CrM
YX1FsXav6hfpeRATxgTtn8k5yVWjgXkXhv7/c8+ShuJqOYk0JtPNEqkj4aZb+2jq
2utXA+OcSUd0jxLy4rvmnV5g9EFhR3ZH0vFPCU1U3bI7Ng9XnTfwIEBANDIlUn6J
ij2sTht6QbN6mtdnFdFFNlIGL9N66+98PsQSf2CydYhtHPqjzo5LnmCHZUeZODuR
2/xbJ8uFX2wfvh5Mn33p4cwKBDBKCqaZ9sxjXfGzaqXCI1f9RYC6ro4jYK8nhxn2
dWgbHhlCf6xkFLSKc30jdDXF/RXem9B1CRJ8ssA/pp7VP4R2ItAx5JEcX38QHGay
CMY4hIgULVdb9Ta+qC33Phk2SLKMN1c6teDEg///YzzTHBcrDGi+DLqOvEwJR6b+
atnGpzs5PplygMLcTPXmVgss4DtKWjkRSab9OkmGgBMpPNKv4maEgcm4k7/cCRx1
BHnIG/waIvpwPPEChaL9VCXKJEXKdV45TaMnE+D//pvWG9Lxr54Gob2NfL3oKWbt
vF7SBsUl0UkYdX1EP8aHTGIgGtNsoi2cSpXsypCykEP2f5F0iJg2ZdlH4Vq1Q2Zo
B/A1QkQu7mU9GFDJwPvXyENNptleklgTvHWowahpWTZvAGBx546C0kWD3LQIpH3X
MSS+npynD4/KVZPaCxAq3orzHMTYi7QoERCqVlLAOvYMSQEpGIxLl38g18nOeYOO
qQSwPHEGhlCAPi+fP+xY5lokDZMmQazzConyv4MzxlLurd0kpVOvldom37YBg6b6
YxupazWQoqWGF6se+wsp9UP7CrlD+8vjXXQZeGgxzaQ8leZS8Cj1R9h4lR/Izvym
NvysrXLm8pRQOcN4kfPljhHxatAtQX1ngj8s3fLlyLDwWxuRmQ1/CElKY5Pl0Igv
ayYqBjyTh/dFNq6ZaBgqba7pFgJKX14ED6NTiV3+jN/h8rMbOi5GXRY3qZ6e7+Zl
HLw3gYsMZupdgESONUPvmh+sbnseFlS1C5NhTc6cso9AlJGZOHUwmnlq0qvbPmSv
A3ISlunM+Mhoxca03L8AjX6VWcUP913OH92+0WpfoYbuvqTtWZGWlqMtq/hEtxqJ
xEH5lFYFZdzYjet7a3aqjc01qVwMa8JMRqirH6PJzcc0uCIWvIyKpdfGqSvZL2Et
4kZGTE0k7e58/gkHLAx0cL3VJ0avG9q34gRkSohLCP0zDTqWlIwbTM8OJapy2OTy
pJcMZ0eY3dg+7iNk0W4zrS9TEq9o5NWw9Q5RlgGtl0X6RzbOAiuva0TKtAC4S/3A
41+wO9Cy7GLsH5jkcM8RNNy9j2ECbtrv/2IlfZ8BO09X6xYgcIvxb0peSUQjKrRY
G4a2wAdZXXZU7FoIFxOYePyzIIvFcg/tj4AMXvrtZs9HABIZ+YDcroXP7MUPKjqL
Scy5LeUKJq9+MfEJf6LoHEvEvRUlkhvQ6TACsOzj00uadiCEbJiswdBC1z8Y20dJ
LWk/DWc5hNZjFqAGo3HZBeoAE+friQPSFUjJI789AYMDPSoG75XbaExyE6IlHc8z
fq7aDQ/mOiFR5NYK8uIkGktKj1LR2hjGhvhE+PORw+7CjzDeW4WVy2YJAEeXEA8F
1PC0Q0z8knmbNk5MhVH1xNK3BQUp1QsyQU5AMZvRtwvss6/cnV+WW47rJfXX21XP
ypU4LVbWXMRTZH3WBxF/h0iPczZhErdioHtI9ZHAPOHxfoJCNj39WK54W+l4ATZF
r0KqjsCcgk0Gl6nOSb7P/Rk1betTxKQOHNJXVerH3O3J/z3lmZ0EGuM4aUlXmab8
2/X8vTNvllJ0YZBKF4yjb+RiFCM99kaL0P0Qm8adjj5lvmHcZnLiFBALlpMiUyUU
LyX5ziCtYnUSrKWORFiKXRnFcCgNKE0uEvGmIPMI+y8hwFjvrb8grhmEXLySF4ku
7VAB4A/MLUZ4UFhh8sfBRjN7a7qRzGVfs9AunoEAJ2qC9qLcj3zh5SEZ08k3biVU
DKmuKqfBESvIT/qflGzpvYfW+ESvz2nXQThVqC4dJvzZrD29uCLgkH4kxGiV4AF+
1wY/2YMOKF4E7dQaI/YSUqT2RUkT5XxEFzk4I+umsNyrKGfNdW252WvgiKnX+PYE
FPu6nHwhJf58Sn++ajT2PdBZEkJO3tJM/beIuXT5U49j7dk+92VDrwfirsB7X3I7
Yrf7dbtpDsoG0CudTsJFu8/I3ReFcFvPdyv7nyjOKsheUPFZLJvp9zYZYEG/2Foi
1xE6F3SuiCpZZ0cXvJPvgx/9OA6EaXbyORWr7q466nBlFncw+5ie67Tram6Jy6kM
36U8PfyZjgz740dsJhaVWZm7Ks0VphEP2Fua6Z83SOsEryqfjyrG4YQu0fFBZ/yx
1U34KIraaAeRGb2YOcEt7rsmYcB9sGYAatcCoGVq61HWbzvegdE0SgnsB4i82ZYx
6JFgmOtNMJ9yErfkJ8RhoLp8LJmT5cN57i/6IGdHz+lfmnYcAclFoYdgKWBGu6eO
4LBxX6GlNdvGz1bT5XZb2lTpi9Pj9p1FKPQ3tOUYbhJcarTT5dCUx/3tbIcxHb9n
ecHkgHYHdXTLhSOSEqRgz3vIeOKeyQiUn5Aa6qou3ymze5TnjULw1+p7ckWx2ynF
tzOv8w8kHCNb6miMCuxtE5HfNrbI7zWko2jVq0RDKlMroyvEFbLhDipdhmhtMoJo
z8GwDTs5pvqmCXh7UuDuyCiXw6oT5Ux6n+64ArsZ/ZhHezfAb9KepZ+G4YSQpYg3
EeQuKlMEpFQ/7QfjnxL6UM7i5P/75XHUKH4ExR7r91m5AK8aSCBT2ZMlVq5Pda8O
Cxk82wsiz32IpS6a7bZmXodhecTxgQJtCdKl38qXgqaqeLINdXFK7Wh92UW7Q+yH
3V7beKoRbsR3WdMLLJHT5ndXmzA2ZdMJq2lKEqdpXHajwvM/3j+tJM51ekBu/G4C
B+j39SUYl3CtaYXSaY/ky9YX9I4MtjGCNjczIeg8EH6zy3uhkcAKfrDR77pM13fh
AkEPK97o0fiz5ydqgqW9LQTAVu5E11NFqjmFglwHt+JcYZuqJ525m47ZZZ35l4Qz
MRBofQVS8a86tss06jWNW5pWBPHTd5AR+gaGxRIXh3MvCFVX5v5dEkmWYNajo8y/
89W8N/0X0CQQBxkVP5oN0nwaLLtQyTNvYmeWoyyVoG+5I5ivOJx+mV4iXtNNRl6C
CcUP5wt5ZrZ6cONklnhX32CJoQH1MHAx0fsHAvu5f309oqVYNkI9HyNed/KRQwSk
//2Iz55NqcVeA/LH6jfTdXzyVJaRg9nvzpXw0TdsSNulsepI+B28nnRkaln69SrZ
ikMoN3/junQg44HSwrmwFvhBRgR5AulF37ec4MTdKWYub3iEgxvHaHMOqGq7jyEr
aPs86dIeVZcvrU0pECjbRot27nU0/Ex68XfVZXMs0qXE2K7N4/jofSdi032J2oBN
I5V4wClIRHuCEhYqK9xGtTteFmCbwRSS3ShscJcPMYrZkpbGeHSPwXSdrLT67Sg/
N0QGez0uKGX0VBG4PQyw69TV1JifcLaAZg8MBM1CiODmrQNmF8MTSBk1JF7f592b
q95FrGwPD0F+Yorn428t7/rHW+8M6eYalQ85bz7nG4wfXbpBacHDnVGOeI0Erp/z
Odx7wD53zrrCJNCY4m+Q8dj8gaL70B0h2DBQmv6IT8SbbH3fk6NAvMHoYb+K8HtC
d/5JWZkAV6hVW9ij4QPI4WiXIlRo+5QnoIly3sNQzrFMzK8oLy/tY2AOa+/35HL6
07xPnRMUQcno/zJ5k8+7B4JLTIajsjNbbeXoWFKtgXzlWztmKAV9wu6ug329+HLd
hDfolMD8dADLJC4p1aGenQ8RP3/29TB5qNKPKXdg8SCuKREaFouTgUQ34vHd8fwh
6IuJasg4Zq039HrhLYl+VsA+qMFBKitd2f0Xe0PktB/K5FjiCAvz6UPU7URkZw/i
aytW8nUY26Rlhq+j2g3P03hxhQczXQqJwRmzlVvA0dLsGQQXPvunk8pa5DYd/1DT
0G9GEbOO9kK+Q/XyBGmoo36/A2iKWfmfZOqI9eRxJz27Q5K8P08Ok5QL3nMXLA4L
3za4ehr4kIEkLWT7AbzipaIqXrhqtQoB8wqbgh1oY7sL/6M5GDoHiJdq3WT/jz1T
UlNhH2DIhqGKt2rCrhMVIlzNY7CHYJJe6TzwjtZB5Yh/9CI/Y9ko5SbiEfNWDiA5
ouumijcUnfcUzcnoxjD/qJpLAub7jdn9nqM7yaC02EZhM01AnPOmr4+DutCfiLmy
5ASVtADlQBNWd4QR4prB4rN677f6Vxdd+38gPI0vgzxT7mGZqK0rEt/0QVS1DpGw
Czg93tP8hSt5UrzCjbtVfyU+cuDWm/zkeaUHEYLF7P7+dcu3f83o9b+xNCPCTNiW
+ampEoro3++zobIS5cgjWIJBXl/ur9hCi5Qc7DpcKNhbnisY/WunUaoU/zNz2uaa
GnZkiXjt5DRs/bur696pvXSO4zwOMqt8OqhrRQ/Ek3Eo0JuIkiPodnR4sEKziVbO
ek5HIWAFntAJQRzhyXNG9GVRINJmCoqw7K0DllFUV9KJytNxcIXTGFX5NMZ4wrIb
NLu2+r8YraRPXFFybtGw4JL5BkYA9huRnmfmtH7GPyKDGJyY8mHRcK1UWCq+J4EW
/u/sv568Fdf7RXhjB0z5PItQwLx7PG7bJzUnUbTM9dMtjdD8aG98jvmkTBuLUbDj
UFhmZvg5WHounKQpvtiT6ZrOlnVgvF2SBU6tmAJf+fYU2/bjjA/U6VCQjSZp/kDl
Kd/CB0WXDlGa5eNYTELLi17VZEyi4571kt7X7AAt4TfHirWqQwrr/wPJIpvqvUYn
BiVm61K+sZrwmjunjr7D07hwMxJsQlPIBLzLUxfbhECcLGgU/rEAbfmb8yRHmXxa
tsXorXo29PHwCkeMmOD3ylCZVtQRDwhWjecCim0Tr9wK453Aw+p/5yLD10wc19yk
D9KSLBmyFx3K85BhXFdh0L0rmpxH2AaP5eDtrhObWl5ewxDUewYmYPn17Tu/Em1X
sIuOojGu0o4VqPrkxj/a1+28j6K6E4pntZ6A1zadGBFfI60YTeGMSan0dKflcO+3
4w7tXbQPszoSMAUi8bhpTCETv2eqiJJjE+7YpT3oZWaWfMatlb7dM492JcWHaHe7
lanaj5WZ1x2T5uiTtdwLMrjuFY1gn2oR9ysxqRUNfkMii2Io9D6UJ9M8Vur8Gqcr
zKEIpml4rAm9PeP6TWpkTP6p55JmLRVcVx1KmCdKwc2SBGL/eQVc0AA4CX51oFMp
myZ3vm0oV+sJhJdZeG+ABGZeYQhaa2ChGzlNupR3MGiccFNDMQtFqFytSOH6b5aP
REr/guDtiM2aTXcqvlxV7ZnsdxzOAM/feczSDnjIGcu/g8dOuIcCAIGGcbRvJYUy
xtPdgj6mHeZEEMGT5dxo9I3e/LafVvIuK6nW0SEZGARBbm0iNf3om4TMfP+OVczD
tkbhPiGSGedAStqldSxTtTQPJbB/32X0+rmz47DU1kcsVr08tlMto5B97g6G5rfW
hzbByW205g3xzkTsth/KNnZCpHZZm+TAXJ8iHccYGoR6gajIzEmjTMSQUjZOfMt0
LWqr/7Ic4YC1+tL+kXNyICWw5EZfNLoyTm8JqX7yTzMmsrqb352H06avYKc5XXU5
Gf3QfgkwuE8TYtX3r3GdH5cCHNdTgLY1Z+kiVn5IlvbCZVJc4M9hj4tZPA/L36/G
6JBc/xMRsNiLw2hFi2BoAkETRo6mLfrqZIBBi8oYPqQfjkUoCHH28evD7ZQUWgQY
F2mrc4AJS+sSKiFOS3Mx2uDhtphrfUBAJ4gRN/2DSVtAZLguSmqH7r8ch7o1wQP8
M3iJdzq51cag/6IyWLVaTfaLukWH83meN1zMxg7tsBq3qLhiRa1JGi3j1mR505Zn
1j7oIhxEmGjXyIgXdMpxLLYM5glIgx4XBV3IlkzOxnD8hYAsYjzDepmOrdyLHGOz
Fz4jJRCL1bHNpvFVrftE6SkCE6N9ka6lMQLUI8pbqBEGQCxzLPZcuQkVeeUip19U
hYWpDyj18pIRYzEuthBOgnPGGOzSafWzsro1FZdzCPL7lVuAi7wT+s5Ov0K+KPnp
P3pTM9eWf1lIffGnLOo3mpGv+pfI7n0Ei6tkNQPnDfNIlJcddIbRq0aMpybnzgD+
Ph1z2Zvytf4VXnx4ZHVvZM+ZkJ5zsn+gtyrnSV+82F2ZjcQDKnf2B1MT9JbDHulB
pFQsJyzrU81P8dpYxqecIu5OxiLWgPsyHyKqpVDIVDC8cXBiDNtAJS94CdDxTNIB
Iwpbw1KJNHeXEbg0xfWloyjMtgT3BBBFFvxtfLIh4UNcxF3bqJmnm91q0A+fnUy1
JVV3yrRkgIRjUsfGkRzHzsFPYo7hj3bz3KA5YVinycpsQuZH3dxcO8t6DVYAlCEc
UOK8VOb8/BVZMdQBdTWtfna3Sshyv4wIvmJVoO0Z3oPzcIWMU0XVc+XsxcNsjIYo
KMr1r0LJBVnP/EmnI71CaPdfM4tQVuJlwreosyqUtIH4R34NV1qo6+8OkjCiOBt4
BbsfhwS3BIK3nsjH2V4/NfWRMbHfxeavr/VceutQFjBLpQ5ih2Ja8HH0SCNSjEmC
DNOU2GFgUJ+93fXgS8bpMVRFV8ZO9tbWCZt3iadF8uwxhhM2GwG7Fhw4cNMaKpNe
/me/Z6E5uk0sR9T0L0yzg0aG2eMxAAzlj+XrgF0lXW5ZFxr0IhdrP0qzzC1vfroD
fNVBiZarWg9bRLyh0LwlpVRpdu7CiQlqXwS+Cpeh77+MCJBYiUFvfXX8NgCovFOK
uF66lAYVjebDBHUwt9aZNCmY0MvPj05t2f6gUxo8LxREg6XoHvxssT9hBBSpcX7z
LHxpOCRQOX4rpg7/ET6ZkyBVsvPr8UI5G7W5/ha0Z3AnPub1pmxphn9ZQPj10Isg
samUNwcwywDXZXpBq/XD+r8gvftSqBLbCd1KURotB9rUwTgI8eeszHTIX2rieR+z
lYA/eY7h4vU7NuRwuUrEjermVg1oEQsHzWVmJ+RGg/uKpfUBjM/SVJHWkhzKomeM
MBADihsg5vLGZx65ciCmIFhMO2T2L9ef5hDzFjPxWrMnNKcMjbPru+Ched9o6oDJ
GnOlyHf7vh7g4CatTJSBW94PQ8j/NukHmJcwbOQz39xNEvoeq/vthsrC91xnc8F9
F5PaDOCu/1aiCE+nA44Y3CPvKD13nvATeOL0M54g7Ilg8l7EXd+06pOvvR66alYk
gkUQBQR8qryS4oRBYL6SjM43HWsDiQElYcW+E7oKyW+yO/xKZ+qC/or/Q+2kJ2+F
4zStjZeTicBvbpfkew51dryUAwtmDbLVAC1A2XcCBRyB1X/qktue7Rxdefm0gdC9
0eBNM/k3ZBRYr+TQ3AsaAj6mhQ7b6N0nndY/TUzsIg3jolFi3SKorlMz8VImaEkH
KC2DXej222uNNYr6VS2XscxSNnaxe3kiJrhorufOc71uAeejeTG1OXYiYYtb5nO1
uRPlU6hq2YyIfA28tW5hxYmY4gTzWlwlO8vs62PhR7CvYgHclecZfuHS700m8h6A
wvrYjC18soT8fQJgO4zEfo/VnZ/x/up8eFpynLVUOBWL7nPMILLxDnJx6MH3aUCE
LMrFeoRvDof62+lepoNOZzkwRD6cAEvKcG5lj0T1noQPKLoQiQvv8iorPEGmnyv7
VhVPbqJehJiZpBgjr6iATeywKxusoHNouiu7MfNtS7iPmuRmOgdCFm/jINIgctbT
O+jgZm6xTzJP2tXpC0Ske3ENdJ5OCemR38MqWELmflQY90nSl2es7lUVijiMsoQW
6URMSXTizCXnuu+sqda8+YdyHIBaXFL3uHP/i1vawZtFhkGg5lANBkgJXy2nDdLE
wtZOf482bsDvTdqmI7JZ9SrBuJENcJe0bVgRdjccZ224r5FF6NDHd7Zvc+QZEl9O
k7y2aAXQyQo9RqWuUhvZfAnaM6AiY0RfDzQ+0HZSChBdn6Z59PsWdjm5F4NL7Jxe
vTekXgxpdmd1bL8metXbBWnwEx/FsRNW5Bu/1CngDwH+XjlfGK/xT5mJkKyx/Wjy
mMnDB0Uu/OltvDwKLGVkcZ1V0N7NITjXYaBeuXndsASWsIwpoNU9f9duNXMJ4Dbq
hBxLOMug5mr7NzI9C5KQAY5oFXu84Y9dJ89CPS1jwzmbtZU4Esj+qCRQuBXC4/zz
Cyr6BEEK4DFCEeF5JQS3vM2u6OH6GivkUGidD1D2cXVNZ2gV9neFEB/4dFoq/Cl4
8w6fc4E6X9ElVeqxLENVVCqspweCEWcZTuow0g/A86GqT0EbGwGpvnv9RQktgEru
uy7EjBpJmbaOzTXWy/bumW2J58VuPTTi67u2O4o102TqeJVcGCsuf70bI/8E/CNA
eeoH6zSktp2cBtjol9E8AMh3W5/O/8aZzYGGx5iBtGaXUca56QVE7uAlBIhRmBsl
ahRusH8UvLVSp5UbUlukEXdMmXUSgU3cPF4XftCd74aO8UXCMi9A6+34GXP5yGUi
DbOpZxUAXno78UGZZQInFd+6JzqG5HYuCVAGaxmcCyXwPCPKbutfjYm/JOw8wVEu
LjChknw8TiI28y7fDrvpn8c/f8k8eQo0btRqYyL7CJwuZYavLMB/eCgRfMnksVJx
7VuddEtQggFbuVzfX5ss30GC4fWzei+1BgKtlZtqNCZF6P2mFOzWHtrB4r2jdN9x
3RvmLt/1isFjUMI8FnJ2OtBw4KGKxsSiLtf7GTZgB7e153hSrnIpqo4mCUoInBft
lvvyA3/GESwoYhWdjgR5ku9+ITdVL1kbGrbMt7ZQ73+NwtlNPMvXcLSpvYQHdQaH
ZvDDNcYPPNotkm0kLEz08VDVJqF+OA1AemDyHmXU4b24x3UHEJzC0c2RifT1F35U
XGP7ttlEpwdtG9i54qCxcF/2jeGp/0pr7Q3U9rVeN8ZrIZO/nK+7B0sQoS9JVJEx
Wz7ipXq/9fUjWBj/pbhw6EyTOMvbU61mq+PVEp9XC+S4deefnFol2GYDN3W+NVwO
az3KPdl9dHIVgCE9XbUOVWxDRqVhp1Y129uaa1kR9GkmziEaLmHFcfZX3ice8kDW
LJ0VSfIzEDIjn0kbIj7neWjrX4K6majzekrK9dK5dBl4AZ8S/cPyt4G/2Ocg8Dj4
fICR733ObiT/1IBafQBgJRWaQ0+2RGLZEqkrwIfkzi8q9sbRExjs9DDKtxsnGPIo
F+MaHinF3TnniGMc1OqZ2CBQ8O1FjCSaNwTMyKxSGPgq3G2NLO9A/BLs1WgrEmuE
vgmGW3NcgyEfgODdZ2S0HOYojszmZkHz738dj9gpbo5c2I6p1ityBX28fLquUsj7
1vNq6Jd2RVgXSXVdnWPs0hKgm6jdPiF1v7cWlx5QEq0gwROCve9NHfgxBZbK2EV4
05JXrioNq/d1ZkZxYEgTHeRWpWypTtfkbzFKGvHb3BWjPBieKHg0pE/r7OcxD326
GMuEhbt58lzyTEhnvWlK8kwU9cimBfobkW92hb4rMkBOIj0XV1PBII2tJ7S+LkTo
HEPRz67yuB6XxsCZvsd0vOirIMlWMsjzsVggWKuhh9ibnsHmWJac8mMMwR8QA/m8
gnpLbvT4BY0dnou672x5U+VlCiip5VZ2jenRabQAVctR19bnkpNttqHpLF9pCXPf
pASCCKVK3c2g+P2WhL5e/IbtiE8aIkmeY91/P3SNgdD75qUJnAtjvDk1qZoyjilK
WM7Aud9OpaFE4UAEvrG71XqXtq2J0WlNmmVQ5qNA+NOxK5kQ5dhR7SH0kSnV8y4T
Moz2F9639Ix+NLasvQ+hFQlJxoypFIjFMh3A9t3BYOC6WyM6t/AKJJz5jxI7q3sn
13AoQ50o4nvzPQoATE30IDPttxjlQdrWynVmvUcAx4/lcTA9IfuIU2azqbMSSzSQ
vFhW7RtyJtToS996IAsmK6aF6g+GokMS+6z60EjXekJykbBLt1a9ywQsXGbmwOAZ
vAtkG5TxizpeczWcd0Kpk0H4j3wW5gYbrolE2J6fYodHrqyAtfnLO065pl3d8bVL
lb+ZjqROeYitIbI/hUXk11M6aDpNDiy7fu1aBX0j9y3P2znwX/iqwjYtm6sAkEVq
2Rnj6bo2+fW5Upi/gN7XOTuHJuw6UMBhdN9CC8PseIssc4w2yxJ4gJFu9KJVV+UM
9VtCd3CAPa+ChpGefIH3BEq9kiNV8G9IIJKu4HN5ssBC9owHKU3YBFpwLur4hehS
l6XWqlAIfhC0G4k/bocdHRsObjpqGu8QNYsSwcg5nHB++Z6FomKgwaP2aRP8/uiF
KWitY3Kew4Pj+TQOSUa1/PR5BD4XWdES9aZWpQg85nsI5qbaPBAV9TwfP+lXcVrs
aXrO+dY4qNlhA6GmEcHUT3sw1VFN0q/urXd5aTS4wwmxAclWX96axu1usU6yFgaP
/Ll/agJ/qUsn1jwYzcogGmZSts0X+5khaTX5ZKvlXLvQ3NULOblDM0kfuMxdDqrO
5RrUYafk2N6zILFYTjbIlUYoQL2rX9QYL9xwPsdKF0xPyt7OAOI2sSgi2WJx7Q7Y
T/Lpo9LIvxOuS6Lr0vL0vMlg7noG+tvfyxD20pXk+5H7dUhBN3rbdr0sylS/dNAc
LJq0I5ktgzynyMzA3vEPo4hbzYBzg04xjLskiSiy/gZTWueBTSN0DqMSmLt/hA8+
EvmJ/codbw4Sds8256bWY6WzePxFo7sv6elDGcojR8IJalIbVDHK2i6eAXbFxaYN
et4ISX7+UDaaEJ0euwLjBXDeuiL1lDeU/t0zr9GL+Io8ETLEFL9dACGEXW+JiuKS
Z4siNgQJT8DsxxbACPwy9DfDoogYhXmj7gQ/8uJsmthy3qEqSGMm6z8QgezrnYiU
yuv8mu2unYEGkSda8QPHnfA+eG2F/DJvMZ/xxPgukojLMhw1jQ09ku93/gw4A+DG
C6G5hYYrY05Lklnoohvv8YVa2R7Q1b0qMqJGDQ2MZRRIRDYLgn2Am197PqeuOUkr
7veMcb9rDNoKRfjRpUWEfP4EdHgq4sVhMd2oKPUFxbM0B9P3qpvBGcVLaW54t17Q
X1khpVA32HjSOjP8jCYGTonbvdg3WqGxmfh+MfAI2bKoHmiuZT1A1oM/4sd1AnZL
Y3/UYVLQW6+XC3JDEDBmf1MyZEWxdnCpwrTunwCijcHzu3MbwEQ9+2BWnmUnZ+Im
1DazXGza4bEnia3Jr7vUBcoazqm6qcstyhH6gs7TkH4u5MNFkO9VSBMf/W5fItAM
7lRBbzuEEbqs/puPta4+5BnOD6SLw5ooh8Vwq9IYPJwy0GsXRZ5rQ29sCi7HMEGV
CGzGV7IweGUSmGfGZdRCd+S4nrwpmX+SPlytr8oe8Wi/V47KBAz/o62bDG6NoGmO
Cwlo8D1sV6HhO75fGPSHv+hOVbPBzIHxa5MgmXOkrYjWbVshjUmuHJ1iFDGAMNtm
+NiHDDeLYVJdxLUtP1yQENP5poWZYMmxtSd3cGyDWhMWuo2h4z4hHtJPKeIhBjNc
JbsePKv+pl86PYZgOzU+ftID/uqZladPNUoKmhVpBMK1qPr47K1laRZp6fxVbZM7
Iq84fgkhsL2rhMsXjqkdFsGvA+yWTc4+5d3frzjXYOEgvm6m8incSMSmvJGLRLPa
ovAkOSmNaVju/VH26dfBSlmhvtYkrHOayfleqKz3C7hbh171rXNn33lfSPNoXk/J
kXTUSWcclPdh3oTfmU8rQaLaWhf8ieGBmBTyww7kqUodQ/lV9ns9AIeSbwJeHoAd
grDUDEUp2CY1k/9IBwrajICwT+5Oudypu4mEMeTw94yC3d11WKFQ81bz5LvNKFN/
E7R2eOLy0aI0/QGbMkgcznIJV193OUaZHK5e2S40gJk7WlL//QXYgQx0tj5v+1gD
Filjs4O4nqVMK3H4jBgi5M6uz6GICObOzzoRMN2Tq8jqciBrL/HPR30wqwU1rhyB
t1Gh+pN3lFOnimA0a9wXfEuxG8BFR5eOhRZ+nH3Bd09YJMBb7Cx2urD/4N42VahU
TTJd2Yk2viir5o513nANnapg8lowQipd+V2+fEvJL+pfEXlByIdJfuPGjxDdgPvk
Nqe269q/O9ZPKKBK05jk5u6ESS5i45fAtduOEiDZcnvDwzW4fN9Eip8xdYupANds
jLF1oPSlshufZdvMKOMCnQ2EMEKdL5V1dQS27T2FdfIxZ1Gy/cBI1juKq7XSmCHo
WWOIeLo6efVpANRhYrGOYbURHDPYS+c1EJB9OCI46B4HJaUMoK+L3kDDaNEn+jNG
FjP5QTfu5GTU89+IjT7bxSDgYXhOQOWQ5P/edHyRhTauY3Ax71LwoNJEVskBXwFo
jalODq/hapGqkNjDOsCP+OIfMWY5XuG1znB7jTMrYSn5JeWD41EzvHgJc0E89lOm
53DhNQT0kp2kGnO7FoM0nRiBnm24QZapovSHnqehlNACisMd0+D9rmyye8G/PF9k
TmfHSm3dTZtfzK1htW0weAU/8dVWVbMJDNQAJ/nZGagNj38dB+Pl3Vu/0Wdxqb+T
e4wQVWG2ny7fFLrqhhF+yTfnOupLKo2ACevFkFBQ5nXFzePfUFdMn2cczBkQeRaN
/4gCg+5HGRNxeDCrZgKFV2jjsMBpa4ewgyVuQ1HPSVzwUHOD5weMoNwE5rx2kZ/4
Q/C7slz0ym9x6JFwH7/kYs0clGqRKah3kL7tHUdXnLpcsFkr0XPuk3lfAaev6W/m
n6bD0R97yp5Jp7EWMvfcQYukChI2s96jvbGkk5LTue534YZXZd5nW0AbWtIdnT9p
H48sJm/OBpwBAydw1zpfIOqNW7NPzjJsi+5PtoVJoX7K+mQ4fkYUzAFPuCuIW/BV
VQDhjc0WsYdoxKo1Aij24EPbvvQM5FvfEXWb3v1bC+uGsTynKKaRkOYbDAGKro1c
L2GoGYkATpaRVegmZncIAKFZJv6ygCleknKaUeRcyuiBKB7cmGitj486ogayGevg
/iJL5IRIUJKWIP+uA70srajBpjxXDzzd0pUXue70FrzEPe3ThV4lWkvzyfafENul
5PGXhrfFXZfQ/ddKDVg0OSFgzuDKvTQsGUYZv1Z8Un56hyll0r4vxEVvvZL8qEWJ
Etgat2UG/Lk6oYAx6yXGbqcyHw++KTVuB4GbA+snBqumqzVsNxWBwKWTnQtArxyb
ZCrOWhEnwPq3sKkIDIWyiIeocZCoROSzX5Xa1NK6mzDo2OJSg6nEAUO0xNA39N88
dgAQt96HN/aoo5CMJspjTSJERoTRbQXGfInXgeiN/t9vRzC/0GjdH2svivtURUtb
kW+QL7/5LjW2cRqo0Gr2OJZwSK4FKKg38uEGXYx0VuCPU2dIVC+AmGyTS1fMs7qu
prucIRsTXEjOy+iZzcqwz5DQUzwUrdyTAdB0tr9jN7X1itLu4peaWXsTjaLN469J
K5KlzoeDfbsHGu/NgkjHsNRQMyJwfjUKdhx9vRSBDWpGkgkUeVsvrF08HVay8BA4
BNYhJtQ/1jFmgB/mT4ah51BK5AzxAPpCWLvHtpDwHpM3feJ6y+Xir1lRdBYa/+/G
9nbJlI2n4C5jzazBpjej3aFqM+Jvl1Kuzc2QSxHi6pJCVyoeiq2AfTfAJfHsgJ5q
XUPo63WKEKeaRjGJ/ZgH3ywzQ283K8hQOWG1OkCjvnxyEqrCKvu541V+k9K7M1gR
sETyBZMUxpbCd0Fyyj5jLCGx4VC8FF5slnOPZngU+uGRBtzaEnmcTnKQhFGwhYT7
puWIBgHZ5cjqsqmoTnq/pmL6lq5F+S6i4ZpGVzvfyBM6gKu0DTZ80Y+UrkLnQPze
ZxZzyUruPY8ukZs0Bo1nDZ5e+Iua7o7Ybyakqzcl87aquiIqXXVeldH1JdG1pSpp
h8stX1JInJf4CZR3nNSdEJgioauQ/d84cKVRbStyQkBCwHp6xbdiEgh97Z3RlYzV
QFPgFrWKIRGjKuBKmNFxIUNJrLaIQx7Mp6d/yctbaqow8cosrzcg9/W44UfUzJZ+
59/jEtKx7K21DVuwOHhl8YlCON4XeLMVxPEkbRypFev083C1oVH+bDYPxY/ip5kp
MvEQmLRCj448JDPqnHJLDy8ldkSiTEAUD/ZuPVV6wbn8LF1a9FLo2P0KqVvXY5fq
4xaQUaE61Y/LPscN17Mh6g==
`protect END_PROTECTED
