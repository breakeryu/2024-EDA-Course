`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDeWLP7QHcS4/koyjIFVHLP6w0g/5msTlfp61cR2FH68TUZjGoKUMLoL9tjPvpoK
F9C7DSS1cImDPAbRJ5kDTmpGrjmPcrd7EosB4/VjjTu8/Fj+kpYYMzHORaZuWvby
eP5edGnYl1Wndz0dFaKTfN0cuhXg/xpMt9jD8XT8zXQ=
`protect END_PROTECTED
