`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SC63Fr2jXnrz6jsiGGRZHBKX6qy+k07OykrEqCZV5Ed96tTIgPIwbcOP7uHnf1RD
AkUEAnWg00Jg5sciro3QQ+W7ZJmWW9uZWigwo/Mhq6nErb/eWGLT9cDKWd3yX8jA
5E1ayVGqruL9pqlgkTxZBkh3z2Sik9xGRzkD9epSgCp4hNPm4FmdFFBjFIPyFjVl
xZee2Sg4MA2rJ7/BHJ0VdLeASUkR9/wT61xzJ4kEo2MBy1cHvuqQLf+vmyvQpBLR
RIkrkjgw0QHQZeJ4Kqvi7TjNUAzsrZGO7vF0oj1DkMDx61cpsBi1JqKA4xpkM+J5
MdTjJ2+/26M+qQtdqpJ9tiXJe6dgesHCliTI2QtJSxplK/iHm2aBDjqZFnZl0CBb
4Ihq8PBAKmbBJOJLJIzEYvRvcYr7I3mkVSqsZIgy7ezf7sqb/zhAsp8c/uU3SWj3
NPVqRwlAjsJA4v75W2FixLv5VmHWQh1cIMthdKtthnND6S25Gam43Z7zamfKlgG6
YUBq/CTXCvPEWRdGpLy0fiZNF87B8e4FrgsEep3N7jm+lsYIefRZ4cLz4zFZCQQv
1reulYbW6+YAUX8ghE5Md/rQhEXK0G35ISFGfKtKDaWN7oQm69iQWBNsRw7wMzju
jxyL6r3l2CA9ndiOKsAldKJuvSIu3zUqwQSokxSN0RyFK94ZbnvDILdqOVTgzGN7
tIMLuJe2qWb/Juwf8JtsRAuPYKUKnvyks82aFmlY2pHB5qbsKO6cIdQbikeyu7V8
I705peciG7x3W2+Bhs6ftnT4vDZTZarV2ODh5HdqUtQXkDxDLN6qCgi3lQt0LwHm
Gh+PGhhoicWS8Zq2i5K1N6NP2NUeMhJRIZ1IM25Wo98QsaGCHebmLdbew6XTpq2b
s5yqbqr9FH851r5kPu8yrRZPQyDmDFoAWjiSytvZavTcnQx7Bm7Jp8HQv6iUGKzZ
Dw01utahgqaFpApYX6KkSOhgspAZrF01wS73kVXZLGCXEKmT1VVci6njk37Ewmmv
23/Bd+aRrjw3XijD/MR/89NfJzWhS65Hh8NZieNbJfGK/v24tMe3zFquvVAb240N
wceDVGo+p5FcqbdTRqttYAvHrO6ExWI+7grF+5X/0ruGwrLqYYH8HT4/02NHtu4m
bBBC4bhdR9R+yJwa2PeO94zj9pCSdDBkIezZWtNWeFlq8NyqEmzUyo3Zz3JomYTa
uFlH+gq0D5zhUib6iFP9nfBsVt5CFvzYd5ZVS4ClbB0xKkdZHZquFwb9U99PJdK9
5oDBLrwTZ9m99+740gMW9Jmbv4rjNg9yojV06PefTZUdfaxU/vac6puMR0Ln550L
mq1ANAypELWsphsl/INhbVQz2H3/H85SMvz8aJJl6ZVs6LjebYxkSzhckilBg9eZ
WCvYp40exedlQ4Ziy3QmLBVkvF9vBDdUfn8UMV2hbeDacgF2HdvdrzjxIZP/Nqny
j54Col2c2NAVWL43h01N1/3VebHngue0TY28h5vKeQvQLyu4QZ5ZocCAdLZeUUeL
X09t3P7R3JKDBoW2qeiM/HCxghWYQVFUCnf8nSGiQQKkNYZFd7bydlsI7BChYg5P
sFSBXH23/oo/dhMETEvzH/hchY6FehxgkDeaQlns6Rh+pLrdFyB2cPmOr9+XiBoF
N7uppA880UUPzO6Xif0xvJo5SLAqwh9uzUoQXBDwFzB52KAKcxR1tNdCpKYTGqHC
ln2FKMGX6avS5FILxA2M3ULNX2HLGrzxpgMvDNxCCUH/mG9zG8JmY+FUZF3PLruE
Sl4cBNlzw+ha+kcyrRzLo5aTWPBiymfBQ3EX2iicE8fmY/qpvlOxWPCvGLQIIIEd
iE4C/j/V4Hz0VJQUU6KxK9eB2CxocE5QBiQhb4gV1mXJvu921QXuxFjPPTKjWyaE
t7NIVp4u2vh3scFLME028qYS4pQfwi8KQ+uWm+9oew/YD8YU0P40zzf1N2Fy85Ny
71994yWEiVTN6hcu4rhgZOjF/qNr5Et1tKXKHO+iezd6LIJ1hoCNNtixyOZLMptB
VOrMDlv0sA+G31lrPL1yRjkuH23Pusw34MtA62joSx72vaztnko1DkDEDxqmuqf0
xuYpk3Z5+/xS/rOtwSisuzPqJ3qgVBP6lKxW8XiH1zsTi+rMJs2wPuSP1D6jctNp
3/oAU3kjJ5n7Q3z/lxlP4vZxMKJnHQBv+WLb9e69zS/S6L6NwdsiKEMM1GAxhS1/
tsnNnUJt0NMg9LiXPTh6WUU6P74asobnZX4lq7wOn2nkapedb9rvASIjB2YCdEck
zqKlXl8xqmaancmk87OWKIWrnIH3gJvPVgYQOJ9wxs6qiCgLVPJyy9Aim+a5Idah
n9Wg8N6pFQfAu3PpvkUKVjxHcX0AsuzIeI2OdXAUxDKaa2evVeXnZyqWIiH2M9qD
B/4vC0xxawmBDpknAxw3aCOGr9ulzJoX1I5JmyNCANbRXnTXd/wZZlSwBngknUKR
YLM40Bkovl5EGBQ29TmLHzmTtlokCD2LFOVIQs5YaH1Qda5jlOzVtTpuFOO5MDPn
5yd8YhzL48Kjv1iobuTGlGgEpFyQnSn12rLxccYWvm61Dn82z2pxvk3qOjPmICtT
/dM93j3xQQMQcB9Ah0W4+MyUdZ++LbMdQqChFsMS/JjI/SrxDM08fKPGUc4LL5fs
RNEUUftnhJ862eVOKK1ozf41s0MEbOJ32YiqA7IN46LLRv/To2YEuTXdVU1d8DMy
/yyE8EFYr1ZbxLTs4NMPHr6/3ex0CrR8EPy74zHr+O2omUzgUB3MdQscFLZDKJss
UMyD58dOIiN5HuqRgvgEm2Ym154uR1UFOGc5/EgTOYvDVBtkgTnTjXF1Ll/NhrMv
vVf6pNKLcf+4jXzztw+95z6UX3G31zxtofIMTH2fQTTB0MelPzlpaiNblxuHQsBa
1nD8ObAldrdEQn+aF9x0j3e0nTUaYUe2st/QKPZertV1I3PA5RUKqXcGEDIMyiGN
V/uGIHTXNZCPtg1Nj3oA//b8i80aco1CMmUUX6W9wmuAbJx2KQ4H4lyTI/+A3fn8
+ziQgEZXHaQ1cFTJmQeZGaG+XHTF1yz/u+bUzKCTEsyVlCLz50V5sQoiz62cC1ld
kI3Xmqh65/69dfNNhjhve4qcUm9h483fs+laQQWvx/mQ3DMJXde6JTWZ/7sKT9+b
VWCridMCX/oqMwdjpogePvSmab3RoPPFwzgGflROH/8GOsgmVx0olA9QkwUxBMBJ
gfRUEsP294vEBHmwXjBymrJYS7T/e1FOb3BBGN9AwbuIZBK6CMhj0xRtTBI+uvC+
srb0opYT6s6iO4hNM3vqQvSxn/AY5TIWp2W4rllQugjllcmNtQTSPNX1c3IrZ/yt
6WnLMOo1ABnfQab08oYgZd8yiPjG401btZEnRh8gWdr95pFSRzZ3EcpsZd2FUmte
q/NBF4+HUzVV8XZ8xAK28HyNLYwzpVz6xOcE5xazSW0fi96hhmPbUHc9+9oeLMiu
kRsIRuUE4IUA+KYKn5WVSnW1SvzU8EExGnuJuUYkNE7cFtryb9xBhawEkOlH2eQJ
6QemTgZgzYqLfXxF/JOH1fG6qiWb9NaI72d8Ti7ZPqVJ6bTw6mpr3nIfV9nK01Ky
VNm4HWbGp8itjoWUopzh6Hd4YHdZjDY6RGSu+fFoZbWlDuKcpxJJl+ATKL3ZlJgz
0OUN2WDmTTh4lWfermvzzpr8p5q52afET9Fcw4x3CS54no+BdHEcZAnnk93Kdotm
9bOhLYd8F6VGMLYYk1fJ4DN5/DJEccvozVpjJY6qAawGhYtAOHWGfn3n1oSsU45z
by2TURwO8Q+qahtGPJBheU2QSjyN83+EdYjip97H8xxdNEqECqbLJKwTLUorfA+t
gYNv4jTut84ZZS/R/YXlcB5weWwYq8/W18z43mzMDXIKi04gwwwjkfId/NHFaY5v
aji3K26JFsQAZ87Y2YkbMDbOponLISWLH49olalLYCW3vNFhTn1+6BCvHulRA4IX
z07FpD5tmoEWWHGNvtO39AyVDdZV/0/AEa2t9ERh22zG7p6WTMFSrnZGaI5NDwN+
0ROjjxJrE0QJsnp49UZYTO1g++yc5zkJMsKtOeq1Gp0yZbOBTOFPx8Wi5yxLk172
xUoOgr898nQExNXKlrt2Lc22Gmt4IMPCZP2JBVXCQZN2u/D7RVOitYSz/Bd5zQh3
ibzbvDIuZSr8Kq3C3dqUF+ZaaIvWcKc3s3fJ6kmWwXG6rkIowGFxCMyksLIIGz+v
QqIRb8rR+ep/ifzDyWwpYYLQQvTfeInWsFHnTzjDitNNqqLsGNil8zNcx/Da0qQy
E7BOWlHv3zFtESqVWlXPSBiwGgXYLlAwOBIct4GlngfNh30yGvXBONgjS/cT3MOC
Q35PqRKF1cxtd1yV0NV0ahAnB3nkS1/2oSfCrnvY4fY7AJ1XR02Xbwvr0Tp6mxjl
wH2u6V80c71X0elbTLP0M3w7n4lVc38pCRhv1Jq+WysDxtjH3jICvV8XtR558jdP
2GxC239oYNRa98ITjrxDcJTYTApckXOIMzUbKbmPmHdMd1uQT0PWGTkXbhvGbcUi
6fdVomx06Uy2gqVaMPZvbiLsCiFe2aVWKReLcOaqCLp31735LqcR+yR9twMC82fH
F+OJeqTmBSjilOQvD/1hQXIq5Gsse+iOXG2e1aQJY0iJdZfuDO5h0linNxy/vWqc
fB2ogPMkF4S73Bx6ZUDDQuT74ZNADDBNhoCX6loxvJSHEfF4ZUiAMETgclNoYS4z
ZC/tWF4DdS8fJxETAjshqiIg/qfbYMJIz5JX7/GmPUm9rSQUimxTUbuoSkysfsMr
WshX8l7zKR+Pv3pDAOX/V90+i1qkbr8PDf8HenCkTSYA2ijtskai9wpXSdyU3rCg
YIeFCG0vLLc+ucl1+Dc1T5kxbvVAbXnBJdK9JRLECLvDGUkmukcNvejrSCNlWTHX
pQJVksPJKv0VmkCzRdWTU1HSJMDFQvg58D92/6l6OpBDs4SjNEmS7aRLfB2PdJox
yOqGBwRcfeIIo0SxsJr6juDjO+bFwEsOuNUWWvggonDF4CMWGErFBBBoeBRdz0Xw
sr/ZXm445tQCFEpglbBV+aLC23eBD8Rti0C3SDZ+XqD3ZfOCKOGnhecQLdVDBXGt
9nBKFBP4b4RHdcxtD5TrzdfNgNiEdCTG8SBn13v87yYDwGg2bm6eIY9LLqgM77K3
VZa0LxRth6Tlk+Xiy3bBiYN/HvyM2Nak9eProtr9cDr3z87qWIL3jKYQ33yp2L+K
ZO0ZC5UHMJLxmz9E7W/m6Wxf1NjPkR0pMSTCbp+NimW8RSaYr9AXKpAZGx8xUCQP
Cy7Et+kNUIKhLeGZ4Uc9waHqY/G377Y8arDK+wCdyahjbUbg5nU0ahAFOnxKe2ts
ADEpgK78FG9bqZCy/4fF3/BUZmS7MANYZqGuIMdWmBkuvnz4wMoFx3n4BD0OXYOJ
HaklaBD0y0E1erTFbbXnPN8mvUyNL4Yj426AuCkjhU+TxTWMRLyiG0HWslxNVBSg
x7Yy+sMKBlXMm+eaIOfvq3Xb5z90XKVBmJzd72ioJ5B06o05HnBaVKWP0699V+F9
ietZ4zxo4mdFUngvm0ad1ZWciGmWdozm7JGvaTDtYBHQKOqFEVjOyKnM/g+Vc/Js
CE0QYYmz5cl6Yw4FIOHdXOrIMStNf2dHmdQahDd6XefoN/WLmNRIQrYI9DiQoTx1
Sy31djYG4R78UInYIzjy6Ibwxi3kg0i+lsA0ZBcXMEzBGXy+YSo3V9BDurTynOOQ
R88d7i48Y9bAIv3BIW0eiSL6zxHR5cx8cyXJpX6VmDDxrmqNnkKawjSj5NA0pl4l
nlT0QFdgqoIls2synY2lrpz4o0f6/sTzgSwDxbwcCx/CD5M3XI39SYYl7feRQdZ4
Qk2Vci1iL7hw5geqU3b1GMj7qonTnP/obPruWoZjh+0Kz99uJylt5McWWoCQfatY
9zCztGxGfuL5OemraaTzdCL86yzl6Yji4HcRKoNReecdje9mfEqV6ylRQMeTbQWu
CpzDteGOeGieewhIuf5TJVbPaOGpZfHZ0uZ4Ze9Rw+5kZyDw5P6NmX1R0FOCix/r
SYIhmrjfTXaWCVqC/GHC3IBOsf6x93tsVpZhx/DHubLUHE9oiCMhsvfN9WIxcKfN
sKoWpECZSikHi0fNT05wR3QEzAzQ7912nFybMNQU01uut9+s6f16QN07Qn9Rn1EQ
3R4JqDbeSnQLXV4bpwahFIAjs1WlgViAGsUA5klAixSe77Gg26xr5SWNQAn7S5/3
57ZQjEA44bNwmqtv6F724P9YlN+aZfyPXaubOZvAvK0cjO3gxKtFG+HXZRMVip0A
KjhzNBFOigGar5FHdrKUl+bm2J9o5XFGuj5WwaI6E0H1Onl9nPiN+D7T0TC792JT
6OGw0AXRQk1vseIFZ2a9kiR7oBJ2+QDP36jvmgWxBNjeMLdbks9D3PjbZA8d0a0J
K2ubb5YACQ+NGH/shQ5ZBBMrEtq4xepmGl6hgILUhg/BPrQnNyqO37Jtv4VutaLa
2tFURTihL3VMfZ0uF8cRXrpXaos7OQgmoANy1TsZsop/P/jWApoL2OTlTRBOR4s2
C9mqUdfuXOhjWqbz3GelItA6K2CeCi0+6LiHE1jv93CDZrFnyprtADY5QxC1777v
qyCxbK73t+PXiebDl5cjKhSS27WJd5rgizFbstgO/DpIQxTB8VqCG6w2zDn9bcmu
9oeLugN5hmdwW2zrLHjWAIfKLcYg6vYzlELYTOGoaGA56tMKxp5wZQGJmgosbMvP
HfK5G62IzEWzw52RU68KiP4R2PqKvYV/aly562ZU4/Sl2HaSh2/IAbcUd2uUZPiy
m726N51adIQKhd0pBO1Z8FoO35LFS/GZk31zapLgGx43pubPvm+YNDYyP0eZgRpE
qqNxOAosFPIgBFTm+O2IBww0YDV9v2xzkoeF9MSDEYy8vVuhAFWw650v0ZI/g6qd
K2Nh6y7l6Mz3eGf0tCPsFnrytWiSoJ42+XEVoLkoDLETk9/7wbBpjfb/2eu1M/DP
MKd0GD9i1mxgz4psTe+C79X2DgDMy8gqkOdsCWcBAeHZ5//ozS2wd7tuguo9Z6KK
l8Wvld9znNP9jMdDZrI5gTqPXJzgb/BOM/Q88uCdltRf9KD66bJMNVoaoIJqs1FO
Ywp4My1M4ZQheEziyoHVU0R/pksCcIHJ1+OUwodiSNCGuH8iv/Pk07QidTxNRBcz
E1jlYveq31PowYUVsO4YA4nGvXxlwkthJ4bqVpxNyZpAz0FqQnUG6AKFw2VmEe5h
C6ko4A5BXAwRLlTUmIloZ9cdq1CgvWUw2pdxxx7/+XNZQVAiTacAmX7RivPCJeey
wAZ9MPXxjDmtEAeNnF0ibuMPz/V44AWWr45A0fx/ZPfAjryZwwHQb2P+hX27k66q
EYgJcgfbj4P1hB7CZAcDXI+aS8k0YucDyBSTvGydEWWDn1XXBHgGHdd65TQuJx7P
exnHxPaThUFEHYUNGTCnFsVHQdWMUfxKSRem+jSPoRIltku1vkxcRUWNZHw8gwaZ
ITtSJSyCxSlSRNhK2Zjne499B3MHv1lr2vE/WdDiCc1vNaAXhlITQBNon1e9mfsD
CTqktUigVwe5Q8I5zToQVZlGCNnUblt8E8RzPKM6s6P0ZoDCOQWZt+AJc5/IfA+a
MDu3D1l+RYIy+ftDAm5Aw1wlfG9xHGaRUg1pKAZUOX3A0DqiUIp5hSDXRux0/pbf
5w2IouSPj33SPjzG8SmixyTqmm2bKfHnYaYiI3I50qq2Gw2ftlcEZYYHEh82Jquk
HkViiMiVeAJd2G66azq9zcAf+XM1Lj1D+qowk7weLLD8R9a9U9jCD0NILz0609AB
mKza2ptTEwg9k+5eVanVr74YSZvGeZd0dMRqIwzoIsev9i6DHH6GVm0TT+top6S+
NIxuLb77Ttj5jyepk302gh/3jXWMcqNh+1HE2YAZUM49z24+oqQF/Tz5w01x5gJT
cglt9vKlr+gh6gZX/Uxl9yxHgIZn3H57R9LduJZ1497MxedWTiTdWWXC4VIr8y1J
g557S4xlcJ8mPmvpkQ8oPujBUhzlkPHC95pRLkBe5dxBwT5g42MvKriy58o+yYqt
uCxIa0ebUW9LzRYNjm6hERLRmNzqfDSkcfkHuldv4xja0DB9Yc+y6t50jYwqCmsy
VAoRUardI0l8/EY4juvujKAqa7XW6qdWbyU2BxK5Oc3NrAVnpgxeX6G0CX5+/b1m
heHRb2H96VV0T27W9jFi03dYyFeW1Ggc9BJGZEX4RXr4x7QwhDZwbEuDk/F2wsF4
FFZ48YLDTJTXPIzV+eXqmHE35Dkac0kNivBcgU9Qu1FUKsgwlzmt3prLxSwiuHNS
zTaHg10ebeXTLSL0a3DLCjgxray3gFufIRYjTK1GS8z67xjL4IeYZZCeAYEIMrG1
MI3Vv3RFH97+KF5BW2YLdjX5CYmq5JEYxz2TFa5WDN37hlu0gzfqV3fUE9szJYxE
2z9CEUfsqH1fyXhYbu+BOwTvetRXDwXmtGr/rrBlStepUYYcDMSxO8E9cC6MaMXN
g25NNBfzI8qjFRuCrBDWLWEosMBAaHg6CR/GDzI7WnGQtY+q5Eehn9Kf0fLhBWJ1
sdbL9lsK9iEE1SjDcvoJFTMQwGRX9v++NKG5sc/84pB5HLYvHBz25n7t08ICSKIs
cmhw92vdwkd5W9C6DUTpRWaQaHp6OQPHu2xaKdOXWHNpkZ+c2tl4m+7LXc4jL3I4
P326WtTjcAA1sToE4Y6JpIJgoB6/cXS/4BXUQMpjFP1LEd3h0PFqK190Hipsrjeo
bsrebyuQY5Jv8ZYPZTTuzL404svCiDc0vI70qi/pMuYHIt2oIS4uevPCgKJs2GZk
P+ThTd5I+mJ9grmXdFRCuy+tyk9eR9tE80ExsD1W1zA8HZQaXsDR7j5irvXaZfZ3
P+rdxxdyR+MBaK5PidCgWN8u837vUUTqqUPljt3sFkBNimFcpR1aKM7cDdQbIYlI
EXg8kr46+OX51VS9FFz/JeCR7zX8gw4n7XU0YirC9SU7wmcR0XTbW5/5kMO7RZd5
QmhMRXs/2ZqwpjCAhM7fzcZFrOb+QU93XnoV7clqwgYrCXWYMFiZoKU1xuv3+Edl
q09/8YNNS80EonodRJdROJLxJy1EUcA1HwGyeqVIngMT8Sygj2870WXY+1IeFe6X
/hOUurB/oB/mBx2ktJ4Jv+s6OUft3QFNlvuX3Ib/tbK509KBF8VeXnNIU6R65g0W
68r3avwRX7Xa+cWRQ4XE4zJbicbD9IBZZg74wyuEoLc0Sphjb5qU0CDAyzjpiLVu
wUR67WozAF6r8d7neLFMJJ94j5b9vUChZjmMAs9vBRnXVZiwsA9dGGz9pbuO1M83
Ob9wq81rXuQMlxd4/xdfmjSGE0eyQjVrO215/HcPqfZMP7kNqaxBySiPXMO3rfef
kxB1faXjJM7/9yYYEuv/zYBvF249nYlfN/rRe84OK3UZDcsZPKgfn8TqRSwVYhCL
fY/Txd50ZLbGwPdVkTUhdfJpqeRTZbI/tOLve4ciiQNEuoToYgKgygiM0ioSSB+7
ibQbQQYZQ4crcVsrXYnwuQSgMfODcuH6l+zbw8BehKq3QN3M7esVMp7VhreCcBE8
1v5YVFQOyuW+WBSeHvR69jMi9bA6ZPqnYQ0P4o67ZV8ThFu9TUyzLivlKQrlD/J/
wzDnBbYDsW7+G+MQKtbH6kLsdE+Gkmiqrvj9jgNLWFSd+xJLa775W7s5NKbpRJXX
pzUXqiRv3CMD6eqITBRuTOHZA44HgXCWY79kmjNWJDSAqmY4U6/zniwUYzPVvkUe
91DsEbNTj25CAzyCCdAwKZYZr8WnfDJR3Ip8/V8RPn7wtEBBU768m3L2J9j+yILG
mSo8cFMgkzzuHaW5Yii2vVmZ1I7/ntU6UZ3XtEdpsFz3WGUGKwf+U51zzxNA+Y5g
8h5rKKLpLJxZiPP61l5/oA4BD4xH9mmx0mqh59gCS8BSb4ddTxIpjU4qOXXPJyak
X6fDryUT2Vcu5uy53opG1RCMnuLuDkNfWZO2I5NaVrP5hrKtgFVdkubGvQf16rkZ
Kcv9qH2uAOPwxn2J1AVKpsWMisep3Nt4IsmIsLo5MFcrEIAOA1aOguryqK+bigtq
Tu8RPr79XyqHmECjzzfzt8P9GObTttx/quEwrxwBiF3yyVDiSzIPYMSQ6EtAIKPA
sJBntHzyREKvNU+PzgTFSg+e2VXAfI+RHlGmy0doV0rVZd1rTJRapKeE/+IL7eMg
aa6L34GQOLKyT4mNr955L03yghYNIB04UTkV0/cBcJAK85d2KIfspHWONqfXR3Vd
me4nv+1a7eT3iAy1ggi+kiBnO4DhvvrKUEjlb6feyJpiLwB8UzZIZvyXYdOKI5c2
c/rn810hJhUECMqbJFga81v5xvoRd3YkyC/wrrdrlpBuirAjDVx9BjsIYR69Ifta
kpAIJa+nGFqQk5PAFmlKlbbtlFHgX3NCndcFSH2ZWPPO4P8hvg9IS6LJsMw7rmfZ
NNOD2LzJ9AKV93MHsG5cRB+6uikWhEL5KUjfJ15YFIS1b6SCpY9yTI1xuBZEzHdq
7BO93BofQhnBoDxWeB+rNktCpQE8k6eIbtS9z8U3fyS124iG/UXCNAfZb8wdfdhL
qfpjKH4Oqm9UO+T1NBTQ1u/FtftPVA3ZMRZ/+d3y29f+7MRvksLjHyWkITudnQKN
9zmNtT/arVf49ThKcr9aJs+UKdxtO8MV8/jGi2Url/qdHLKCj8riyQJycSfYCcxx
ZqRpDS0eu0lylw4VVdewZ/d2yMaAsf1EUBYmIXUk+l3wHkaQDRetEWjZ/QWYVbFE
g0Vrc5mlkzK96qsCmXq1ugkV/B3KTuXdzrzwGAc4GPz4NgLYBuCMvsENDvEwBDV0
lrWZXXk7xUdpXxwo7qaS3lcuux4VePZOizuD6qf3yI4l3K8L1+dM0j2HS+KZoNUk
Nlbk1AmJWgCENMcEdW1idzVcFc6ybXCwbky5sqGR7g8e5k4yW+yrkbg6YNujMewB
wtb3isEHL1jdmhO13nDxMqo7PfwZHbjcFBxHXcYANIa7gbwysXSn8FcISd5jnFPj
FaFg+bV9Z0w4gb6sUp2gg1nfKbMCBaSHjZo0WzQK9aKIeLHPksklzYzoOqIVNL/F
U70wwg6Qpu3D4F9DJUNT8vK9sxOsSXKrcI81i44pyxHlkWfqKgeBMpzD+4+RuDVi
LxDV2HIXwFFjjQt7TAWmvQlgefanj9CjZHOOEEBg+pfI7R+8ByAtQdPVYuDMQ80r
kaVAICqH+K41vdXksc7DVNp66pl1idKqrKPc8dWwyx35Y5FR7SFmyoO4QUeSSU8i
y2GGZi6c0aNrh67uxyVR1Ju4ro/7k99jLBfprxL6q3zEdbcktXaeL8iBV0+WlbtP
BXlVaNQC5agnldvqnwprfiETBHdqiuiOXgOz3dP5PharMOm3tiz0yw5zurn2Lp2S
GHHRZajPBG0copwhuQFWXKL5XXIl8NzPl+ceZzBYlwQuygAmaRxxeA3iy2rmJyx4
TbOpovhxRfv+1eHGr5d3JkajiG5E52YlW4i7J9Qr9C66491S3YfnpqlmVMzMA8ao
bLJCGq8yq2oKbNjUvAZwtiyoCoXgatW9/S8JGLEdgnx39XBwyW1cguX20LesZ299
yoCHKcf5VctqhNyV147OngnryJ5YjTlkN0xsogfmqEXwQxYJWvklQkY7Bx1LLwJL
LxN5uQveCVlT89PpGjUqayS7kRdb+XdTeCLLNBY16TdnilmkiVd2jlFJLXxC+MQC
KIrrucSdM3SbGAVSkIXhrN5YxwrdJ5dN81d32A4CWv5xYYcYwOK0XQ3uJUBEtWZ8
yVJ+p+U1VU71hsHeDsxuFSVgV5wJogE8aRQIr4I6yCY3/BbinWpz0TelGQEQNkJ8
HVsLGbvzzdHDNRn8YNSPJDEJSycMoaKCSpbmucZcBN9LJ47v8HJlDVqDamZuvjSs
pZHxXweRXYdDqR1bf04Ay0ebqXyGFEbRAB/UgZ10cJWbBpP0UNZPRsLCNMdEFOPl
RCef0wpc+1q7mjyDjMoMZC94qcRhRyIc9F+yo6BBiu+uZ5W2wLywI+gv78kt8ZZX
8HlUoCMzL9EN7cR4SXFyC4L8CpT7h2KTXHVPrWr+OCGY7/udPvEqc0lGLbPDs4e8
DTo53X+sLDa4J/f6AU057WR7jjmhkBEvz66i8dbA104o/afSx28V7GLDUSfNRWJR
p8rMZpatV/9xibk9voUXS25iBbNpz2vhbOo5fvbi4dP2MLb0mDYBa8Kynr41urwf
4RDNaeVIoNy0491cT4TGx5ZTax10QpG1cX7yTOKugawlsRtyZhMjw9CpDMUIKXEX
ukI/LD2kaW3XR1K/qF1+CisZShgM8OHis/rutzecyqH7TnWaiZvE+hgQRFXc5z2v
Oi/T8a2V6Zp1+gr/lI0V9j12Wsbqtyy2K7NJnXh9xvdxW4yCJUjsev19ya0ZIqW2
g9jD1sfky/SYbH3opH42MIeFUTUHnOmS8nNRzfvvrxuaZdlzfZDrKQxM0G7ollgA
F4R+SI7F1GFMRyaAEv8o2fgVhkjDTLYSx38DkzorGYhcJnoMzpR2rW2royNOmCKw
6woP1ig8q5gTHYxt16B0sYcNLpeO9EbaNmYlozXssGVTOTAE1vdAC6NsnKu4Koi8
5cUivJNMz8Nhfaiaw5TnOyvPA+DGuWjSjH2Yq8Qsk4R3+JNY6HvyOJfBBej5rOHb
WxdO0Pj1bwyCuuuoP/1i9gI3cshf9nLYgZNnj5nDzQZ6xzYXHUqRbxPXCFt9toUD
ZtvfcZdwcdkqwFW5+HJ9sFuAbrqlugSyobP6jbZ/QCwf1jUnazectqhGp4NAGNQM
TrdwnxttfxJ8WIz4VmlL2y2JGXOwSPUOkJ1GKa4HnA8cpP5TglX/yA/hCYM9GODG
VkmJ9FIkA+4g02j/I7ZcIppvSa09s9zSYWjnBNgJUMXCVTCmY+1GKZLp8LkvqMPc
w60hbOZIYUF9TnEamPn/WXDEVrNMuqpGavh2iSpQ/g4MbN2hxbPYAk9FU8AAVxtc
eH96LtUMlleLrf4ndyhea22bAsNUnt5zDCviHOM0p7xoB+YRg/jrCYAuR8GRIlHR
En7g0CWLV52dXteWDnooRXUWgX/2gGXu2dy/pNfBws8+lFaH63wjkr8bYvGkJ54I
/qzI+tOaoBgK3aqO8am1qbKMfZLhR+R2aJlLwPa+mfkc98GCK5ZNyq7//mCY1hNx
M5hHbvBpvM21zDIf84723+SnsZ5dBJw1Fgyt2MpHhVduoB9NGbojoxMvgS/+e68E
g4T5HxnSDYbrcvw+CtaNRTkj6we8G3EJSBfSh+DH46kJ6JBoo8mBjHuRbD3dSEVO
FBZ38PwTacIGOOwW9BTssHyLpJRO4R7CjtemGAl+vS+Hh6xn4ve5iE/dIXy4aeP2
vb3OGvK+dfFNRC9AcPZr83ucZ/v430ALLLN3uvR+P+hzuC4lpFqg+/n9DTYsWR76
5aTwF1j9tf93wTM9cq37tmVmZnqG2sqwLMigLyrt3r/Met7Xn+c3TqEnhrIRAKus
XZ7fE0YGzBzXH5k3xAv7pjcvNXNhhRHlnfrgqw0195DWsb5JDrADuMWebR9HA7KB
2IU26n/QgfSm6yx1fPgMCdV6jjMVykjSwfMTGWwVAOmghsVH4vAEHOV2nye2fByw
tJDqbXYKy4l4IpESe2N0r5ASlVRBPyE+bPkNw45mXZAtgu0DLDWfsQ2lAZlqVzdb
scLNpKV7M9BN9fj2AVUphPF5dTTh09+PQZwJ+NE9vPc4ZxD+OBjlLZOsgXbJx8xT
kUOxrvcW63pM07jZQJdh6rKn80vYy6kTaH5mpCk1NABqgzkjANtvpGqbPcF0tdBM
RNa7wbBAkSUMw9WnjBvvUCDbENY9cIy1qJ8+sjspOpOc4n9rOzSiC1hmhPjiv4pM
xImawUCfdE7AeJHk/TPMBG34g3vAOT2vRagPjGyWntBRUsPK8qLcXZiD8X3Cz7d8
4fKSM3bDsJvvXBTYw41D6q6TtV065pVTtfiXX2skVlZTedd7Tdxi+kSx8Cvu2lll
2eydidql3un8kYnBQsv18AEdba/sbtyCNxnMwarqSUtVnXKymUGzpKTH10MyNG2G
Ya/yNeFj6v9gc4sFFhjwbSaHTltY8AwMfXXPopLT8HHMWqQiGVfINbVyP+tGh7I0
V1EzIyWMehO0OaX56IGFKpUlUAcrVCHk1+AYQmdTML6yIhhTGwi5+GBTLGRkmLkT
EP1hef5p6hbrCJODWwtJHGd3M9Vcn9lcZ2CG9IfGvGYrBLQ0L1glJUNMHFHAC0W+
Vp00tcXi1+szQn09I9Ns4H0MIlMrvBSd3eL7Mnai0XuYACANAfZE4t9slNuc7Cju
RRkMMjimrRnQfY6j5hE/nfMTi/RG75mof0+OXqIqy1huaPje2utv8tvyD+s/Yzhf
5i4VY4syFIFnNOhcHgrPfsf1P1E48Lt5EYLxS98E7jPid9vW92rVvI1terRFY0sa
DfKtJfXIuXYK8qkJqYFQVklpH3hzJE8p8ks41JeQPMERPL2UJZJ1b6UYb3tuAOa4
hF3fza2t3POD/MxxKDeiPndpovxuk0Y+xg4XSRjvgUqWPYTBwVNcamaIYFrb7B97
B51e1uTUiV+it+guLLcpQszLQK/YEfxX1ZZkM1iDPv5yF/RL7FXz+M6qNONyjUpF
5WOY3i6L/XrZgivyXM7SQeI1S3E/ENZnJQAYHuhFFcBkBy9mxsWCV3MU12kf2wW8
4J1JlVsx4BENN2IyOivk35NZ4VEcS+jdLQju0kosIw/duWlpZccI2JWGTAHBBxe0
albK8gQtyH2Qu4A6Ra47HxE2GWKSCtS9cltvRx8V3jCaqcJEsF6EGMIgYjOfWDF4
KOSbh3seiJW9zAlZOsGxB9HxRyjGx5csWv+G+wl+OEUShwp0OqSUK4H3FlP94p7o
6fuGzYHlL3/EDe+TiG/oR614OItuToxNjiFXYeKOJFWLk7c3IIGHiBUPG1PhcJ2O
9FKKuEEX53+dCfuL8w7tJRBJN8UwJoWXUvnuADnlmSTGWCuTIMGRBOFA7YKGM+0g
CDNEeaPpjHJE/6HkaesiW35dfauqkuflZs6UbMHLKndyDMRaNZ5A1poUUcn1i6vp
7xBa+Nu+RK1OjY2ZG21oDxjRK+get2PYy4PZchyWRhuALA0Ac2+oZvrra8r8IJiM
0IBT3pYCEsFHxS84fi94ZC9XKD6+hKTeT1qI8BlQHGNB+l1SX0s0TbQQVRlAknld
lJr6WkcB/Av34zqbfk3rqvctYT4NrsQxLLNNof/mjw3poPgVkDk0y9rARuwBuEOQ
8AhSB9C2PbeLh9Kh8e2x+evxorV5stu97cwD+SB/iVGxMC9tAkux3+Sa98Eorl9h
3cIqOy5nMMzcaoca27NV2dJv3Byk4CmPZmWw0SasmWT5r6kk1v1WeaG3qw0d49E1
Cfdrsqj3pEQwg3Jb5k4syDI0Xruvd96fHR/AjBxyMw0wbWfvFPPTpyODVau18q3C
/8+rHTjDpIia355nEXzXXqV7Gs9KzDCD9cfkeQ1X01V342tVEU4nQgOgY15hBFAh
XKfAK42Ksa+WtXbLuln2egWT8BpawamtP7BopEw1ixE5gqK0WBj7hCHFqQoLpx5K
N5ZvwJHi6Lq0jyURNQ9qkPD8RvUDzHwAyuhIHyr37/5d5ZG5ii91v+3IadFT+jt3
KWjuwjjLnIiKZXKWhezvtWsfBYK1ZK7loODkVLmdYl3RDkoYnuWn++7nQKhCCzCt
1pQ3ldNpQEk4fIYTaPPtAHffhlDOJQoa5ESMWxo99lJ4exME1HDXUnEO0nvxm96W
o5YfE2wZdPaFvVqqieUVDNvLshG7sBr03g1R+KrofKl0gAbfx8377d5pMEGTD6+a
SSAM6o+CTzQeocbqBGx5UJt6rmy/aE9pBIbUFdY4sk6Kq0RpHL/eBQOoPD0dCUYu
oJzVpE02adNHGZaeMQ2HWDmYPiYy9MNmLWyZlvnnYOYOh+vt7d3ozLEVchZQ9DNF
X+Qt4jnwStVLKCihZaQ7BQiAVBg8wZZRcqcKHkQYDnaoKGUhHoD67C86iIMZx49G
2kgd9KhKLrqQSEQNnRVc48iKMcmbbUqV+kIEoe3xV9Wz1I+yo4Yim5S6O8KKPIxx
sxzpg5/yVhzf7xcNAg5bxaQBS8FD82KmujrSCyzydvHHLMt+FoBWYHWeyTL/G9x0
yFoI7MX7wB/xm4KR/OHbOPdp9My++pEu4fD+ejMgUbSwz3WL0uiyzbdmX2tL6o8L
yZvNdhDepB0KjFerwt0Eb+QvXmBq59dI//XGEovWxMX1DXXjSmRyy6Hu+rlKEurl
bFogcQg7fpmyXEpq+ekADr89MXVHBtlhGFkjZj7dB9Omy9Nl1Tr/9ngdHLLj6ktX
Uc9lff2djErvZquYSVTEn85WrWW1X0EAJWw2DRe0vpQswaeyc57d1dnRq8KraSFG
pftcyu+fjooky/7mQ0O28OSocvfPBN8NgNni4+1DWUxFUx88x35W2UVmhZJMmxmC
VLkUkxyET6tsdQ+D7Mllf6u3rurG2VXYXmWHKnyIeYkGJW3pHk0FsWQ5NrJK6bD0
u40RjzZ0aqcjV/qrZzpgeq7F0X8d+eNf5bsjSBfOhBkqhfJhnxfmy2AKGpiPu8rq
ahJtZvv1jt5jYdZHEyU2iRrcW7pjYjXHjT9ysh+scwa5Jcqv9W+vYup/UGeasCxV
joS/Si0YgO8b188OMGjjHybkJ2d1XrXGAR2CkRBJeAvzlKes5Nu/l0xRCx6Xdxgt
COUbh9Tj0jXYg6eeIyIdcGN9pE91sdMWwn/dsbAycDbTo7NrFNyKpXNIUtuVKyGW
tSTCMq0A/sNF9pWhNMWtayEIuDgOKpxMlzCnZvntEOj+MALlNZdVBw38K4xvWDaN
/Vbtqv5NBEr6E78f59EwziqHQgk/zd0rVnau2uKAXx0Fe2N1fJpcNdSD0j5iREHd
nV7I7h76uDoIHVzS/TFU3+cqHJI/bMRHBNLhbtt0GC72S38Heg5VOIwhvDx5CEM4
EBDx1nUdTcs3Y4zoC5TdqihL47gpuoKVzy44epePcWS2Bhe5F5R8sRdURZUljqgw
cQHeObe+VKAQQU+fPAaC2T3XC9OCXvgpqNmbYiAlnkpLNlCBQd/JPYf11SjSBT0i
t1ZYIchMJ307Z3L+SE83XZ6zOvhARyEXaCuv9j4wXul2ZP25Xlk8vvFi6G6teSkg
C9iUkczxGOJ/tG3jwxoUb78bd6hF0gp2L7GQsdsBtAYOF0c1fZL7Bkxgc3RkI9bf
+GPPjlrK8oBoN5yFWSU6ZAZkJiLxjzvoWLdCEhnjteJKdQNIlqR6g6J864R2msN0
0HjWFOA1M9mTN0ZENXszQlXN7LXPwW/ZdW5JTjTIwCRWN6prI0kloPDjDjhVz2vm
IhhYLove7ZM9JklK5G/w2OwsbYQywYj5/EzxpBPCRR/17p85p4F5tvlIlkqChDUO
gDM0l02SBj1RoOYbmv9ht8PWsIvAH0dMIb1n738pPiyXsN2DfMPMJZDP/1AeYH+S
q7Mr6wHp407m6eKr+hUFMkPi3iBh6Q9FdL68zBCFhmJ35UfyVwj4W4g7EG0bwEZd
xuGAIzCte2MhfDgeI3Djk7JS6+kKLOY+Ww0CUIbKS/Ecy+Op6d0PKdlYbKt/vjbW
nkS4B/f+6ZUnVi80SA+aFYDjzJdyC/hP4l0aP2RALMRjeFY7bUgoZF6ymPyzUYsp
L5d79LW65VoBDP3zJOziv7/FG5alQVADhDf7NolepsX2L3zYRCx3pva5TtNaCPyn
BNSyW35OMS+vwkyiLUCAfPIf6VOVHobl44Zi7em8W0T6k7f/n0ycbBoKn4x9fsCS
hEXoH0VlwTgdDBIZHVKHlAoOltVa6BjZKeBIEodR4Deyg8YGgxlvDYwZsvchQ2Ij
FmAHBGshVnKmHsoFBDvNRJYGi5uzKi9JJgV6s7F0JFLMXXyXS+T5w3AAtb4eY9Yf
W638PoJHK8O43WtWt8ghUloGlZinS0sn0dOVre38DVDYJEH39/W89WO8+kki06U4
7FDKmyLe9ys7NwVc7PciONlqF5aFFN8SdZQhXSvvgE6taUCdmJ87dOoAwhiknIuc
JG8boLEPvup+hgZpnWIMEkkjsDer4bo/N5reeMQC09bTpeMrRMHEMCTS6vd0b6/5
aeXoBdMJXbU9+ynlsxm2uua8PX56ML8TzmJBVfdqf4rWYvQMz6xePFX3qSncQvzg
iBcTvy+bKpqQpFteu+qESgVoHORtxKjN9kBrgXKIYoZQkHtyOWWg6i/d4OiqtQNQ
ITvvc/OICBnYQ8h6xkfDf4M/fBsoGPeu3gXT6UxJvRKhEdRnK3qKlZ/LnoCeRtPI
AU/O0S7xyaRoH+pogdqc2FnpSd1BSEAbAWFtqKYINPpRbduGuQ3U1XhyDGo3vv5c
9GbU0p7UvXFPBKk+4Z4uGAyDXbbwmmHqe/WAg25aLSBez4LuJaztQASd4+5hUtfO
rMdVUa6rWBTEnXB5zNcHm252rU/bPJ0kuX8eEiOYmYTd/RjC+feLtP3Tqnh/DuTZ
geI/HxNPU1RwbY0qI42ttpt1oNoOFSRcMrM+1JMt5bnj1IbVrHYLOb0dH6jt8af1
fAvqg69qzn2/r7i/quQ6O6w/4xEV1xHD3l1XjtT3JguQ/ptr2V3IkA2F8D/9srZb
Rl5IR+kqY5LeijtrbJ3SHB/3CRhP1+fSQHfH8KdOevjNjUyC7oIUIriwpeHQsOWs
r8S4a7Z6jNkT4v49+cRSSvIJCA1M1kiQZprFczwfsVssEOkuCV1jm9MJvobaoNim
zFovv5sW1YdwfNUm2nOexPT5Vbh3yX3F7PxNVZSecGDicq1dvmxw4gbdczu7TRWV
xVPabCLL4HWK7kWKd26ezqNgqAQLHuf4n1lKoAirPXcwVOTq9Z1SewkuLTtWxg4n
hYN4san9mqzd9S6IBQT1mzKziTjUQxsFzCbY2ONebSgBWQaTO1q41pod1bn48z6E
O0SXxVqu4ADf85dPV4vxLXDQCkC590+u/OPcoLQ/io6ldwLVav5RDaxBjEFU5xui
caIuM4d7zGDWeSJAcKTs79ustj0ZWh7pq1BxlOACC7oR1tRcbrVq82tLEylJIlKT
HSJBwv4JD1XSDq6LyWPqsFhmQrpRnIo7eXolhQJ4mr7Fjo7KMHe+hhqEbAY5ZURE
GjWwXSO+b2Ix7JSckU2epQUR/3vwhOexck5htP2t/zqUnbQk8fm8pgUfB1FeB0MR
cZe5OMS+Jb3IBMprl5MECNLGLWXfFcWZzTvHLUHR5NdmBR7Lw14SP3HWOOpAbCOy
GwPWN57GsRL/0hRf1AFcvnaFCbhiJRPR+usz32YJHvy0Usmz8EllogSPkNSmPrAZ
e19ny11pEkt3tet7iFJ3y8AhP4g19+tASLJ/VqFidyno14W7u2gm+EkD+3n6GGhq
N8vBuCbQzTHQ+FploVX9IED5uW4x6yQPNyh86oeSUP0DT3drydssm3Ki3P7xD3nd
vnMyFY9/Hhn4XY5enMrIVEQq2jEDqMs8J0lTEmmqoH4D2QAnLSXMYzRHnPcgfsOq
ovqh12sN8X/Us/n6hv0ANK25OtkgerME2dyfClv4YD9+2faWJlgSPYwdmT62kuwE
s3P+1qKG528k7u64JtQyF0H2umXZkJfIBTGJCbTH8rZ8FRQm4S6rerN6kKk/8V4g
fT71sfwBkQ8H4/h5hjMxculIx+JsfscgzhMPYlywkD99kUVCUtQiStFlMBoQwld4
LikhcUkCbAMEaNF0jM/UqIPWC7a/zyDOLzYexZHOvD9ksbQ+8TwbkJtKE6g0ao2A
wK6zsLnFZqSNxBjagy0sOlPADy1GCrM353fu6XUQWdAypaf760EqrjCdVioyq+IW
JeWXUnlkfSMeCiYM8HdsAbutG8hXJPfugOeX77CM88+SdFVZv4IrzAcrEPYjO6q2
tALXKS5D1BlkoQgXrRj5NkY2PQUKSi3LU2A5UEj0OVLNaYVzSq9iKXuyGqJ7GQ8C
/HNrOwCEEc13uoRtPEHoPHJChN7PO6dT3xajrO6HQxH4xRqm4InIdZT/cGlDflOT
Trvc81gxcmyovzLZ9dsd5n9PoJHsfaI7CYVuzRwLj9A1Ky6ZS/sKXwdKDuyAf091
MDVDS/BVS+qmVox1ONp7uGQw3XAUM/P3iccj4WpkbPJYykYWbd6ZAJB44WU9XQFU
XBvwEAL4qcGcoLAcHR61ilXwWxOhRYDTTf4iAOX8sPB/Typa5lEzrNK+dR3vDVmQ
bxO4nyPdPWchwwqxPE410bzmPG4oKt+2Ez0AQpoqiTURff8xwu9eZWb8h+souXh0
sta4jM8ist+vlkRdKqObdU+V/nntxBfYCCZ0rUXOTtIQ2H283XRbXPGTHs3SI7zB
W2l/NPqlhBCSwxGLr/KdbRJs2dD0LD9aKjM0h88cEtjItb7poLYLMw8y1z7Jk4z/
+/hAKf7XpBR++ZwVnHFfbCZakgpWfgXCnX/fAijOrnilTX1qS98HcBtFGO5Ojb0w
XH2w/IwiNlusmdz+zVLJW/GatVLLWzjBScb33H2Mk1ocsGm8ZKqFgeis7EgJUPAk
acWQDMmVpst4lDKYjHtPJIqLtEanqzbMe9ChVWVHKQTwxasYZ5CQW3RJ/Ht6Y4Mk
if3fXBuDPuKp9mDUlQw9ilvnGsQQsFRyZrlPb2BYF0WztQhBfvk6P3T0j8aKhYmB
mX4riMtOVmBBsccUOI2DfohAPGO7LvUSNI4z/5E5Xc2v3axUVBpxq4tpjiJ4PRnn
NuP3tfmkOt4wxSW21M6X7ji1hmnnh95uZp+MrPa15OqbsxT6SDuWch0b20AkgbA3
D0flRD9/+DUjRFkn5xorcSbcW+mFPTjN0V63FpU94hTVDSnah+IOZGSvuIG3PXIe
WcxQOG8N8woNFegGS71Y8PJnxRMz7E9YHwj5zdyd6TDGmsjFzXsRUxSj8IG4+Lw4
rA7tXzhsmGqSM+kl6iLV7AU4IqIllthVyW4DcQXJHeApb3QvX4tSVYSlx4LCmSpW
a2c6cdQuAFDLtgYAiU266Y0kXo44+ebIyYj3PoDbIIEZVaVn5awvVgNAtTd//sGG
0VAslVsS/fMAgGIZsYV55+665+AjnYcyNDywchHVE2fzikvaB+84HlIRKJ57tsPK
hgUqutx8yHEIgP9osVjxCttdS18qURMPQwYBXtlQojyUKoxyf+A3RIBkdvypZ5dl
3uWUXuYF7jNIYA/yU0AeGqG+i7sqkjktATONlqjfMWI5bpPs6gqtvhDQprYhY6/e
ERNP73JTZnj4IoHFgqlp4k8VPrkPOOIAziiKn0DCtvEziamkaqEbrTpp/v6TB+FX
TpE7mKQsvieTBkIG8k6R3HgLV0f/TLwEcRU6ggavGj4N6Ra1dwBxyWgK67C/APEq
iX8gr49X9UDn8cKHMUhcCRgsmd0KXnHF8uYbSwRkqsI1Dsh1pcytCZkkafO9jWCh
EQicg3vhz4N85uQuAQSQPDlG62ZB8Rkml4czU0/AcQPbAQTnYuWR/845OLHAz9Wu
AXWhHTXk6/Ub7TQUImL3P7UBTyBfIbITy+EmBtzkApif03x+svde5dkbkVZeKgAL
kS5yyvdYzCibk6eZTgkWyOSvM+hGZ0sOXTWFSOzsGqDXsKhcaXpYD1MwRe8fbEWb
k7FxVBc0VtAkGjrtmUet+mnFe1mjuGuD50Sd/CiY+XmPW3k8t/kNFiSde39JuWOS
j04lJqWhqYyTTLL95BNWul3rzjh2ySET4eZu6WsVSrdKtmVuqJsHLUUvw4AE54U/
MuCg02c3W+hq5VD4zkoRSh5PTnEOBmHSbYPMwVAjkB0cSvRvNvJUgY+NucPSVBrJ
0s8MUIGlloDrvD9ZKLpeQRQoNisrGd8zOkpN/RZVwfu1Lx4czf2ByQ7WIU6CRhbF
DdBVSuwzuNtLKqpmJMXZhWCQK3gz26VZHnATVGUJj5uEdXHs4hXANW08ZihXjsld
lJzNzlPbH/w6YcnPaCPeUPtaoRU3qHaI58h2m7SNe7QWcvok9+S7eik80pigicAw
IKHlJVcNOPO2tJ5j6wWnhC44jX+hMCnm6tcotuTMdcd/AD23WAWEE1PAEy7iLUvh
RAi/gigi6S7LQYxyQLMYuVJovpskeES44IjSp6b7ygGMtrvrXZRdqGOvKw9wL+4L
NNits1c/dMVmJkNrkcTRKxNXxW9fB17Pb40BzI7QoPevI/2lxxBsKmPz3nS2G2vH
LFashjknUWtPYAL5bB/AJFL/c0RjaFG04aVf52lZw4epFQuCxIxAMpbcUvpXXem9
kCOmOjIVk5vK2vG3zqd1m/gUPaBCo4wx2ITfz6UdPzbUgHQX97vdzdam5zxGUMhp
bgHujKSn018pyYAAs00CQnNR592/cBDr0Pl1ZzEUTFDM0HVa2GgqCAOl9QHxIKdX
pXCUgojlcRxlO8U9p1B1nUG0Lk99mivhp7usIpdyh8TFggC5wkcthro+eFt5Gh8W
08OAXomTHsB8/B3v7DyROCEWS2xBeR7rRZb3BbcHgjkkSlJ7J1CXd34LEu5y+cIQ
aYpkJWkG7UhfMIkwvJqpwb0XoJfHedPBYg+3OZK0uml9I+aT5MkuGaFKEvuEDKG+
blUukX4aARlEUtfmKJKGLK9OfdfNyVulU88E2v1fcY/kpJ0ztGcBS94aVdByCNYr
0uHy4Bf6AH8oBzI9hVjwbU/Qg2O0SMGuP0A6H5W6OJfWn2/cjoyQyz20HJpC/pwN
FzE7nDL+kCkIU3yYGEHMH8BEmX2s9mZxYzIH9L/Xz9+7d2jBewKm6nMmzO76P/L4
BO+2220dkKzTAmOX26ylXU5TmG9eu/XFnzBaNW+LS3EpiAUc1gRSPgY0VykHRiW8
PzL3ux6BYHwwX10VHS0EHh1srgGBmKJSHh27ZHuQQDQ4qQ5af+dHqyet1RjFOFyl
cthubvF4RP9xPuCg0A0INNecbx7KU+JJFfQJHbcADThZDCad4PIAvT9FVYdVPD2t
w2IcP7b2iKeNGYiu/W8dlO/6DsDlrqYJWqD+Rzv4DnIDfFuafOvDHcpFHS7Mcvfr
4WEm2hwOQLecgMGqY+NxOlCTDdCO7uYN8/hx0cjps62houM7q4B3S0yREs8FVAaa
VVNjKi4TFZ5X4ag7mBVm20izooxc2S9SKdj+2dU/6Gb4CMN3+pIIipmzjpwH9tHk
lQdJ0eJx6r3ZhKB2gG+W4p/JsSHM+XpeG7QZ/UUiaXqgxQXJSRuuJAXkVpvEuhdG
B+xYYg0IsC3RBvLGe5p3oqeNlEsYfE/MrhwTtlR8CVlXOHFoupUycP5LopNqsZbi
ToIyDb8ECCJXnJnZnWW70Oq9NXuHFAnQehiEsiJ7+vHzvsESnQ7ixzdrG5Cm3g2e
77kOug0ckVgC0P0mQA4ZyABcDNzlnzjcQuTQ+qLvVhNkFg4z1XBnIyDPr9xo2EJH
DWlgnebH5QmxX+QihrDErlZKzr0QG0AOLuMCAYN8jFk0QTtZPDY/WrzyWuFqiuYl
bAHrzBWycSO2KPPMDktoi02C4ElS8uLiJ/iODb2XDxdkOfiaoaRqfYyfYiVNLhRu
8hFzmzDANZekqBbf7h/zwCPHkdvZ6j59pLDwpfzN8yn7NydRV4JOnZU9Ol4t1rRP
jJwM1uVO7BhjOhmYVVQVKLoB5NIW1GAlzRdZSVqNtKjKeOYVfiZ+bQvf5H47t1hz
K9OIlNYm1v0mp0oBuFBFMDNikTHyn761+9axfCOZbVtazCDnbSsFC92W421A9BSg
Qsp2UfVz/7GP5iu3PlQm+lIOV3bQuVqQX8UHtGB8678Fd3YzdmRwvKwdxg4rOazU
fBgfzidru4a3iWoyFPBXOQDJRzCgNhAgnpGS+SZlH+zYje7lyxgo6joYvQR89+/i
ofjXmgY5ZnEF79omUSt7jwsAWCDI/4VzqX97vOFKjxFWB41g4x8DVwhvlBJTfwY5
o/rvao6vQFR70yWqX9BDchOD+bvRX8gA2SI/BzzrSJfJT1eHoMzkO95WyMEdkQk4
otVZ5LXCbZzGz3G/1hpPnQglqBeCGv1NQEykAhapAGBOfnVS24uOQ3u6Hc/rT6Ze
54IBn4x+fHla+qO9XJMgOZJT3vHObl63thUD1CHbonT0HmkoLj4fyjTQZL/wqffy
kNJoCGIIlKNF8UeS+PuqR64i3J6JooY4FSvurmZGxBPfVC3sl8ye6rUBXwShEw37
Kf57DmVvs/OU1rhMDpX7CcbLnU1rcyg9v4cmIm6pZWgab9RRedAWU7dBJ3e3vHCd
0Yme3+XyJlIr+XjYtQEzEhlXBz5KNmALcC1vEDyPVfZtPNCnv3sQ7/k0ghdwis6k
L/4HCF4JxFP+qvIku1jVD1J1qllkQ9BoQzBrCw6n/4Q6Ey2ZfqROLh5D9NzTCEL9
1lf3ZCIeQhQRLSkPIlHxOgz+VL5ddsQnOYfJze235GfqKF51M+KdydtwYB7/wcBE
txQIYoZ1J3M76ZRToC5/rf6/c46Y6vOtRl9UzXulIR0KanhUXsQhOM+vRSUDlSmw
XsxT5acDiX1zt3yLTUSPudlYlw4Wy3Xz/YxfH9lJSzwZTMiPXoIBd4hhImnST71W
uTqkrVTTHsUnl2HGVaAcK7Ywr/xlNUFJHg99AEVZDecRQmmPJUGP68xwLQQhF/3g
x6BIH1zi7hgd5TQEZ2+ZEsgMEOGNx2363veIC83AIcwPg2IR68u9haFtFbfsMxA9
3q3RC5xZTCtLCpQdN17fLutIsFVG3I56e8yRKKARRiU4hxAMG6oV0YHkhZrHJnic
aVUxaSMsAw04aZNJ9voPJ0riblFSC7iumoEUzsBEV5rdPHuikEEupTeT8XbUK+Ha
8g0A8qlgBB3F3RD894CcT+NbClhnsqZf1kMKh0b4F0woAj065qCBe9flWa19XcIz
Q0no6JuMQB3MPws99UqdYocY8fhm4KHp5FNCFvDoeHB+TuPT8fGkGQCIPgGudu9I
401SLLtzTuNyQOywIuEflcng4Js/iWtr7QnHASuRjQd84UTyGGzGQo8r5tm9CGYa
cNbxOQFRBEVQiJ3befVxvwYr9xVSlVes1TclX+e5K6qR4AhP6AJ8vW92/DxrIwit
7rsSiNHgAB5I2bc3gkjNRqd2z+bbe/uYtVszO1AMopoWUcEtBHOkJFGQvfvsfYX1
auAh3SFLO9cQk2oB94z0qXtfNiWKYpVW7ylPQoEWiSq5O3DgCwF/pnxs/WzWwyK2
DAUEjV5TnE4TUHLL/ewtPFqkgeVXy20TYNp85cuWjHplxRFad7zjoyxTKHTa4cEN
O+aPQy2bewtRHr9yOjya7+vxqiYOwLdkXQEHSDaPHr7Qp5VVynhuUaRdsHttTTCM
TC5d3PWdsQDjsVdIoK3C8WdyCZiSiaHlvGoHDvqfnLRXgbh3m6mGVVHS6SA9C7+6
87ZHYgQ6Xm77J8dUGoQVJXThWeFLhUwh11Bc9Huhta84YUH41jWj273YKtpBfKfn
g5i1+YnL3ooWNVaJ73rh1hvz/8+M+rTtFOr4Zmtq/fvq6CcuzUqtNCXiScnO1eyG
Xz3McERaes7L5jKvzedcSv2HmVXJA00QKtOFn87Bolca727McWwhDWKtQuMDUrf4
dMTp2+QPaH7na5SGTbVxr2iC1OV5u2us5sx+4leX7riRkegqNv3D/DADoP5mzCke
u/1lxW6u9MtJO9wJScoaw0uCSskJRPY23MmZw5Qh3Aorwt5ASVbqZ08I1o+/4niG
T7wACs0qFvR5QMJbBBaz4tzj2P8Ji+W7hDgMgg4/bazsso3ecaLU4A4hWXkNjQ3G
S47RZTzvbkq0ax8OlxEEyCXt1QRCHsc5pPLMZhE32f9QbpSOdf7lntNzYReOyFrH
w5ZcexMLkMzy/2YhbX86E2OG0eA4gc1aDu9AJbVVIGR67iE0mpbVEGIuq3fkT4hp
epScR+m2AzT4JMbQ7biprfTGAieskcea4UTluBtjmdyGGyQ7Ijf+owkmqhPvhGlP
0ZYr7JN/23cBiCL9OKXp7nbC8AgmOMcJqcuqchxBOaQd1LZ0NGUpVtqGRbfsLgbY
Ssp/QxAlfcWg2D/HOY7Zi4nd/beJf3W6KOU0GZ/+H9rgM0R3s2CA38fsiHnzFFbh
hsfAxJr3cfqhE29/uuUb/w3M8V2H7a0do2ezG2W8JoOSpclE7Xz9d7q/y0G9UuIp
DxfUR7n9kdxFWEHo4WHyhBqLw9LoaliCO0LJTx0jaCKm3pNrPReO9x93hlv9GHaC
ddb0k3lscHs242qQmYNOkjR63XW4WmMCD5PLfXSCMIsC0Ei6eggD3zXBYrYvkFvK
YCp5vdo3a2UXL3Uwi78fmb+qQtowAiWPhGeGmG5yDhxZ0QL1V4Iot2dIKTT6oWek
kv3mwGaz0ZtufZq2Ma+24b/SZx2lzdPEq+lHsaorKebZvxSQxBbTH1TzRIDW7gDd
FpEsOciSXAjCTf9/n1+kUOV22uVLR2OFQwJDTfPJiGKYwykmHQtjzciXbvTGkcyq
27uFCoHju4rCOlQMJA518GI6dWN9YJQJ1bOeprrtXrJr4vsx70a73kvDQZH4EuXY
8fkB6X0VDZE9w6NZ//URR2x5VntOjL4u+6fx3lpnrThFnTppve3M8aHjTqyJSgv6
V7Hh0Zag3PnE/Aa7/nPH+tswWINXX4lhZ+RRzYcBwqEGkxVXo3/3B2mVZ/WAKMzp
SfgKI8V5dvcIN4PPno88OrZMzqASYUFWDR6amTAfKrdGW71g7eESkyfsPPFu/vKF
LGLFOPCZb77yU7bmu9ed9e6Wbv6GdWVlklxvDD0sCCcGbC4ARXGPlFQuhToAANaS
xLNX+RXMMTimLqJ4Vvg5wmH1fVNhVWKhHpMG3lOCf0yfcd/2E2dEK+B5ovh/0spf
xrUIbAJtObhzxQnEhw/B9uKuCeYZxHxLtWkhrpLi/pZW8hZWSmuXYE/n/E2uzgUV
XAymFWfHp0mU/C1i0kNIH75H0jVNU0BaqmXjNOdEeOOBR8UQDB5AfldnYwsrBlL+
8i8zLazuQSRy32slIBdAoyPqp72Nn0YHAWFoAAI/p5uF8nvmoD7DggvAxtl0ZWtd
BCSCTUPsMpCFLGKEA3Z3FcQKU9vCadiH/bow03aMrN2pSb2XhNd8KcmOyAqMAZjB
3tp4RfqpHrJHLJfMnUbTZhEL/7uDYl4rKVQtEXG94bBACtjWoLS1rOcVWsKBRMV7
KVGIYQ6ErnHNGq2b4f+/FWM6m/CRjDouWnWTtUMi1wAvlpD4s/zV1I85UXp8OxZ4
fgmGsQi/AC5iwWjFmmdG/lkZb41oc815wQJmsziZvYQ31flDO2FR+QgZKJlT5xzh
CY872PCFSFPyuNDzGbTUyYe4vEzCioaPSHDe0nBqWbxEOOA52lu4hu0uAS1CrgTF
dnEhOPSYxyvhiUUi/ADCKYfHW4Rsx5R9Vwv+a10VbgrMEtd5C2wJfu29Cm4HBlL1
0VT2+wr79xbZ13iFJ5nHvVeG7wrr3/2AMbRzANiY0j9Fp0Bm/2iAfbi4U02FUlB7
dEDbjPQe0zbHXgVm+0RmcuVvu6iwsLDurbFMBk05oRJLx9i8CgriDSXXfitEgiFe
KBegLzV4TTJ/b9rYToNSkexMOSV8tAiZHMQgj7X2gnPwXhR86gGWNgswflXFJMrX
6EJEnOGMm62IHWiLD19OaVHsA5OuNWnVCSaVtI8XpPIJWl+o2BBk/PcPvfGSTydo
XfTWeXTojHI1lwPIUr1ZlM9jGOdvOd3XB6Xf0d7uOs/RsNX4sQ2oTR2MnnwZSl4K
jyuQuzyuDQ+1OO081PLhGQZuK+enfNplRBcg+JysHEdWrD1SceXcHWS2pu5Kqyfj
vLwF8cAKtYVJYS5RxyvFadgcA+7QXVfKQo5fa0X8TaBVpkxjaWVpYQaT9x48U64I
WE9p6xTIMmxhNgsZvTasXe5iMYPZyktl3q5Z1OPglnJFemKWYvdKp4FAs5EOlMy7
VCOTNZQQIfrKTXm57EsIuTs9W6gVxa1l952OFsLYh+yShEzDg/wRAbUxkbBTzllO
qlUqMX6dNc4hQ8TjjVPPEI/i5d54+VYyiCjCTphTrVVetDbmkIaOAusxDX0RugPA
xG6aKpGoVZMG0WUQtRqtJzDUw39vu/v6TM9V7gKrbIkVgxgP8GCxPwinegZ23/du
x61IDfSq4ymiWJy/h7Vokw6XOTCnoedS2kwVWRJ6st0lYtEggoNDWho3WnIJefUk
qyM1h52sHMiZUXZUCRzho3/gm1j7U02+7afYdW3AVyyV/gOTI268vViYF7MUu8o/
gf7/uOol4mcUExHaf0LHwBO+JFNtZXkgWKvko3v/FX8Bi5AxA19rx+Y7BXkOZc24
iaWHtmNhj+GBWR6eVIIbqWkVFtT8uDP46Z4I7V4eKSD9qkMZ773fF35Ra82yqmGh
84lQ1qfZiumxAqmPtSnugq2DtPZFuk4RarBfnbpi+UD2R3XsDIuzQ3sPpRQEIslf
jyHeuN1Q06fjXcMF9m0Tb87F+GxrL4Q2s6RtDFSmUc+/TEqk0NxRXiqjH09pvdDg
hbsOanEDlUw+lK38W7G9BLTFFpHMEj2OoxSCyj2IZyHrzLQi05wMpVEj9H0LYnd0
61UN8DCcKuu4w1VR27LjA5/WRksQl7K4+wz4iuEsnGYnntn8yfJCfFwVdQBvIBom
+XKcFO8tZSPqM8LSrcUip7IkcFCpZFGgoz/1YvP3ljiq1MdnbEMtDrdBVidR/LwY
JFkz5gqaO9dHMo8QDSsNukkNlWzv2xciiTBUYrgyyBcRebTdhtV19HlibCS7g3ca
nrCkidJDZmn9JZaFrWyAFwmiNwCKoZDegG3IengNNtC1ao+6unPCocfsk3FjK4FI
Flyr2qa8O5PeJYA59IzPpH/YCqBZKnx0AfQYs98tYwr4GH8SXPRpwoFXHm/YFWem
W0bwkvw5zrx26BMQhmc673Z/2sjWHQ1Kh473zMpg3hRZKLXNTV/lBDhcIc16u3tj
9UgP1FhlfKejOglRc1tHxnFJnv0iJUc5qVGrVMX0bNcEzLoI+QDcnoskTiXoyGd3
1foj+qZMmfRhQcBAZvLCc5EiEh4vEFbruAwP7zOaj7s4a8GggyNmwUy/3+X2/w4b
B68Kv3mzNk7j3SNXbiQ0a6Ul0KeA5QAzcQ2viWcJ3kb6BeXEsNMywD+/MIdgLmHF
WsqBrZrHtpgp8+DpVVUAD0rFSGrSNk4Q/3ONdu6YQaCgEPSuT6wiZVlB2QjYV56F
mnj1jmKb6KlT1thhS4b0faIvm//whQpU4xGs83R3ZUck8W2zfPxS7ESkU4obu74W
xsTzHfRSYH+Zl1sF6MevUBK5ZzRSWyXKklwLvWcSI/NzX4B8Q7MJE2AXZHFI7uHl
xpNnQQWYCfY6oZSCgBt3N//WPktThj6wyRI7CQEGgznBOJe3yPpO1KO44Mb/9wzS
5FBJPYQgNoLkB636W6mltOQlshYQj30cGy/8dOLWdbkQs2cg26i6DkpsZG1D1NV+
Lpd9z6JCrF2MN8pG885zdkY98v3sa3ye0Sonarymzvyk9ShV4NgTsbosV3BfyiY0
SQZK7qdXpyjqUlw01oI2SQL0q8h9RjzgKS4gFxd+QBR+zxSQ71agaFO4PfEyna6O
y6Y7h+rArVmehvAW4cQJpgPmxdGnf/kAXlwM3BmUchv8ezc+7kPE5T0NiGGDpW7x
oCoffoW6IaNMD57lQLkzLAzdYpmV88Cbewc/imhhHgUVuxrdYZ0PcYLwVRanJeDf
alLm7sJtG2JQBO5L4xQ6G6PfadK/t/Tm5x9s1xWzumdlVRnuAN52ZvuXYYQTfjYi
n8CiWILbPc6VEjfRYdUYwP98GjENyrrkxhKfX6rmPh9/guupBp1w+3zV7AOuhxW3
iE7AyvNtHPdEMr30CKqXVgCeYCJU5cNBIYHo+YS+8PPxVvVzARXPUne1oZ2065X8
DIReVPgsrKh6qhCI5aImYwzPj3W64t6sB+DAdgpO/yiYmk1sPtLYqFC74Fxdnrc8
utbdi6YNx8cGB9Xx3VsrrpJo32CJpe5qbsysRMl+/xjFOTsnWL3cI/zGaCyBF4Fi
vq8WDbABgwGRz8iMfHKu1r9+CH+bBpG6vKRaiXkdS9v/uTtDHdxavOXaL+iArBnn
+6u+YAox6hZXFdq7QOSxfX93rEXhy5ast0opRrfx2H+6pWK5VvKTH9O8WfmoHGlE
XD2o70L7q16oXXZKgjKgtmduG5+boPnnohxrpPj3Aojbml3wrgkXyQeUrkHCcjAN
3YhcSFWDQtBOcqie6fCQBlUASLfq582tK3QatOGA1Sne5sIvXV/YI3Z83xTE5yAL
7BqT0I9unpMLgzhw9WRXIqP/pGjcr4cjV4INX/uCPGbACVw9H4N6NwwQtf8g4+4x
JiK28jOZsc8ebfHmvdFFNTAbAB9gG0xsOizQQVLxKztpypKTqOw/mbf4gQM1r72v
HJrZ6pbbiiAGOQI2o/+HRviuV1fM2ZOatIHJNGK2bplDyxv5bHAXqirNbUXIU43d
nYc2Edp85FY1gWfEFbkG1igi2apt6DU7VALbRZVU/hwVNIVbs/cwMoS8lnTs2RbN
X7Jq2KQGIKwMc50/41hHKOSWeh2RuFLlDScbbjBWXUchq5VTAUdqfP0Co+nPUheN
SYpCPiKP/6y/juCJqPPKdPJpO4S6URK9wRSkCHUdyJdBbba+EpwreLdX41qumbSd
JS6lr/s7Nsox07gTKtEeL+LHxoq+VCwD/e1GgoUNRL9ojdTAnso+OueCZHBK4BSX
PYrSBvEU3k5TeOZ6j0nJTpeL8tMHmXF0MY2yLMJPKS6Im4Wto2wc0f0JvHZcdmrt
JBntITavM5o2r97IgSoM5yFQEWghF83juU9Z8tSKEPKIFoCcB+rtl/k20lZnB3HJ
IvKAQSfyjoXj5YoWHSu65yp3B1x1ci/3J3Nqwsd5AYLejXyJiPYyAWOR9b7N7bYI
PBAl7Vtkhayri1dT8lWF1F8MiTjW3gpY5ofcmpNTcyXktmxyqt6GmXfUCmY/e9Pa
+t7LM31hfgKYZyniOhCtNSIVimJcTZtqTE277QndBRNuUmaZRO/7t1ExuCv3iu9H
Wn7jYztSC7+VBIsOcfpNYzB3p/E3hgPRlOBG0A/on52dnaxYGCTGeb30xWhsqym5
1gLkN5l9GDtFkEt9hMtlbgdh03mJtUA12WMgBd74QpJAOXZojHaADlglsNpY7rB6
VZxsBDuu684Y/XQuciuyBtP4h8xvjQ2t4IJRGxvS9ACojBTTWhqYT0qAdZxYrcCm
HE2Tq40TUifpPMHzdvmQTmElwzMtllYQQN59hLOWuyUdeHv6GLtmxF+KCjXxVc8S
e6v0Drw8BE5dMK7fLaKkLEKB6TskXH4GmzErN9P3LmQ6yRzc3dk0K9PrhnURrbmd
auO8/MM8EmfTlYHpG0U2iR9ApKGiaWF0MMHMX5acD7uEBTk9/S+0YiE0CbGdAdWW
k60cTiK99lXrJVjzfffQ3cn4lKy3LUeC2l3RLFmM1QGQsAGOdouhW63WN+HxZ+J0
znzlh5YAtDWG9zG5yk+Kx4KZQb6n2r57dwMYq3VLg6GxufQo9Jj4nFSsScLLWy3B
noMnVKXPE2f1oGwirJe0/KEtGXsCSFi2vAc1XdFkzUVonNURcR7T8T86N9+NAiWF
msakV/gJpU9evDplSioFtFHnZNkc05qMfOT2gBwf+0deKrmoTEXA1rutuaaDXcoW
7XLZhrB2U6lKcdGSvvZlitAAQiRyEnkuQwJNVsVCiGKdF5S0Gk5LYUmo4uyxPyIu
fsaiPrrrk06ZPrR8H0d/kLYQAVRqc2eSLBU9sLKcgJj37L7zKBIRXizBON4lLHrx
fpADKG8WXCsfGME8s1dcWB4uy8iKveyheZ2ZpPjcGh+xriOjSkMWGaZn9aWmnqMn
AWisU8SjcQWBMXZs6WQthci3IcS3MRhZ2FUwfR4PcpX7Sqo0eEZdrq8sj8HhZLgf
AXGrshwTGoboBnO0HWqAjPoEfZOsg634xooj/nkC7sSjL2/4PU38QG9mLFsMVW21
v1ZhHfStUh8xdOAcR6Gx3848aLYAn7fyaTbp6F4QIMuQinGyw1Mi/kUwIysLfN1/
gD4KXIKyIS2ZDGQhAzH3mA++zgy7wH+VKnFE2Z7mfdUiGBn5aLPQFrVFxwTO79Ld
0RUtV7EhM9LKsRUVF1z2w0ljq8rgFlndVsjYNpuKJ55980M25lM7Pe891UUEkudB
hC+yCmJnOKiWOZExbx520H8oqBMFrL/S5UIjoce0uWOorqpe/zEPsVygNK0teJ5d
tK2sJkg1pYGp3l63myNTC5Gws5fJkUBxdvFw5YXe2H1jng9x/0HSxvtJnfrz4A7V
8NJz8PjjiZsnwaEyFnAamhAOH3RojjIz3pcAiykEsuJ2nWOtWq4+G/yq2uYUILk8
JZUsRzJMJ5vJm1El4yFcgYEDTf/ohPuiF5e6GCnDGt6f2J+Eq7OPfmMeGoUuJXEl
5IXMFctosQWyey92rv7Gr4p7ZlnFLJuyprgpQOFRgA1X+H/eJiLPh2orxJc/PuZh
SiXKUDWmqSZgxAEwRwpyHQqg/1GE+bGTs7+ITjiYPzNZf9n9nzCy/337jOOno41g
lRfimcyif6BIhQiUxvm8IqteNyEXsVJAPGzfePL9BTeaN7nroqXZvuoDsYTrxiFq
G9R+wc1WH1lXZZaBrP1ElwaB9x6CNFqgQkx8Dtpt8/G4X7NaslxngETltD0CgIv1
asb3IXlJnTkCAiFkS7iFUSxUnkVmnVEiplZK2aD7c/ORHdSAeyNEyTFITxJ/vLSR
Wl2racR5gJnPXuQQSKKAQkb4ERPE3AD4H844Mqjlc7EJwePuUGqXKVfdg1PT40yL
YKodzao6IVkiA9waNDI/LdryJo6c/uWO+cCXwGnBqUgBi87RHB5ghaQTbd6mHjZ7
ySa6LUU/3tjdjzvO8klFsBMsJXGRQ5k3vRlNbTTVUuzReldEbpqsY16Ck3undSPZ
fmGvQgb+BxOUj2atKKVyAjQADg5V/QDUumukOtPjQovAFH/PeN9poLUFDg6rbgpn
0GcaARqo43APTFjYsUKHGxvxMfZQcZOZZyoDbgCZe3L5butCfHJpgz21CN1idOYq
Jw3vuqOHTkDt+46Ho2XT3fky8tdHpNUQyQFCN/bBLBrJ9rL0yrhu1Ix5ig31o53f
XBSr+DyAAM0LY8VyzQUnBx4ZTy7POHzrIyVaYiNw0/wvts5pPDXpJr58JTu1BfrT
60MAFTcMAZle6qTJsX/6N/oRnzCb86ZlE1FJy4X40XUITKe44+w2+4kCXcgA4Xqr
LGR+spoNET2Kiai41dwas5jUco5hCJfAvCHljW96scqNjVt5V/kejGkwG+6bQsKo
Spx7rFLCrv94TRYDE+uMFaEQ2/l72hX3Eb5QK56UUD4QRFjvJnNVy7Qtxm4aLlxG
nFjTkdZ/RrOIEh8RJPdJZzgb1s+PQcnbPWtXOEIw2o4RYRNUk4JgKuDxkFYTPHFi
WawEdOq5CJnD03r+m/UzkdmkH6TgG0B0nddHowerMEqzozebXvLbKvsKpiRa+33D
EkY77HnwhZlE2XkHcrfF+yy2QDiq1Sl3SkvaQqrW2IfM9XpACnK2mHcUjdGtu8n9
YW0Z/AIf9CiUSvEsqa4LY4/RnycW14cO/ECg7ETgDscK7jimuO7ZETsWFU1COOpA
SrCcSFgo4SAoinz0ITjFJK7URp/zPm1P4pyDyf2jtmcgIccSadBwXW5snCTB3fw+
onS3IYRJqP+3qeTTf60gkjSA50XCX79oTGCsJ7/24hDF4bOwnreSUREQizrSGYsy
pbP6Umv1YCEQDc9QjvfPoWCNnauhOooS5XjuMJdLoXplngac1nLBfu6e4+biWt4n
vMiMgnvElc+1S3SLEZ0PIN75BAx7KVyAiLyldyrAkecQBMKbeBZ8wV85KAaYYM3T
w+ZknJRi5ges4/CJK/s7O+xlg3DnJUgytzVMVq2ZZYqNrbrPHye9nAvoDu98oGLm
c9IbM3LN4aHncS4i2YqcZqnYssmGlJQquVtc6G9jBJ0ejd/7BkZPjn7E5g4RRmWZ
zs7H/B3zBy5v8ddw1BVAWirvrnnoMz8rDKei0eWKQfTMUO1qP4wQN7TWzArWUw+m
jSlx1knK5Hle1XWwgcPN3zSiGH3TH14G/xiC9D+nOWGh23OTaYUYmpty60o1ZV+X
c4SecYAFWMlShLGEE/lGk3+3el7CkF9Gzr2nJT6o6EU3Hanv4seAOcz9ymxI49cA
rvOne89a2V9F0H0ZTYkFxTdB7AybjsmDjp+FlXb1UnN9QIjIAqOTcsXcn0fJKo07
3iIPqArMl08GZCF2qDTej8ZdfqOe1iRPIXDV9HCbOC3gb65WU83yagTPDzpg9Bjw
AdBsgbpZJZmZ4KgMplB7Db5XqjskMvjNag9VoALavmx4CeUQWaE7/FJOsHDtvzBg
ZMMxq183QRbFPl84ZhchUDt7TnqhC/K6iDz7WCiaIg/akV3PXLxfr8fHGTG0xsDb
CohHMVZQiEzGNn51ke9HwtzdKwUdpzgkoZemvHuZ1rphIK/adeW1WqirTMxG+UM6
cl5KhSaa2imB3uu33mpDUPdVT953YlccVqMiWRfV3qsvm+Uo28wivXfqhtiZIUvL
mQ4ercqS8QtCLDBiLMUHn7kQcMNL7UZl9XGl3g8lhiJ+uugDwFRldB+X+EH84QxC
mFwniI394XxPSi2b0umtzE6vmQUY8dlUqU9FLwDphtQuYrlZ1NoHbr1xHM13QWmD
8Bx4SOpKDkCKDeVJLTrCJ0Lq5mSUmka8ON+gqATk2c5iC5dqzplR69raB7riKuwU
xWAe9/3pUKHaCIMHWS/DTRp9L7e98DFp4eJZNDgzfn0lhjqRR7tFbFseIWNOOPFA
OAI3AIqSAVkg+CVAngYBva4UVy78XJghUfw62oSjqNpZAguaJGAYEw4KZVk1EfU7
+krVQYxOAakwcX2bKc4cT02FH40JXh7YOgV1VFvVlDca8NHcQirdBFzo+Vgs+PqC
WXZe8iVleuZrEdWSuQqERRqhOzs3Pk+H+viFQnW2NIWhE5Er6Ly1QI0wJBT41ZGs
V8yUv4MWcTQiGVOtu9gXp13krvZcDnuZOKeLpezjsFatYalTa35anWV8QGCxm8Lq
dJKORlmDho8JVegG/IHd3fV1866igxKQqYZISnr8aRtyxop9Lmvhpdergbb0jQ3B
Tx0acjMcXePhNml+3o/+Q0E44oUPZIYeWkJPNfFDHhPDYlg3pdUmWJ0YvPAUUw/W
d7OJehBhGClrtyTcwhMb9uFdKthgiHBrBu50Sv2+FPPwRUFaWnH93EHqr9/6hGxd
ZKDUrdZ/Bi+lbiqNguzX5EGNJfiGAmV4uc6SCmIrqKKM7o41HugIMLPibmzPdFs7
K3uq/akghpuuiWSh6kDe/apjB4v5/TOypMgJoDBRVMzelBSPHUUGFkXy1Ug4lmRK
LUSsQgo/ZQ36hKk3WJ3SEtk/7WGUX3czNB+Dd7EA4hB+bpABeAswH7B0wCYyLnGp
G/Pmgn+JrcwhRIXUGUe4XneNVp2bJ12HAJXY7E5n4HllKR0SRFtR8krOsjMuI+xx
IDFZou8Aie+GmoX/iPE+MbrSbRxbmkk1L1ySAS7mDxiJ1p0bOSVvsn2POX7hT8gd
5RUw2wDvsA55/QSiyEgoG+8EjdQ7NEDg2TblFBzBeJrotbYPdzk8IC5pJOHrX/vi
WaVLZeXy7qDphYBZgCNaKb43fkvWmikqPUkNcmC0q66yLIizP7dMG+0dAyw0hVUM
55Vta64IDQ7SVGp1tnB9mlg0If0WpYHvi+kDMhttmM6gOAREbsnaa710LO5hbHpA
6Ea3hlLgQAynfo7RQ6ki8WAJ2k5hwFFu4E3ciAUqwi4V6keQp67E7bND8z0xvxzx
JL5DRJJcKmUvClnv8XlgGwp24zJm12qIK0JuL2fNBw9OdddO+jrlph12bnWyp4Ya
/MIlmoOVvglWhgK1nXwgJLWUXpQ1IwSLjqAAiL4w1+uiP8GdBcFJQ8twbs5i102b
c8gyS1+ZbD6wyjnx5CVd57K1NdVmEoS6JYDMohiglXVlfKGNIdei5Pn1Ovvsz5YL
s64UW6m6VCY6rUG6CKOSckn+bwHuS4oEaP51ZaZ5IMzXt4bAFvOg/jx8B3/5AU6J
4e8hLfUzRkf8KRIrtTnErArueVzu/gWtK+V1PaBdjz91WVZr6iVY6KddG2hUgLpg
Nox0oLirTTW+G9SNQtvmCurymZOJWm7UQiLAyviu3AELJhcM7LF4rZme956ym0P8
XtVmi+Yf8RRf6YyyIpi3LReNwjer1OI1lyHn7a26Ln70fqGoQkqZ2kTQ6vkxXdPi
a8siVhtg1rpbY/uaCs2jljGrWpEx7fY9XxZOJRSlll8sg/6fOI9Ji979FL83rIu2
z8fv2cWq1Yv9Qsouravws067o2ZH5oiFKSM7kVJ3nCNGkgG0+wIehpOBor4kiZz+
j1umxLFadsNE1oBqNNwPZQp5jQcfGQv36YUlum9Y6d8ORzLAW/DRaZ8PpfVfjRwH
1yg0KiTnuOhIuvBqs57F/OeBs4h/XAoo0hfWaPbcmBBBNXpuRNsRSbTDwP4yYrYY
mMjev4fO6LdJIXeUnBKF9qqCdO24N8kV0CfZqc1z/59xYERz82yRwicXL3ekeMeJ
hagFnaJi/J17M0GxmJF12q9a+cYe6cKxOFoFu6A63KR6HdrxSUQwMAcHOwaWLh8W
Gt2Qgmq2E6iXGn5LGLG/ViTXqhfrzow5afeidK7e/9T+60Gp4USwB4M5vcLcv47p
f/lxm6yvWsII8DZ7p+pys/nQAqkiDoqphpicr/vCu55ZjRFBnvLg+3HPVIHpfkfq
G203etkLlZ4dzg18afXs/h8pH1XpyoVl466WbD8Tf9/5mOC3/H1BcvtWsjcaG9xS
qrvX4GsIIQiSFfCS6pQxIX4zmvG8ihycn8TkwdCoz0aH/ijusHFttOHHTCp2ggLs
InclhwFIuJGm+XfAW5NJJOLi9SAidv//YK3jauyIxXFr5SBrPvXah6wzGNnyFcvt
SYP6N7Vm+b7Ja9Oe4O6JqA/IJeARdpccF1725maLidJjAC8ouKmBAOJYHKm03OJh
fYRvOpDn3o62dFdp+LMhc3MgNZ4xFDzdDP4HrO5bFEkbco+n+cfc/YjGOWvVHov2
fk5oL0tjsICxiHcLs8yrWm2ZnjmTfOyXV2wDOxgHqJiSc5zMTFwPDjzWRDfqtb1u
eSL+cdN4k2yWPUohnIHGLeacIg4osPYvzl+rHAMfRe4HJxZZ8mpjsPAkI8vFVRFA
9MQ39b+Lp4A1CSXSMaZVWu3eMLHicXGZk+gxnRtVdHnJBk3DZwNDjjoz9Uf32MZw
UgfxnB7QbI+PnN87LYGcXENlqfBWFo8lcce2law9KoXIQEl2teBVuvdTuKTCStJC
kuS1FyN27cPjY9RjPE8CeKdsJ2Z41L8Tw44jWDTSXLTUqQc1HihxW431uQiSr7+C
XREe/dJtEJA+Gfe/4MfaX+h4mbxYgUurEvAGUFlaSn5921+5/kIVaIRaIXaOuo/6
Z/ZLiqVrQV158zJ0ua7k/zOBurFTe7CBt4oTSmk4ZQWfr5cLgWXVlRhk165hVmeR
FAYZqEiF/dphrB6IinRpFkJ+Ot4x0pA19EK1kbJ9iEG9Hbq88v+kxZMEUt8KDL1O
Zww72zNcvf3JuAfSryoLPSHD3ZAYUzUwXd3UkQ5LUQTUYWWIYYMmbn3NpnjjfDHS
3aSh6fHfOexBrHLIhKUl9MCnkRkQyEqwzDiWvJu0X1LDpC2sbfGaPWohuk/cJIP+
zYgRXZqHHrwKxcBX3fQJ6/rRB1QItVd4fmRUEzWH5V4K7difRQzMlMd3qkTDEvtP
mU3eEFCzItaxZvZf83NDK4RVvWjGNRTiGsxM8+ROGZxPiJZalEz34sUnP+u2aHOd
3BdiL3crvrEFqpQPtRzbm1T4p6jk/Uvc3Q6OancjK8ub/h7j2KjvXsWMT0uYRl9k
MZg037WKSmMskvFO+d28dYYAyyV/VYb/J9sHuPH9Sr1FYXDigKO3VkP9ZgkUO+cL
FUbbShRpvufqmMPCJ2iIFih7GcOCA3hOwsbsGvpRsw36LxFYgiRU2WfOq4BxFAJ7
ieUAT6QRTN2OCxOg835/o9DMX6qojWcjWOFB8PogWl3nxs7VziPALiB8+Ctb9kYr
YO4yFytf0Y4zSrn81PwqD57j7GgP8c5XL+yo3t12CyvEQ5HQmPdGYx4Qcm2gjciO
F8RNhYZtZHOmZWDJaPJtlDT9lvYIA/DY23XZHuQPEedcOyhrFpxZxdBDZClTUpSh
+2zfF0YHnu2s/z/OpBtKr6XtiWyFPNhGbQVibeyPppEMILAE+hL7po+OyfPva2bE
4nCVDZlL2WpqteO7+FYljgboazS5okDlaSPJXbD5wVk/JCoGR6zVnarddJ2xcwjl
Z4u0bG+iKgGrlX2dkQsgMKVlGS9CesJ0oSlIu7Jdl6t/+oy7y8C9ElhK5ac3xWbj
CEKQ8e2A7YsWEXJahlDAuWwbBqwLenoHK923AR0SBbdUo/FaHfSDAGVEC5hPp/d7
4WgYyddyeZQBO4DtJ7WcMBRuft1bkx4QecWzY06rhQaX43cX1QeA7loN1OUEJ3EH
6qFNWKY3fZjwZoKowCIjihZG520WvCN7+yB9TPysDdwit/iMtdQlZ2Bi4VJI8BMg
HsqtvidY885y6uNQudKSqJQ2HsWP++FRbMxpj93cD2Q1X3c9YcwBiG8pfcudltJ1
86LrtrYux1JDCCmuI5xbI/aycDf0soTe/uNmRcEdGuUbIFDD8LvEkFxsQ2SGFDx/
Wp5k1XzAsOKBCPf2hLT9WJeJCLm/EJKSio7/NT3dqvYtLZEeRyqqYf9/qvS9itfY
bS2hMZYG7/oYk5Ojkl1auHzjrL+GXSjq47WDMId7I2yhTNEnGW5i8YBBX0vlzOoZ
7V/BG7bq/ZNI2CslLBMaq2XKE4dyewrmUpc01dnp1+4HasD92rhlI1HeNiQo9WHJ
5KW+zSmd7MWoeD3BT7IOIGB6zwyIhQbGiLAwqTkn7OvfJIgO+055x2l20HEnkyV6
qIu5ZbxgCUDV4ARq7Kzpn/UEhf7oef6d3Q3TIJPdYI8+cEaqzWmpqt/OC0smzlfJ
Y01FYmpR9QKXvLo37otUtmkxdLEC1a2hiSN8XV+YbD9dtI40ZOu4BHkRKMWLNH17
Houvt0Q9IVh+qqZqFbzwS9wsd+sPsbhgNQn1v9kE5KGuV3yKfBgP2n5Y9KX9Pww9
GvfTwNvrQmO5XPqyFi5M7GIH+voUvQ/Z07Pz6mbzRBiSsvyZUjpiq1yjshN1R2mW
EMv0/8nkVS9E28vpx+hmDXaSpsu+z8BsajRLkAqL2uR+hwIVhjp82S6s0B37OkQ8
Q5kL35gslQEOc+lU7K9HxLeot2NCNU9J4U1HyCMbJUuNH4yJnLcIT0a45Pt3ZCeQ
qZGpm3R9iSD6CUEIB47j+PMnx8SexTM4uUN0YgjstXXx8XHd8EkYYk9AhuO3S4ZN
tKqVHcq42XlprOOvOyWUFTPfv/rBnly2vRwHcnvWGNxkqSFaX3/CJ2z/jQTTxO1S
RsGvUDwUolRlvntF2/XKR5TWNMhADH2ff9+upAeuOcyIT0Np9hTtPh7e6P/Fc6R+
15DAg+mluS4XJW7b13a/QX0jhPnVCxPu6ublgld2pHcISguF6YvOC7LUcuknPi7w
8JGnh8yQzlZWRbM6LMw2bYVMySKQVq2Kt4OLlW7262ymRFcBEVNKmwQVAG0K5j6R
rVLkQi76He4E3xXxYiTXnyIodxMirZeoQ2op4kOUwFzkG4hHrmsESfef4Sn6QeFm
xZ+1z6nn+xWpa8ugg6uunRs+o5yG67MEJReJCkFi/qWxV5wP71ISAIpGYFk3NZrn
v2FsQrhFip0nsm0ZtaF5o/6YLNxw7dJ9UHbBQxqj+dEuYjs+L4e4ve/uI7XuMnSZ
pKrbrqtUbEkIvPbnnKMpmPTaawlLb6ojeD4TSL1GxFxbUwtkpaiNoNW7ScDRe8LR
AcHER4S/o/zN8gLEMJ/n8CWPbB5qQaIM/r9QCw8snntAb8OD7Ky7VT3tLoWC+rro
/LHfavLvxfcX21xpTXw/qfWb3R23URtr49ervqej/KAJtQ1t2Z1ReozJUJm9szeI
TyhkCt/NEaiQ2gaNyyIiKePrNqHGtfoDKugkROVPYzexpPntLXpjpOdQZw9ZMR1F
e1Iosw2+z8H+keQGDmNv43b6Y3qcSjXEukSh/x6YDnLQOa348/hpK5uLoFRiJJLH
pelbH3tRlfbcnu7TOv2Xc9NzQZvPA742I6OoZbHYhwtk7ofRgJiyxWZCi5PUNJwO
CXCd+APWWf8RxEzj5q3Eb5zpkQmFp0TO8hT0oN9jiK3mMkpdR29+Q/vOnlE/RPOJ
DcLchh8Q27x1KfLd3G6islplWCN4SHzGvMwcFASD7oLp6Fh1UBB5AxbWQvkIK1xS
UO+/pE/3pZVsgXxBau7E05QXLZc+bZ6FrZWrdSlaBSwFngy4j1kR1PqDVS0GNcgf
9ehFL3TuzlpKHX/33gLaGo4hgKZvJ8BLHTGoAkLu6bC4kMzZVx7MFm6dBOsTSbyB
lifUvAlsQDJ8h+UNGPcWiDpjRjlDa7wuuCko2BF+bbUYSx9kJwlSo69EEjcGWwqS
Z8ei0UGr2sw29K9+PpQD2tIVp+H0OsMh9qYTiC31g8skDj9ckkz+A50DstrkrEUp
ynRaaln6b9pOGN3LEWwZfieX3DtK4aHwBIFz9eRwTDbNzaOQf/lUDCLw6Syij1mR
zFAOANHgwyWvExJOrY6YjfDlMDjhZAe5Sh3lmH3PsfConNY33WEsOimeEJeBX34b
1qExdqcl947gkEB8aiPDN60NQqcT4kNr05c/WxgjT2L7aXo9VRMiqtgzRZ3wNF7p
qvbkGJ1FNHEsmJBB7wRvyUYF2o9OEiy1cklCK8ljKfGCRWPBStDaOyGNkQrRCUPW
rhtcypnfaXXvmy7hSLGyldr0HQAMa0ySCIh6qzV3VhOmwelsvcAY54jhA5Cu0kz7
1RYvc+KaoSF3cW3RlY3Uspr2gfY75oDCUQuY1kgGiyVWjzVlxTcFmf44ai9FWkd8
FgMCACTEkPabWKn6mCMyonbJ5nVBRvfuck0kEkk2Dq1CgV8I2yMFaMIKqY/PgLWn
4EJ91KCVe2M8rLboVBXbs1kracpd3YTnN1ebYniH0Yq3jJ/MkpGOcKa/rYH2c8se
GE2XNjtlhrdzkybGr80lB+/n6nX+/WMcGH5g7nnOK8MiNA8hAYW8yUX8BSYSTUBX
nHY0b2bqT0psLCjI40Q795f7mKEl5w8VUqrB/FEcPctnwSgE63ALDENpq8Y78CzS
DElc/Ppyfd5ISfVQ9f3Erl4n6V5i3smVVxFYh2bK/43/CN5XHsCncjqWDSTAP8Ip
fAcD9CmNh62z2QBnrmGlojrnZTAsKYdlxm5s5DPtg78C3t4vLUJkG3UNTlw5XyW6
RekA83Na7zMLu/eOgYe6hhUAc4mQOWMSFAywARlYXjdsPGnNw2vWJqKsO2o3AiqC
Hb/HQwiRaDuaiW1uK9gmoMCN8ck/VKBfxmIvKZ7O3fP+v4CgtLD4BjGJfShl8zQ4
hObuE0cyYEOXBg2kM4PWjN6lLH2mIqEbSZyhTDFXgktvN9eDXFf4Knsf52umCWin
ixd9KCIH0qzwwKru7bOf8Og2N/5nWJY5LfvfjaTe8THK5eL1tYimLok/K05qmDP2
Sh+IBK0fOd4o4377StPUXHVkONf7M7lVrI7kb7KR8hE7oto2tblTr2HIs6I/h42k
+MSWw29W7o7gTMSgyrlrh4psrsZ26kWx4aC4iNCeeAwwJabbx099cQUwgGfg1OI8
oBffUIXtTxePB2eSYBLXoo8GG6fr34p9TReZvGkisOOJnKtE394Up8u1WkY3tERA
UiP3/m28eEja4WYjp9bjrgwsSDopKJqjbCaaFuolSXImXK4LyntNGwGhy65PhWaz
d5p76TSAxWR/JpzFl3bUDo00f/18dQHz9RhDalmkXpWyT9+X5XKJIeNFzv3ilQwC
9I5/FO0HTduMgYePuqIb2vzkKDMC1LrMIQZduPJ9XUR2r6tthcBJIL8+H9vJIwVL
DwLikJMlxry9DQkh9KeempB6Y5BFIHf8kPR/5WAYDPxIiANKoOy6/7XAbQU3zlEP
Ep9+NSTjnUUAgv85aST8QiGgCe0nRRfR3qGHS7GbD1Zj/Lotj1boH2nLepNJPVKj
YIAHj09lsWUHfN71GJunyT5HAWHePLG6YjnuXj6jH7EA65AKe1nMj7lQvp0HBYVi
igYzCzugYXg4Y3/Z2ClWUElcMnYz4ZxJaC02jvsPCoDZyvk14C62GBYubaoVEYGT
sbqvuVp8iqCAtFeDuA6AcbJ0CaFNt3/nsTh7f6FzZ8nEs/sgXEY3TlJlrQq1eYes
ke8lDxlI8CSI21OkIkW74zbfFFzdAZI8L3874rrVEDeo/QlJ1xnapLnmIMoBehkM
QUKsVhDgd80k/n65rpMNS7VZupE5hFZQd6uvuz41mlEphz4C5d+MJRvPU7q7N0Jw
KAXyC7KiolgXxZZBIZ69hme0+vnuPghK7UmN3Nrx9KJAD+jvtGsDkQQ0fS5KaTq6
ru+drySyrTngsoTENPMpAMvJQgKc+hYgvbSsiW9jT3jwsG2gLwrwlUXeKsemF6WG
ac5xjxvtg+ww1E6OLaK6Bv/n2AodiBOq4kIABsLUNBWN7CyikhhkonBVZ3u/TE1F
nPAZXoNh05Y20tLRdLH92Bc95MFkzQJMfB42CneNYq6Idb3E4fMwAIywzBGLYrDf
u1lu88wtssRqtPQwcrDssv1VEddG9kZq5YHPAZBlqXkRNam21HNbVcHN+azuL+Pw
z6eldiYJoDsxGypPTFqtOevy4AM2oz2BizplL3wRVgExW72scySJEvSUY4Y9NjVL
3voO3t+vcZeEd+A8W0kzjnufHfvn38rDanTdAzW5m5RNbdzfzk4Lccs8fDFDm7Yq
dJnwEEoO3n6NAsgD/37XEey9gv5X5j5JCTHrYjs4LFRWbUPbTrsyAOdeKikHbP9n
mW8hpZMPveXkxVWL+d19inRygLOVzXz+PVd3JkGSVh2S+ge1BJtID3/+StccCY88
0qVg8AxkTROwZGkdMBVT/jLQaD79lrHy3sTYGJE/AJ1mVUIrEmqt1zqVjJFjGt9F
adP8RuKA0grdnCDD3KOkyLRcIExpPTYJlJeG0585I4rqK25lY14nmWB3KHF8L/m3
e+5mBeXkjKmtTDI7aN6nqJTAEauy9b7Lht00jaRGNYd69WSwhEH/BX3pY94SVIwe
ZUntXUnfYSrYmLcrdFRuMvZU8ST5tERFPmNED2b72F1DGncosI2pDg8VZTg+946J
m0rKUk4Z1odJfgLrzOPCLUd32fJi1UAbq78vnqnpOzsMTnizXTZOZVarif4pX/TO
5dzFR74MOac2oQcIOFr0XQ91UUePdfFlAxxGUMsa6RRUqE55PMlYAQoZQEu4melL
Q8mxqYwFYRjJpjr0tB9LjSHZoJm7YtX+GWaFLDlVah8PHDTy+6c8NWUNuRzh4I4i
1+gBOJvPOEcZdjo27eUXq98EOcrtcs6x9lP/00RcRTvfvWPFNdkbPs2N99Q8PH9t
uF0jBTqwq6Kr1wA5hBWSzSfk0V8Gb4U8OUrA1gbNvUqWPYgUligaSfX5HpJam06s
adqM7z8waqNyvrLZulbdMtX8rXMaaa7ur16jfBrDOravLjbHEOFPTV2fnxvz2wHS
iSyVvhGE/6EYAmytbLPcDs5417iPjs9KcT83nsEW7BdxEKF/TsRFNh0o8kMnGviR
3/Y37Qn0TpECWZIC/Xhr4SsH3WneSDlWudeGA77hteG4hBhNkWcRLWL4VR4i71qN
B3w2C1cv8DLcDDoHJ7AMgsBYxSX0K808sSzZsuIdfBh1NDPRZOM5Bc0lwxqQQ1gw
R2lQIgnSlEWtdet8D3hf0PcuufAdvjqtjBU7bEvRCjRYlE6WW0YpedlZ1loaWBsj
XOMEfBX8JcgrP5OrZLOYyRFprz+6EIaTFonGH+nSDJYe1oeTl1vUMT+3DMIlAZ13
IWwOsM3HDPm7ECHmzbMPmWu2ndAK6oKpEYF7a4t2tzl4VdSWK87lCVzBYhAigueW
VvlnidAArX7em1JeRlqdREcK2yPH0Ox37xh0sI45VlIe48NdsqsB+jhGih9jhyoj
hN+nQkL5yvkUOcythAdzD9MUAzP4hTvY/NgutyYFGka51esOJfssm413bpn1DUMF
+kEBrgUHPs/YNMZW1gxszscfwlOt6/QZ6Pg5FXcqHsho9VEgbQ1uOLvguS8PQmeM
4gmLX/wKJb39bXSquRqSN/Gy5pIufqjy4oxdmFyczo7Bl2Wn1A543F0hJpTDl2/0
JFGZQn0W4VY9J9W3RarPjUtRl1jAkbU6tMndYPSjybvs6etL9NS7f9LdPwiF7eIr
wHWNNrhTtynT6ULqwGvQ5LimN2OVKsbg/297vZrPsYeGt/NQK9a5AmLPJ9a8e0WE
lKVSDkGGeBLjp2c1DT06MTS9MDpc/4ahOCy1aNnp6KREUOQP9d6nzWjMiwnreZb6
kIP3Xq8kyxvzVW0ZQQSUSXEHLRi5i+G5ctcm+PT9rouml3BucOkv1yeWf9T02m2R
yTHBTBN75cTKruJGDqItzmkVVpUqhpcrDlEE50pP1MiGMM+Air4oR4o8Yjp3jVSp
Ce/Q5Nnt2tNMQW7Jku3U0ZycJqrXhrCUQ+9ZTolGi7aOqrGstySDMOMcef1exQNB
y5BVMDBwPemQjSMgg5LYZP+iwxlqPKesYzl04pFntOm+UK76PcZ+YRdg7RZWy2cz
GuzlsjDvKmNAZPRPL3Hkpulsf0iOoJMbqRvk/qT03SLw2l4PdQ/pdcplzHgWYXEo
WCSsdOx6ox9WjkXMNQyr2U5fzfST/N+XJ6XnxsCIEOEbgLglIXq9srv/N31L5UZs
YHEK+lGAngcs/0qmSQ1goHD9Ak/WA+8Qs6IbK7Rlp7I7p0mzvzw0QBl5x02BNZpe
5zMxcEjOr4XuZbMI5d+lGvmfXV6kUwY8gNbbWb7BjW5PQTDZihahxM6BA/f7sTLV
cJZpdjpAvRUR9PajWUwtdpbFgMP/5K21Mk/46APwKn/M9ckSTpnBeFu66hOYZEo/
10Fjn0xqg1M8EeA0fqkD4lZEb22iLjGwTrfmR0ToEmXvuEVPDX9MLhgbFbQPgtyt
kF3RTHl5W+SxMRe8w3D2gnFwq/7NpssE/WICDGGW4j+xX+lmmG7FjSZh1JuAcPhR
IEwNWO/4d3QFs6Y8w6N6vAg0IG39plSevYMbkdEYsADQI7AAiorvgytv3tluJWfy
aNKiGcBWXrvX0kjLUclYRe7qp5kkskhRtInKxu7OaQtcC87z0ZcvgYEslfqcyg2j
TDR4jAkW8tkrJBSaFOOtmUxS4Y+hgdJmLxGXigor7U+0RDNEtkJEazhnBLAkNn7d
db84EDMi1APsMRPRzuQkNXIlPciVKxYkPqhoMgFGlfmZLaRwKd0LY0IY/ba2Idkm
STsHcDHbMIsU+auPT+ocoti6qaxlzFZCVMXzuEDbkZKKPEHrJxGcFizbX4igJ1qO
cRpuSo2yBraZsPh9WMHEvZnjei9/imnpRS8WQp3bSLkBQ2jIAyFGJMo491kL1XeV
36dCJw0NRMKgNdtYseChTcjstC0vdc9DcYH0cq337iTmPGwMbcDsC5C1qEBBB27e
owrFuqAjl8TcCy7/ewQuGL9rdNURzaxegSDuYC9TSxqzqyDeesbFKT1zyBUAxdux
g5z7UohUefFrn/u5mrHSXpBLPqx8ZQ8TZl8uUNBJq1XQiOoaUbiVITvuC6jf6FMt
N+tLO89oXOdQIULd8GT47yzne+j16xZ2Ug96qn3GvO/B+DwIwYUIOgTHjhx8KwWP
i9/mpQclQQ61fEs6R0Cmv0I7t5pRhw/+ObWwnQeHwbTtemOY4OhXHcaChgWEK49Y
GQFEw0ryf27242I2CIGDDlgOqUrp8YriaHejIANIdReWFj7OWhCNlCf3AY/drsFa
mYZaKNQjKT4V192kZBahCd9G76UDLeHoVQfvBvi58UsHhNH7bQ2Ci6UPmxSsA59Y
X6EOrdXKdGioQiQcpxOBn3Ol9jmd45D3NZTUTR4eCWdpw3482g+xTGVgpap4ZllB
EKgANioRKPIVJUjmpeZnbrjH2n0AZE15JD2ZKzgCCWKxYJKq9MnLftvIhd4EDGQo
UPWmKGvan1C5dynJjZU348Ftk3qHwaI5mSmT2urJMlM9TDlwL6kSuOPJsPPraEw7
JCfNt2NLWpOT/nBq3Y/hYpCqo0u9OeMQkIFb/+mFc9+e2Cum8bbhScdIEiU4bl3P
2mlZS/DtIzBAjGaSwqo/edBl+DtDHzxdfFHFw+tqjzl75D//SO5w5pCWCRbW2Kw5
4fCbXVBANhrleU730CR/ILAupsZNnUZWv25Y1tpV6x5wIBWaYAx6EqR6rzMJgzys
BnqGXxGHZU8Kn6jFMoiLvmaZ3nt+hR8KgnYqzahT5gJkSNrVIoLjjky2XSvHzzZm
WuAwkacYlbZrQFdHONIqgHZOrRB4tWaccIgnAPqn/O+DEMgyuw6aJzgpCHNfV8WL
VXgBGCikDVVfqXGwgRgFp6RJF0nFV4Po0GcCklIu1OTbf3aTGQ/y9vR0/et1DmcQ
Xrctx98kKJzbN2mtGofM0O0tlP98E0UfQpBhjHazQyg/GJdG/IZYQfHbl0P/Rc8R
G+f0vqJdDV/HQKvyVAOrTbiRLTU+Q4mraBC5uusLdl/sYGZFzNDg97G9Xoa6RByc
J6zvWvSkVsk0WoS6sohgRFNrjcbgoPsT1bpqs5bctyR5Uv631PNM4Y6PNEapgeZL
qnDG02yHKg+ydLZSyibyue6ACNeLRnEsVKsbvmtXCAJc7/vCD7TeWRkempxbGxaJ
cBkBcMd34UmJUi/6/vMZz9/9RP2pBo5assb+Ye+zYgdHkAb0O759iXDMnOWC6lxd
hDwhQ4+ImnLuZAUpyNx5i2ftA2S7TQuj63bhOW+npu4Y9X/MVI9kJNLA9uJ+6R5P
8svLtcR+PojQs9JB0WH1fOnw21WSPNrrzbdriDcrItn6astsPwM9Z4xjcO3pIeGE
FyzIMt8o0LdobJmbIfZIrU27pHX7XjCKTh/0O49UFB6rAyS1QXTaEYZxT+x0lg/o
zG8xnAHtVRrQVICDNZLaEjDRZnpYqJt8oYBkRVGwvRyV2n9ym3YCRS3D+UqkZXul
jEfvpKLKsedOlWChoIQowZYXjXWZ15c2+cavjKa2WZDbtANVl0fda8KoRU7mZaYp
R9XNeMRMqTd142IAeFrqfQj41r2BQZJPvtOr7gm1PN04hVe61ZQYp0Mf1N6Cm/+j
shT9a2ROSUQCCpjLxrzSU8KcRUZ8C0hUwyhS96AAEvXySsWVd1rP3XKtK9uXsuQ6
kaAfBY4rSZJiT/vpWdUnsLlLm08jYOUck5vDg9KOUsKixldfVzAy1hyZ2bU2oykb
P0lm5nTrW3C7FwW/m39nkEza3+brbTDwnZuYeB8/JFfkpS7I9Y7FSsjjO8Mb87dF
a8IBW5ioy1LTMcQvoD37fM0V1OxM0vqXAsFc01qxZbsx8JplgdLOEQUeQReDBNNh
LLVbxsNkWtDw6kqnf/Wocx0zgiJdKPZQWGJ7sNi42h6S8GV9TCQbObIEFpc1kdDJ
pHkhdUXl02NmQcBCtMqAxburXpf2PKZFCECOdGNZ8MHmqzQ74ZBCuLFmo1mtnF/R
WF7CR8oI/o89rujoGTgYasSIuGUXOn4PVAIodIhnlml2CT6UxJRqPOIMjeqNmeUC
Dc4WCBQ+dclmZHLab7hA3bpFV0Tuz+uTixNODI08VuG6jCA/SU9ElyCdGhW2CSBn
1mPWyuvz7nM0/lvg0vP1uxTKJSAAL0OMMp85EEaOAG/W72oUs9U5sHsdiMsiAKXj
R2pdt4KDpBOo4l8TMdRTk26w06NtxPRX6iAUQAm5kGGebFisTqrBWLQRVB9b69or
l6BHKoaO/+o8nycdHSM4Z+A49+oR1Dg9NN3JXt+AeUz6Ihbv9RNvH1Q6TqVU4KDr
s1rjD+BCZ5xeqOs1ETJmsLRUhw4sh0vUU4gvGCz/i69qBmLjwC7qrHtnBw/aXoM9
6nWmgscQRugHOJmbJKwvRVPYeANm8bFAui5NOdf5KDO90/s7Lsc0hPqaYUth/kxJ
LEzLFHYcpwdXBCLtJBua/WXfQiHLDcjWa7KQw0xBl/w/UC2KmpPvnKbf/Wm0jKiF
U5PvL+vRfXQx50llJNnt2Dkfzi0z8ZVVy2KgqUCIDIrRonxx9zSyj1Ttp83jaa5W
+5YBx+mA3ys7bTe+yy/MfxJGo+Pg5XZncceetiRzNOIcDUVE1bMHm5C4rvbFK9bI
dqq9HZSWI0HIqJBOYvWXIjao8/BEf9Jqll36GuR66dOEIY8+biV/6QOUso52Hl0L
vsYFS3Qm8D1NrZogr208xH7zPB9gL9UdA+LOpZMRfukucnU5hqnF16qxG9ECcClw
vYZ5py+/M0wR6+04RWoKApkjMzH4+8mwFv9yYBuPOdMBDG67VUxUGmFA/LiqJwnz
2p9l9DNE7Baq/N6S6eiahM6ufQbUZjFCWi6dr2qRZHYsf/96ZNR9hng4hHbWITK6
8qe5auUVuNMuYAd99HEDQoxzH2sQhn1XF2Mft627ReEtDP7nPF7pmWt5pKxO7dnX
Dp7vyn7aUxCJlPfSLv9Xl88v3zGk5zaiN6hGY61e30+HYvNw7/2tG9CuAyqxEZjo
N6px1K+Zbaif62LViEDxUCTWd6QEUqg4HLC/1uo54KWyhQ5xI/H3Zx8vOKVnPE7e
Jwb6RzcKcSlZvW3CEPsZ0o/h/Sa+FRtWDH2Zlas8XW0nWcdNSlKjraoB0h+thyNR
g8DhpW1mPcsVCjR9zShq8HUqSJktCyzY1ShtRxDkIsUtCJexVMaJhOZwX+unSIif
aayxD4wxMBnolOswJH7ftX3ek73GEGjIW4QDMa1hiyvox2lrE2HpYsWQU85l3tDA
gymBatoWfx4L+hvXovLL3+OBi1BoXi/Suxtco+c8XM7zH+EW/9GpORZmJwdx8mBP
isxOkFeJr6DlqgRk3tz8Q5gXFmDxUREqNTVK94FTubUeLFJHdV0hgzow7843qwhH
Yele/m2sjC3ahSpfwPLog9qkDQaNnG7fHTKhkckipBNpyWqPn8WPMCnTWW+Gelq6
8OQZBr8rDLi7AvsRCUxEFCTFW4S01A/tET+/m852oQfjMy61EuVtayvYADxw9VoY
A32xOVk79uBR8tYCXXKhoq6atLV1PbZurUZPHQWs2OHOjOrptqwECYJmaXk9cGWd
TlfEDxyxIFr+NzMAezLeurHUwub9IbPYoqYnorptpSDrQRejBYzJt2+kKFhvdBVl
5KsFdUs7jGDppioUIzbEUTRf42p5fHEXxi++/85qgYUMhYMtaY7nyvFEPEsPOKuW
DWnXKdtoUu+ITG2G9JFFWH37A+KhYHdtKZTHy0QfUTBD/ij0isHY8bM0HEt4Aw74
ogKTH9FmxdoMFg8pKf0j9E/hRJMv35sQZzKOCKysQEDcHVhINMsLcpESzWSeHblU
CafDG3/9e/HAn4pGAU3VTom2lOzlpQpxkUvWtelesqRG9Q6eQ6mNewUQyMaHUvp7
+xrQv6yNsmf/CG0Uh0+Dvj7zqN7BDEW+dQotsoMJ4/fmcSqNjQglcE64rLMgEaVD
zTNka0xuBmAjpH3v4YKcT0Ua+9IOCb7TJqZbLX7kO22mbTJpt9lG1qz84w58Ty+Q
Vu4B4qeZKhDFfnbvJTCQ7Qdx2t6TAmDXOgE4yF/PE3cLJdE/6gdFlbwfl1PofJH4
frNkGzflClDLhWAK10QuZLfvhWcMfdZ57BoQe5y9Xb4emHKOWlp7WZwlB8m2L/e6
jygvlwGt/vyac0v1RSIZjyp3Y6ynoXCfeyG7LpWFuX0H/PlPoGuIhhCWqqMT+NfP
O/zva3+eNwY+x4CS/XUNNRZ2+aEYPF9AmVPd6CEdBdTRFqQhMRXzee4L0aGWEQhA
n8lmhCvQCsU7VfAXBxm/OP+F3Rd+kOHsT8mt0UPiQH1wiPYzUTfSArHZXxlexicf
UrfilhLRoLsnMH0WInO5YX4eThX+56F/FPfjg0syyiHOZq95cptZlJcZzx8CCGnW
IWcOhSYTFsQws2wJpZih5CuHcj0MVdKPUQ8VhMNy1Rhf6pxTLX+qlvKWr1nhrutZ
Wp6b9VZC0LDzhLcQMLYRhv4OqtJySefBaLfg4WaUXtE6X4sMfErXfpuI2qPp2TBC
Ahe2OT6zeXA0YeD7noj+ST8JDOkfsvCW5PphwBVgnAe38hFEx1HI1XToQhjtWlUe
4EBPQYU7DSmaYi8J5Kr1+Z6e2kp43wFegJuXek6fRQ8M/b6VOTZ3ApuWjMQvaKqb
mQaT1t7WGCIC2bWMxrpug3WmfrOUf9u/Gf5g904qDnWaUpKBhwpjHzhyaJ/TGsoK
IxFuJmGqGQwEm0iAtzHTnyy3HkGPlmVmGXch+HqVY8mBa8o+1nBIifFHTt11Z3UP
2LyamOp3zipVdOmJr/m7Vt0R+x/GCyjsrvAfpw7JsWqD0c7xv6RYyYy2UtThmuA8
d3LXidOMWtIx1OeC5EGjcRf3NTot8NKNFUL09bKQ500KYoi5zBXD+XWEMmaPBVRb
YZCNbNIT8/ctQm/NBheEjrxs3VebeiEB/AymLxk19bOnaKE4w8DpmoGOgNJ4F05f
ID/gynZ5eVRlgEeAuRrPwZz/aQE6yltDlOKTb17cnGGzfCAw2r7ikGYKGvlcm9lA
VfLXXdTjCaa89+sAl7hJNMO9K/jitrMieyPmRn2ezA09tw9Tekw1+2Ohm1XtWRao
TovZDLmjrfLRRVDH2D7u2azODuwkT7hKvFa7VzIUupjDmrd1gGoCyTyPdDjhBbfC
O6kGHpNtnF9SWIkOZYWmZ10gLeOnWfW8ORZ3RVVaJKqIuimR37NrIN7iffecbbAh
1+wV7OraXnS9DCUhxTYLRQnZvKRktQ26yLXZ2ThcPFbUeATOQfKT3anXGdc2M3kW
vlgeRK2BBR0HwpLUEAg33nUbA+MLgUWjC1ZFgr9i9RR0yTXefAXqIw5ZBYjnqxef
ntVvZSazrR0qVcNg7LXHBEK+Ms3yhPx+42uEQ66vZ/Rl+O2VV3zCCRjYYClaQoQX
RY3E7mMJzM/geZEb/3fbO8ruvg7qxzWjDv8mocusAK+vJRJN7zZBwLoKlN6mtCSI
j+TFZf0Zy/zVtkE79YrviwOuhSfMBLDV3Q0hM5I9HMDLS3vFVYWBU+nv+uSWL3mR
EyI5UQDIlJvtZ++Mnz/Rt39atq8QYv/wv6Ybdd9noOhwliHMqXWasyspw2ivoRaS
sRziIAMLYqhWu06PbT0gSSkjJxTI0XwFTvs2D9JQTD++nvMhB5Ob215SIqJ9tF1y
lyROGAMsAbuBZxdOMiyL/qdUPTBUc+DqbHjh56UpLnMLQtzfoEdNZHQs2ujQhSyX
lTqbu1Zz3wh/S0f7yDtFSO/kG1LWl4nVc6hT2ixritUim43ndCUoAjzhrdtGyQIi
YXeQ1rLG3pzdec+nywiKyZBaWphBh++SnZApnGWb//cxMzto5FHeqgI+gFS3LKXz
P21zHHxKi6+pyMeVSbq2HHa0NcXcEwuf//rhadIJgF/qX0cq5kLf6kFtD6K1fjH/
HHHXU1XHf26xBXAUbHbB+DdZ/dPKtFOgV81OBPKBcERCyAeCuAY8Xu9mgEZGcrg7
Ht8Fx5+wG98Y2mY//+GXjEGayiM8xI8iRVspkOJv4vb8zdG9HPC3L1PBqXxoZDXr
u9JU0uU/MxmXijYWp6s0Yf0yjAciTDh8X5dx0Zh41VJ/UiTxRXrUkustuHzAeaYb
JNYs59fdy3N9mYhnCy4rFUncADaepwDoaN/avIceK0leeKYqRm4P2ThieE+0Sass
WveVL9hxH0iyekRo0LD93CddjHwX/oum+QCEPw5XDqLh2HoBPtiyc2Rjn1m4Ph9A
6qC3qSET0jNeszFgzSTR9qmwZvRVt+ZBtFCYbqkaI/iwFjgf5ab0Wl8/e0UNP9ZJ
IwR2evKBDtmPB0h12b1JoBLOQ7eU6itexnQEaZ/+dQFco9yIzTHGysyzFq4T+mm5
A7f4zunKNeJKoW20x13UxBQYX6dqFJkr0qc2mRd4L+T0zF8CnI6nNz+aGJGOOkKu
+F6FsYjPR1j4Jd9buOESnsCghWwWyEi6bqH3mjBGnd4Yd+pzWLBRKHKzY0aFjpnK
Gvn74d4gNntAzrm8dp4cV+D8TjrdGbgkFDLmBL41x7W73NB5fF6zqSujlFd2BoNh
D9xJdlvvmu1YoZH+7ZlGMD3AhIr+/2Y8GOd9iGDzBn+RSByEAm847g95w6j7Oso7
5kYWZlFlITQ2hzb2GFZj8aIjgZ5XvuNMmRd4fou4WjId8s5CF178klTI3oONGLGM
zlruSqLvVMXFKpMsdmTVUxAoORwUoFJlXQDTApfZBcPyzkmw5ekxyOkZbfFrGrR1
q3AhPvPsQ+/DqQaj2t13bEuYBZDcBesc91LbYGRv746WsQ05LtwuMT6jNcdGVP9P
LKtbusMgSH2gu3eob56obJDByeF0ibO7h79b7yerblhSbeiUkg2LBdNFISOrlKb1
gD0PFc6aQkCZFY9vHadLpEHX01uIV30PrDwGlf7mddwwDtV+GLkSPBZxpG0IuLbz
m+l11dLqUwF9V5B6lxloVLfph3YuRFKxFCK8hVYwYkGQrNe3OTlFsCG4OuvDYPgx
8mZ6lGrVseX7ER74GrNecJ1gqHswwTyTfHt9Q6TPsQAlXMIEF4EvkB+GLWYvsgvg
mKFJysR4cE9vB/73/tN8n2fzOGd6al7b1+d1lHDx1fNWsThv9KZURcPgwJwEzOSY
u8Z7z3PLreSk3FNvqqijo9BR3O0Q4d52KLoCx5Z88SkeH4HeDkDGVFi+6hv1Vyyp
Id7gIBvuLJyTDOwzalxofapDQBZz6u1U+1RMBnlBVPQ1YwRsQf7bNqwPeeOLEg7T
MtZVzuMKnQnHTZXKb8vyF8bxbTPpAhrd5W2BvYjxUU7Uulz5dymlPM+ZTlWSkN/I
MZg1isCMKsusDxXtMAAoSxojQRwSvQdwMV8JvcM2aCoktydEX2/qLOCmKewa1L6c
eEoPUDPEPL1PmW51ZoCeT0tK9RCMRLlNE2mZUku0n1fxo6bVJWjCe0y6v4ixJIiT
IMg6RFgBTx9vXWu3+GvEunep1tZjTEPLdnL5i5+uRUq/ELqrAiVgiXohiFLJkAww
TnoVx1USLo5divcHptHO9+AsMdlkOfpBHZWKweOR1Ppc2NqY3JkcWvH+U0bd8iu5
NzhKacmYKuaSpwxqh96cpoOc1AcAGZqOdgzop0bvmSn9FH/c8ldbGEMjSVXab11S
h2tV4BtSt+by9vlgb5/HJ7nXkEE5D++krrot3QEoJY6ZB/zFu8gdzvW0x5sadN8r
eYvwyL1peDBTGJfekOWUOzJ4vQrSUfKvf6aGMQT3Moba8KWWKIxpSpZMGICCh0Cr
kIBxSNvWHP/hcfVMWC6qttYAW7PhirmYfxVeBOWOjJ2LEMDDbabd5sXstE1W+o0t
vj91+nvvTx/fy5hkRvSzlfjgdJzDGU0z31rKxQZBBQHbbxqkJ/X44HtVAPlBEDcG
w5TW7nZkct7+S1oSJ+ALYgP92o51uE2xqx0T4V8hIryldH5G507c6EVmD4X6VN7J
SeWSjhZbXgIOFE4AjGNpexu2OjlgYgrHZhGiH+Xx4KE+8oZeLJ2tjDuDMnLLSam4
b5tv6qVBLY/1QjlK/cOhRb5mlN6p7kc1Q/NFe9tRV/fA677tMAfq37DykF9xKaCD
qL0vih/FjtQ16cIOkEVsgPh/9ctWczYD14bMGqNzliQzatgjTqVzbnSoR4YFPBK7
pkRsHyeSI7MfWcLzeGmk8MXRyGzgNROjw8XLaliW1iwG+SUF+MiDQ4cKfISA5uLP
lTgNreafwAgpovgyGWRMbjJKIvkXSuWIcQo0WLUqIpoUrhLwY2ss5Ja6zmCiPK6B
nkNHVDiwKEW6Q4CyfBeX+jIXsGQC2iXAOqBC7lZgwgjMtLbHFnFMglaKFEJl9oFR
0WZz18Gc/zjr5Ftd5qzyokN+b5p+HDdOckdSnM+Wu01Qtg7XEN2Cxpqvm59dik6d
/UrlyTLiMKmFd+6/9SdQ5u1NqBlaL3o6vavh3oaznL803mv/0kst68FcwCtbvXyG
4BdkLfhrdKcmY8apTZfYHHaQkew6HAqaKSfWhCLs45Gkfw7L32ROh24sEivE4OkW
dhlkRhIUW4rO8cg+sFl6B56T9w/oMAReH1P79OXI1KhFSvBiWZmoDk2Euhw0Yysv
IZQDSUx+pt7BkIbbtFNksWVG43/o3Aks/q0xeldLoFvlxd8UjbY2m2ixeF8BlifR
MeIw56FQ9nk85JOJnBI90v8/TFOy/SDXtj/4NusLoj7R7DW0JE4bG2QOgL8LSRHt
i0SNmq1gUlbXTMzKV5aH3v8/ytSCDvYgUR/+iLMITxOhBoW3csppPK7+Vuh5zWnb
atumWmDF5aR3teZaG9FZ/c2yq1RS2TosvJfyRXXOeCYOzU1PvAPDcx0iILNck+qT
RqfWHRiosNd7EZTGd6ytCFYl2CBUJSjV157ptKz3MsByDMDgt8Owxiaxmm8cDAhp
QCLSV2NhjOKD9kLTWDymRoIm/2lmNtY0mJ6h2q1U63MuGeC3AdvV501YUBJwEco0
rf0MoeRStLXCVG29WZlb5qDdCBrV3d1FdWaiXA/7jqt7GrfSrq/YavsMagUYImYP
qQAUrfGcHnfJ+/sALfCXPM0Pfw9kuLpry195RCY8/9k5WqAbPKSkXMpMW8GhIWJJ
ma858njQ02f1tzVn7HeV0IYO8oaWQNqqvuzWDROjenBhym3mT8ooGNaOiNpmum0F
WNLuyuYVNUWFBMfj8necMrp5RBxym6ZvejneFcZ+DJ7gqacfPMNBfe6Qbf1fcMvq
0YLcyaoXkuhx6XF/I5vNJhSI6HiaeiecPccBReOsZE47nUm9UKoWKAid9sRUPxt+
kei3BVg0BDAayHXKB6acm4qZWSuNZPjrWRT0xQLLPZxNyDPpl9FhfyhTIMEWfudy
OnPBmveZ0UcNoCT1iu1mZ3u94l0kiK35/qpIZzZO0hmFMzi3T2Nwmsys89rav1I+
FlKBxmiLz/3nShDsKRdTwdNCe7SvsYxixuosmDR19rfOc6XFZagreYEcosvj5V+2
XqSR00SpqokD1qWzfYAfFFFJ3zrR+n3PEOAdyvSFscJIcyfwrQvobEaY+0jvEyJo
6P2ihU5gfXHkKPSXNbQJL/6rmZDbITnnbFsnAiYxUNvAqYxTt8bFat0rrlWCn2bO
3ywABJ41xPH42xo3GCCtziVFchkU80DItZA9RidLUJkQAZTQV9cDwBzXcDDZHjLG
vY18QRDnDz+TqWWvpjCdpcAl62gtJJfd3phNu1cMs2j9nBNE8FltC+S21EJBECZS
ETgFpN1YCiFvU/EU2ZsYdmWY9B0ymS6mf9cUxp6Sd/B1AET9AJuKcRteWxAO7oGy
Z0m1/nlMQ1POTXjx5q/l0Tz0OXSNIHkxxeeOvKufB15GAiW+gZm289SrfPvqqBAg
mEcmPAbtkKYgihogUESjXcIISC8tf0Hr3r+iquiRG8MoIY3JtGeUffPV54pew8Kl
yulB/htRHRzvPOzuOj6/0tYRoL7Sk3jiOc+jXXp9B1n7v8m9rgQ61OQPCiwF4KtK
nFbwy/S0Km3HEN2+0MTu60dFpqF9m2GOTDFuAnUFexN9flwDEoz4RWyQyzcOfUfq
dtPUGJBfG+tn+MPg7AieFdEuB8+WuCs8vJ5y/xReLRwmnqpKeX+ZWF47K9q+o8md
DlkS33L0vqFinyS5+p7G81YYDlzA5+yUW/gl1V4JtVuYNGgKW9/+17kqI8Od/CjG
bVuS+2CL+hn9CG7gtf3pAjXmbzVgq6NgNz/tlpi0Cx89JAeCp0WA1KAqUcgkBQ3Q
2Yz62OyhIyx8s5dEJ06uMUXaFswry+ZBxieRMYEnepHYlsUdqSAVlpzBLw6RQVzb
c2de64LkvLGzZXdbl7ZNR35VFjhzkcR/AMpNOMpJ6vFIzisvjXgkNWfu9/jtMGXl
pYgawt4Zyg1NJ1jjv1IRJQv7K/mUdKcfOLMma+Xwtf9EAjn2sDgZQzJwuDbhgeh8
JpHbswAt5l9y1aOfTeV5fJuBCO1TLJay38KQQtd1SZHxOJRrZRb2Vjfd2DmmIDV+
7CjvgfSiMPdfMIN1vlJGTz/cJj8Mwh3qEpJKDQhcNwe6eAp8dgKg+2qi4R+2oF5M
CbCba45kotG3xwm6eYgvj2PtzEnAysJD4KGBKCG3nPe6eB5v22/1ivIhGFAVXO2Z
GO1OJD/nEHj7WEhxzjs80qAze3ClkjRpLN/zoN+4/q7Siz+cObVp9SjIPbo/j2nx
L8NKTW2oEdlyKSfp4ndhan2TmoRgR6zLes945Dw1wXZzEtGYSWKco6lrsz1gJjte
c2HUZbzwmu4iIDvi1tkmg1BHO3lxUiydOQw4gAVud7bW9nLISfaVhFbmD5NbO1SJ
wM3WVyvT8p4asRDY8XKNCdCSxLx8nmjEz3HXk62ueov10ua5lAZ4c/v5t+QRVs7b
B+zv2YRJOH19fdYeYmcsHnrwZWh2uv5/kaxQoFuxLYxUd1s2xwe+8ZHkOba/nAeX
kHHJYgcCWW8lII6l7RpLi0bq6vYfx5fD3d8ZCpmlF9HxPjbxa5tGt2nlQ05R1xt7
Qe1u6C2Tm1UMJfbsU5Ah+E8cmFpcv6CJp/vUswuFZDt6wDQKNGascpvkb8ZH8IVA
/pTPbIx1qhvP4K00FDCDFY5gXPzxzl899cbCczwjB1fyrJMpyYwnQB5Tl7+2n5/R
aIlFn92XHxcbMsHRwIlcjOlzuXINPLP6OAC2RSWLNrkxnb4phSjZZUksvpsf0DfK
nOOEgRDqXGu2gJHi2NvBNlHgzWKwZBNnU/+2rmK1+qWJekk4W8t/XrDGlajoLbpD
Sw427g6Kz4UxcdRSLtXSbYGKUWIVmLzR1ovBqN4nYJ4TCe3srIArtWidEch4WPBf
WtgiAwiMcxUx89vJ+8nme/Z8jdc9m1HDcujlHfqLRWpjLUClLkEOsarPA+gEJqho
OSb3FlDAHdhDG95a9BXzi/AvDC0nIwZPCbfxB6b0Z7QMqY+UDx9aRdKTZRwZ9DHC
ApS6RQ9Qi4oddKchveg37qO7w6hBa2JHghw4gP+RX8cUFV5rW6C4f6A52tFxDZNg
f+XxNGuibSOMuHyQ/NMi7rf9ngKrHNbJbXJWf+HVySi9yCyPciZOKqk9UMFhl/lB
yYTDCo2uZgFkzjWXfgNqYNlX3g7ICg2MUjPAdtlptf9X8mArb+qO+6CGuw1O5Mq9
GDf2d0bhG1QMBr200jQW0SVHvwniHlzF7HhUtLd2zMqHDh/RMRYjU++KFROmPphc
53YX65p8361Nh2bNFuzM7t3dkKOwEpCWZlsq+B4R/b7svLaEM3S+/fSDh/DfIEzM
RQPE2sDnfmNs13jbTo7mkLpIwlboVh7aXc55WzFPPlPl1bmekcJk+zqXMqhQrW/C
F7IdvKuXWU5Wi/xDpA4maxuhqT+brwT1DAKf7pTInAlDQ7bVs1PUUxhX2mWA6GY0
1HmdQ6IWcI3MzodDzFhWagScGtzTSCiwQPafO5zg5Il/+kmT60h4TmHn9G/mkdW6
MYGwz2Bj54bWclSLoZPWN5wP4U1WsltEPp+iXyYTgl3sHeDw1pfvDZApw2kU5yLe
6FeHjd6jMzMplbNKKTU/GI4G35YCKjp3Pey1bb8NNSR4HwwjZFtM1WzimgFd5F2c
iH4lKbQAPQXwaVukJlguGWWjez2RH/mHMMWeQ16+hie+dw6IcKECadb/xhhbBNMr
lbUlrA/+7ERgDKll+Iy1BCmOKKhY2IPt/eOwHKk4hhbHuznCyvIUMWfEzP5IDVly
MA+2KEz6Zk38JJvyCe0ua1bkZNtXEjp44hi0Ua3JJSbOp0LUdP5yCU551CTgK0bx
p6ScWGPTgs3gEOeuFmAubVY46LskSzzIVukrLT/AuG7VGiYT1qy1ATHywF0xFZD1
C8wuLDIh29ZpZBtUQ/MypUf5RQTKHkZbVHKW6g6vdM2rj7HQm+/LvjQrLVpDZ0JC
rBu7tBRtQSKhs/+/PmtMMzn4SYIwbhdyUgfzsLowHGHCiguTQeTB4X5guhxK0eY/
LCadThJ1pdCCuuz7GZhs/N7gI2kML4BXWcgh77hmW2gcSyxPygOTgFaadRA9tOz0
2m2/UENoMftTWeqRcXabUU7QWASNB/K1ZjCcSdYlv75c2DlWe/r2QAcS0CcoEQT1
tmoXQpWxXLJwU7ozlGibWnNPMw/kXX4xZTmoSmlaaPHU8nhA4zlUEB6pzZeRFtL+
90gxJU0mR56bF3jDub53Wt3xoDXXMO6bsmb2zWza87R7W5G9B1UujnBo9NeeDz0n
RwxvFbPGWppjD5VvEucqp191fZ61tttD+K+4zbIZ17YLhggYmMZh+V2bMS7b9FWw
1hD0kEH9B3Ae4QgzVgy6pETYDNM1GFup0V1TX573wVvP0sDnjR8F285fw+iw2ooc
9t5Ew+Hb1uR7PuQjm08xXZtFKHLxOTZSfy5qVwR5zPvd5TgoyOJhokV5tG9+fonm
tMtDdrnl5E3BtDtpKjsd19oP9w1RV8geqOqFnO1CMsbaA+p1vku8y/qa+sR48LW0
3ztTXOWitDZ8PV6vjNr8K7cCxsRjtwbWV99Y3KTbZ50k/E29o14lFRnvTR68zXGt
LGNfYmW7aGULfflx0Ojp8gIrxUbQSMRGVtvXEaMDeEQRa/TuP6TIihZ6WJ6OWpq+
TWmvfz69oT5lEM7pp8+aUtCQQSuNj+fz/UitJAVVdAkMb/rHRZfcvpXs1DZYXC02
jvJYwcOIfo4s9U9XEU97mjSoFkjEg6lr9/GmYZwIyUcSW7MJAfZF50+ep9Ud/RC6
YTyDOYfYD8QsQ25BVYPnQMqBPOyQr3jXu0QT86RKPVcSxE1yfrFRNshJ+NioStXQ
Fz/6Z+tPx6dedsLGH4NzPYZZBEZo0Ze8heQP/dngvHu8z40GBwtJDXZc7Go/8IY0
NHhXYUrOBFxEx7gy+ZIGj3BoupD+GbifJroCk45kuWXU8+cFxLXElHXpfjA1a+W8
5MjhD6VClEYiK676AICr/131afhmVLS2rwWU64GbTkxcbLUIvSvi277/mJy7hAjt
e+2+KU0S6TYt0aJc+fjZHswQrn8QRi5Slcjt6w8BS6xfoyPfWhq/Ge3jNUOipkcG
KepqYGJGX99L6BtmxvmQdJfcHBE9NCOeWpF+sPCsEy9KSnvuQn9amLI78+nGN5mB
oBPg9LVQaBIweRt3Ok/aJx77uJS2gayLe8K6KCDj9qfq4mdmKW1zvDq8nvFk0w/A
6Fd42FAWlFaq1wGx+Ex5J95+dtv2f+Xplb2/iwct1LkP3JKvyThjH8Le+dYMjaFT
IKeDbLqP5uxHgtRYFkmAjPJvjqlKYbdy9SIZaZVlrUiF4rZwjGScyqgvilrUfIlK
J0NGcBXlorcPIeKSLg5JpyCjb/moB2ImkWjPqNVTo0jkbsh6rtUwcD656htgpBzB
kzzXQSsqdBH7Wlldr8EqgcbK73TuqzoNuk570QMkPPyGegP4bIt6Rk+jWH9fZuDF
Ru2/UjAvTjUBQR7A+T7TlW81fx8L+SXXLhXJ943TeAt9QqOOswmLRvzD//yH4LrZ
HNlZFoWdhRAsG1crbMjc3cjnt36PnsZNVLWjOZ56Zo/aCIzkvNsHKc8ZDa8X8LcN
vEFXiFoun/GNvLrltOEA5wWdVC0G4Jh0XXkLzMqoErGZH3lngWbeqcuaZwLZ3b7W
SenJK7nuKuGCZnS6NHiCJmi9VXHKOPmIFl/9dYEDzINCTp8+RTI4iN3BIn0F3Vh2
06kavEZgHrJRhGgCII3mZUIfCgCTHq2e5yu5Cw/HYkngrPJ/uXjsMp8746EHbpQ8
WaJQv6LIls2uUSeA/QxBE0/KjaneKUuIxzPAjANPXBPgdV2Os6em+dFiQg5pmeZ5
+spV92DiHQglBf0a3FZt7pcGAlksXzI5KhGKbj7X+uLDY1Kmd678q51eTbTfbiqx
E7AA/rGt7Aru9kMAKdBRuOKCySZ3l4uUio8WTsACZ6ZD99URqdeJYXqBFC+O78ku
OwiqUf7NQJ63Cum0+rBZ7LVdYsYPRKXw5D1yqKJ5jOOnjBNYFvyiEFk4WthnWDof
JjIcCK+93bQwQ7I1qPY0xrX1uwVNDTVfqNuhK88/5WfgsTTUvy99rPrz3WN81nNJ
GoiWu/o4xHQ1cGKjrBFa8q4gu/O2fkvxCzghZ2dJqK/I71c2xP2DdYRX25kjK59f
zClTuhqRSg7wFBYIvlfcTSCdYAQW0VJM2rc44erySU1jkKjtGbxpLXlJSqXEP5uD
JmC4D0+fPFGOyLCSLStqvI0s14SwWM0kw86z6IdDyYl7eF6sNtHl4KGkSKnhFN4h
11w3F5ULKOXl+eHenVdMxz3j4aXbiUAKoIWRlitjZSsfR6QCoVRgabqAiaUAVuZJ
o1DhYWpj9M7rtxT3IKuETiW99tEuTDLE7a7Q/u79xgz2oTcFBitzVSSSo+uS3JcQ
AuzYGJesjWtWXw5cCHkOgUFxb7bhtaxjSL86kHK2s274uD4OUEQZ1rmXdCJ4wBbe
bluXYTrdx5IKdLP6r3hgrELSW0tll/R2/ydNAnvSizK265VD4SF6CxvQZ/pMTTKW
t1C5iTh92ITYADB4TkwsMs/EUoQyEx5NTGQpXS5xpqxU6oSdeXVsMBycbEtKkM98
Wg+7d4ieNeGil/X/fmMNiHyc70hrL9Tx0bx9P3r6cfdxwfjrkoyGTBDWQI0FRoM6
IpI1+OT1jkRbPtHYnjCOdePX1y+OiboqYcITGmSftacrcqQ7NZUcHchcBDigtKPk
8gg3A/k4GHA/bbCky+iaBee6LLJUN0lCnac/Y16sM255YJ2EfAKKGgwNZzWd2ig6
NFjsGLBQyHbmjl8vZkKxouRG0VdC8lO/6vQ6IYXY+K10QVQjkji6y6vSfeYl774I
0tIlEQWhr2ZDbLzsv9x4233rQYlz9CtlNmL5R/2L7q6ZUwX509JvrCu4fHxBPl7G
ZTP65XellCNoWGRX0FLqMt33ul+XTkdlyYTYpk8IJxlaWci8hSS5RsPg3XLgC1ZN
BEw+Y/3Ejs11Pq31JY9g861m/MMTwH7+wRLMwA7Y3F42SBgDHygPO+6md3nGFkUH
GMtg2dhY77d4c7c4WqpwhhA/BEKE92u1tAXFdnQeJnYnfA6GYFmjZr13OjrfWQgg
LCB17MDJjVpPIeLF9WjQus0r6GTkqum0TyVc1UI2hyca7ZSeE+678frNAqAWT7Fx
nkB2JSIHOWM7coK8MeSdi1PaeNlFTzSBEXdvJRRDyO2EMw0XdOAUInIuK97lB71H
KeHJfJl8Xsr6s6WGEzUFysG8EKGs/+LwQtDnctITJUUsvjcj3UBSuJUFhfoLjGB8
u30Vlu48R6oJDMSNgwmbTSIuVbv+DVtqqZRIpjYPRidEtbN31/rkNBqp01t4LZWh
ajfy4CwKrxJaGGbk0yP0FGbfFiku4CW36S7KyvxbtvkUtmymknCe1Dr0ZhHAVmrt
ts0JtKCblzElZhAfimfM+w1gmuGKguDpZWGzvSAnEDBiHTaG738BFGegZsEQwxFt
OJhquMm/cv9OREG7zCvrKFXQDssvN8ObaVHB9yCHMOjHU/WP9b2tR6HTwx103Cfd
xDTIfBcxrtVbwFngXSImKfDFJPQBCBKeb18+zYU7IOttOLQ2b/WEVlrpO7JXqk3s
gnIISMb4bsGvG6vr31ZH6Ej0qlECDBVTXGXsPA4OfCPm2qjaP+yoHmSgOuBizA4w
vq6ihLNPhwWkrkybydsagYve2HIMKLZilIGJo7exEBJJzW6oFsKYZptn2/Dh0tjq
oDLhEfg4FsszWgwYKrOEFdkVJVq6uQZXh/tWZv9KgPF9G+wi3Bsu/5+69QbqE1qX
5f5ngbFhjrttIeX3e3lt3/zuTZZOZINI9h1+/ytUXY8GmAeujqK09fI+B2JrFDNT
YO4D+PLKQN2Zc6SuPtB6X/bFe7xnLsZTTwDbqMEZcqB0ilZqdKz/+F+Qbc94cDnK
iCMmNeOHKQFmQXPND3H86FCi2wtsekU59wKP3Iw2/zsfuCJ+kZUL3xLR+gA9pSW+
7yzgCu+rcgS809WNU8kLzxllN0E5DIFsuSIGjUIDdkXgFmi0Dg6vWNtNMyitdUSD
xo4+bQokaPz3jtTDOtwouOBS7Q7Z1G8yAJ+phDud8KZgTo2Kv1COv+tDCEwrUTmj
kCZulHiE652ngCu1NyQsADSPq/IODTlwqaPE2TrPn8Cmnc1fe0DKvr2P4FbnYzII
UGmrH1isikXch7rpyKqqCIKOosjoGdMqMIV2E7Z9JO6DIC5ewV72DFi2Vvh2oM9m
TyD/ZGx7MX5wDFVdfOh6+GK1zBXdZg8AjWSYJ6GVQ6iY+j8+1FuX1/9afldj73Gc
3LoeFxXvzT0Vk1rKTFtn/EkHFlCsGTVMR5QlTucjtthRzvrVbl3USvy9LAdXyIhB
g5VCaQVFtTjIYYFL5ccyNFHmlGz81Z94BqhTnJCI9z/HiJvkg6+nldgjGOSLQBtt
KtWc1l0eFkEpj7RRokcK68YiXAxfE5m4ESpwxirDa1R55NGRVDRSZ10C7elBA1fp
r5Xx5dGD7kmUu4L3aHsVz/hAjuy4yoOJPKO+se1ssrMUh/27tU6A2C9ojFjTe5Bz
KIS15SlQECKsSbXu1qWvrG/Y5bygtOo9ImA/UrbVfdyqsggwJkPJlXky925FaJea
oJGj5GZbfazge1E73ZeVpjtWI+lbLys0QO/mnlVPvjR/YXJ0QXaEpAZHHrKDmZdl
eyZItFZrChdzZpYDAsetpsLDwqtx6K5YvinWoD4aNoDKCQoYSQKn6xF0zSulX0ck
wSuz1MRlqLBtwVhoaXgtlP62whxnzerTd09fZnrjnQMh1CI3fRUx83k0DDl8Qsvz
eulFsbWyTbPLQM9lR+XTUNUI0iXhdOMkd+b2j1h90OevTZEVlndcF0ehu6N0u9I8
K8WYCAR6+nFDqaHQU3KZTyU18mSAB3irkfOsx2J0TOQ4JRQAJVhFxGocQEeWqAuW
IK8gGrAl4CsF37P8Z5Jl6sAYOm/021KDR734w5SqLkRUhdF3s+7bHFopHNY67Kxr
e8EnBO+ENQfmD0jSRSA4Q3u1LBH2ntrOjgI/2So5YzGJfe7vP2pOKzwoVYPXy14W
q6El+PwuV6JO1SV6KXOlCsPjhS1S/rFsQVWmPKDJuwredFtixDVVeY9rSucKQRIy
f857Mzwk//L/TvAwZAA4ue00wh2UAwab70g7G5taAuR4LU9+enUJI+uoT3NRe7aH
+uzNgSl3m4sosucKl/VD6Rjfw9dMRpMpuY631d5MPc7rmoczSg1RuXvpsiTP8dmj
S+fimwvFqxxEGf3Qq0XvUK6QkKjKXpkL1YS1AFuCZAmiJLx+zY2McdNESvev074U
voP2mosxHZnAZEik4tl10S0hiQZGVzzBrYF9REjleWZLGafg6hNGPdlsyIeB1w0Q
bi3+/VRZlNG/bMoxjhcA3dTwsrHYH5hYI9+gxYa/4I9d9uyJhvqk7TVRxDtwrtEG
Qn8c9p6fM9dwBhidZYWYpjadLTieoy00mZKXSqtInpN43JTKTl1LpPFP0fYJSDtL
P5HJZvzUhJmQXbtpxynf9EksDfAeisgnUwvdn6zve6ZNaIq0CZFCiLPyE/f01JbT
LADZ9H/6G94qTCZ1ONQdABM4WoFklsi3MSquq6qTBp8IERsszv7dnXWGR/R4UaM6
Tmq9oyyIyJwNw1i0KsqE7csAYnaK3SNBv6tt3vLM/IekS809P7++859A07zlPkN4
gdM0md+HqAidPjLWIvk3EUTSvo+qh2c16GREoksBvqA4v5XVuWqAry+Kifp1lLdX
xHpc5Fw85XLA9WlSV0eZGk4Mt0VefXDeY2DwiuqeOf8eh2Y7etBrDodi/uXvApY7
RPTkveqHcHpN1vTSTdkAKMH1Gp5Gvk7khtrI11qMFHBNcGKcSewJWR4eIj/NjWCK
Lykr5e+dhVyTrMxtS95XWqegSHPcxD5asHEXM5An0Oo0nFiKGNPG/GjfUd0jHlXg
1ES7+6rp88LsP5ffvEqbfc8h9BEB/YuB1s6LrXk1Ukyy2G+pCtPawPCcjcZyOBvb
2rPY7zq7eTLZoBAFGqONnE+gUFZ1f+atv9IbZ6M9vf3WkKeoSQYqJPsKnoy8rijn
u4/zCAEEu3prC8GZb+KjTs0Y4MGMmO7OIFS3oIUF5UTgOS0L6LHzP37YAN6V5KBo
ZOhInB2kXKjxH5+E6/k9cGwQhcF+ullMchAskeKWnfpRsqSatKusmF/0GzykDBsM
tN6Jyr6NIRbylW8xdAyBcbcxhAUUP3JqGMfNELMkKjXCf7eicRGhKxe9Q6ucYKV5
WbbZ9t6uFpJ7+zSQRf4aVcQJhJuYacRDX5dGWzZTFAXAD5lIFBNjviI+PlmhZwsb
gAfbe64ZaqSIsEjV6ujxisn9zbP+IyMnxjwSUvxEYjnI7zMjWYyBGVSg3Hk/CD8N
0dNHuUK3EX5CMJBDPHlR0ORyz2rr0DPRTQfDFZ82wa/n4+IKnQZtsiqucNSrjmr7
tPb9i5FHP8kwx8rDnBpl6rmAareoePyPQIr10kuwU44q8OZWruFeCPuAv8vMyNMS
Y1J481/5QDok2zcBKVNNQvOpuLIe1xA3229BXYq1R1xVxbfjYXiwwqv4O+6iUCRF
SyS32QBwZaRjPEctNmP+87X4VDVlSiiuzx9ZNc98vFMTG9QeeImj6GGledqJ/hyo
41oxHGyqe2ug0bYDAVfZkztvHw3hwqskKC+FLGKOJ1N76EFfV51T3NITPxvbi2w1
gPwVxw9FOh5yiPHKj2A8sGljIiXw3bDgHD1Pj4hwiDmK8zqFAf/jp3FilfK/ze2q
sTDaAT1N6kYw2765M3hU1/afrmxUTmUFfWge/3/N+qaEbFKz4ofTsD5ZtofX1xyZ
5NF4rDtF32YxQx3ZFeGQbKs6Tu6MNIybxvWZcNP+At9T843caYGkz77cYnVImfo/
vfY3rhze5lyVCUy+tZAXFJX1R/TcC++ZxglRIMIe/pquSC08A3mwa1lgNENF4eSm
/CkG+qNVoGe/7e5MpChWFdQK8Bn5j2aZfNxsC3uw7/r6sPVfHN/rJzDM0p9syNjK
vkEPPN5vgz7nlDeIGdoAYcuWPqI98Agws+apj+a3FwJHBGxuGCyI6BoiJj11neop
ywM40h4VnhYGNvfECvO8Wh90PWu5xk98rZ7R4g7OQYJ0Fonm5i4/wf2ZMqDxGycC
coxeM0RIzFPIAoc4EyVvJulxVFA6szV5niKAdQAMBXce2uzorHpFogFpopzL11hh
1iw8+8dfKi9PfdXJt25RJrZcZeO7J74O7jHpAqU0faPcOqmW9F/K0iiKoaQZd0Zj
wg4l4VXTIPw00AS35s2G0Y/EJHPbYwj06WbuAiy6g7HqZB6wUnKqF09deaffbWsa
D+KAbTqMWB3s43jlQCWHhwNVTH9IY4/hoqcUG2pIO5f86qu3sTm20wO1BV9z+7OL
5FFq42XAQOM8A7MTS9KZvi4fC9rv9O/rvx8n8M7CdnnmOUERW9acevdgZQR+HxDF
qYovzF+hCa387Q/si7ytdl2F47Gm94fXGEtV7BvMYeTGRKom7iJM13bEmcQifh5q
UxWpjcT9m99NbKfiAbST/vkTA0EgVlvhj6a7LTjEEdJgdvzldgN1hc9o2GUstOLI
oJa9v2lJ3f2X99+bC3VnhBN7wqlwV69z/YgzE+kSMwvZpC//5dS33qL0frgL1SEi
J63APMoIwm/RVEmZehPCOZAqOJC0kM9EhEj2rD5wlecmIh3os0NYVUahqJwvTqC1
El9MsJjIPDgDqR6QYlPSxMLxGsfCxWXXHX7E8QIQAwS5kAn9iKrH05NGiF/etjNp
7C03bNHKLAkotn1Ep0rTtVKEcwQKlVfWkCVMkzSDctCZVAbYPDghN0zh4bzLRivA
uCDBSpOsdQSWrAvAd7S+wJwuyNwb/+97/NB4jK3yuMkBminGakWyJhROcIgwTv+m
FBP41Ykzrki3W1f0yfWv6283Dt3zSp50RZPJqduwtMmc3lfyOraMmZUTBKESI0FE
hVEBO14reblCXFaTm3oevwWOVHNRym6N4DMASv2L3tzsJHv5Cn0FjbCvTW3xaX3J
3q5qT2Ce3vsrFHgvd8qoKRKInBZoYhKayhhjCSWQMh/0EvP9M9c3j0gUL9tRbMM7
X+l1W4BFjiXAPoDBbM+86H+Zn1dUPExwVCAJqQevyY66R38YsgT0uHxhPIvtpzOq
UyBxwoE2MA04wBUH1tEERFCsTVeHQ3Y/LDh4OkBdkU7oKI1o3DTMZnsCT+IGJLmS
RhE7kQU768V4k/3Ke2UmEunPM1JCJsaN2/ZsUWTEk46rGDwgUqpZVcNeXMX1KasX
i6ozVBqBByCzsXOHxdy/qzWacpo8jn4eDrJbyZujwVnT29sWppd/ejf3grxmSYmI
JIW1WOD7La2G5ChzbxtVp9RbQg/y8KlLPPsIOgaohMDCR8eRNBPncXRjj0uInshB
sDH2UZTBHioDIPwUk+ZGztB7QI8OZbwzz5tMZPfJ8vKGpPo8QTm4YJczKPS7Z8sy
3vwfuYjvIx5QXOoENvN+O2FLDMdMxrIHRVUnfNEpK52ZLoYWvUpruJmhfo5Jb6U6
W/UbFsmkjXnIwyPGho/2SI5g2VDPLh125AWcMMUcagGPcjPNgaaOZSREBjsvBs6Y
u8Jaa6FmJsD/4QIWm/nX5hBg8IWnG0giXYPyEmiW5/ZMEjxLalaODXrtpBMTTZMq
l5XHLMTL50K1W22hDDzT+K4pgOjXJXj3au3DPLHzGiB9wtR05L5TWgqqCgH721/F
ZGfLW8Hj4VDvxlRCyy0hmYwhaRDS9xbfuTmjxAjczYiaK4Ze1T1SAty3Lfw5kLFK
6Hsx4++15hvAZIL5FW8NPv0u3ASHSvXOhdKVuEswjjgkcNqQBuVNR3eI3UVIsKAR
lec0O8ZvCUlSih9mMlrVCOrZNCSC3A1tEN75X7GVFK9D/dCHk9KXS4XNPyQG/u95
gtXEhynaOdTjIwRGVsEz/HSZVQMAAcCeOPi61lVdP+H+VXY6hC7pKav5fZY25sF8
liF3z7x8QbJLcPpbTRX/uzoulOop3GOuJCiHEwZ8QmpwE51jHFliz4X+OegXTzCX
WxrL1crKKPHOsTtGlHnYtprtpUinnm1wOKk9dAl1JBtKxsMFnxNZ6sNteJNxEYVH
Ab22FZa64RV5wfdoHH3lt59PpyEK70tuApTfuMj9BN4kEXUPRZ/h2hvBX9XGhtHm
l3c+l4rFBCDLQxHmsuv0Ca3DXyN1AcqQ/d7cQYeyfBCbM1QY8XBP1nUBHLu22jfu
GHJ+LMyfBTIgzO79iE9swuSNEjeIXhWT04VCsSJK3DY4NdduodEXfa9mOCdVNbzi
voIZ4VEmoBuPzeuvStLnX8UdS0gO712DkqPzXa2mI9yqWA5+cDNMGL2ipslf+x5a
j2TWvvcdnhk5XKrcAdvsk2aiBfzgD/z/+xdpF3NxVBSYwtCWP4RVRnKJfCjhHEK0
Chlo8omvsb+9BTh2vlE7B44OvMR51ieA1guvTtn7spZhOrCqJesQYBKwmkVeyG8Z
ooNMOfhZAE1VZwP1+iubZRRHYx1iIVkXKTNuLQlZoEeKAP8n2uZSEU3sY5taq1uW
lVevXYWu/Qg2OiStFSSI1vAZuPmXHIkp4JKhLNuJym1oBHIcAAjMG1gsLEwI2gpu
q1AhaALUAeCbIhCEPGh+Jx0qYiNVx/4OLBqVZsrIBpqHr1cKpOGn1d4fu09DUqMv
5SMF/nIwsoOErwVKB3wGQp8U5XUtdMSDsU/IdPS/vD9z+joEF7y72ouJTqeAb30n
K6tqMzqJ22SkooOt9mkXyRXd2DjNMvKyiT2iZetqVU09As9YkiHHn2pwveSObv9C
St4i70Ey2JovKsXnWtJZ53PVfTl5NPom7WR2ZOEAz7ANh/V8YIThKZeUcaNVk22N
Hz8joC8OiLv3LWdRMiK0th5TBEWjo0+++GVDv+R8tUkCOvbwN3+oNCKzKzNWC3uA
nTkyFJ1ODlGaCGI5UHO03quzHAI+C82xC9gnDgHwGDqXP+Ehrz8aiFmv0SVf6CQO
34hgpmZAVUh29JmbclKfpfFuOgbhOFCEQ0d5bpX/U1aAbbiHWwubicnpdGKo7n8k
PKaDceH392wKvekCspQCpDwWejSZG+8rE765zeFKi+OGQIE6ozkAr2W2M9IXtGF/
Wp99ZmaTGY0/Tve6gXaymhUPP3shgwVNDEDlM+9x17hHOzSlwvZCkddJQQawM2gi
/VI9jbIaCJckhVDXU2POrQdJ3q1onDbovpshw0/nHdDbQcyJXSRby+j3HDaEBuvH
ZF4UpKzN5p/kUEvcqN2eziAO/X3BD1j2bBLULTwUw6THvigWxZVm4a0EX1MMPeNU
5D4y3us02liMsI8+r0zogaVZ/KDf+2gd35eOD3JdO+jGJqdIO0cCUdva7ep7KoJa
ZGLZxHHj9xt6mTu/DAtuETKZczy+q9jDdPm0hP1dB+loWgHwUIUHcvHZ2g5w/fWR
E+SddSc84TCT1q43sORrQ1RsePPWYuhrJWw8N9R811JDxAL92UAJxR0ILYZFc6Ng
+74ohgYLRKnDxgz69sLiCc7Vsj0kJnRXUd1sakkhloM/qhRczmdrdHUAfpNO1m1d
x/5BtnJmPdWbV0AyCEiJRKKy2Z+uVPoBXfUU996KTnDb7MTdzOpVD5ZXSrqWKAbE
gMm5aTAtXqY7O0TguCaZQz/F4xvRUbw1hwX70zQiCqvj1bfolqJyQle7bp2ysGlY
5vsNuaoLHYLU8g7iY2THW4zQRd7baqBv6qD/UjLkac9IZMidjtP6JEaf3GvWORKH
BbyfXSK2rEsIxZiimOaPKJegZLDM592QGA49Mxal57+svW3KLpIkLSp455nhsB0Q
dpopTIuOF3Wt3CnQTEoQSbhKNDdug6lO6pAdwCKEg6tI/hfgXgNeYTA32e4mouMr
3R6OmBPeRq5FaZY65Ec89uOwsEmXhzT38VOm38xPXauIHTL3t/YvzUSudQizsJ2G
JoAm9ZqJ/0ucJ+bJ5y3fd50QKbjUSo0eRFGTjhEwsWiD4xxlOzID4x3GztAyPLMu
pKrC2AAytrpdcVmevK7gPqsdwyu9XTVXz26PrwhrSf0RU9HMaitHPKDuG633xnDu
1rLpMKXXcJT+Y9fdfnu79vGLUC0T2agpCgvU3sA77IzKUKxpq9K1QwTxq8fyB9e1
e8M1q3oXzHLqYMclGs+TKPPpYyFWuc8J62cSlP3oM66KmNzD2W2gAp29+6dAT7hh
GHrf6c1b7bWj/dJ7ZgjGJs6HntrAXvfRc3yMlBNkmVD/wHB6KZesFaVA2YaFszXT
Ds84xYTcfqzNwUJfi60aJa2EotAWDJ4Yo9Eh94k/SNvdJiSAe+w39dV1DmsJMa13
rhMmXJYrPws4f++1it3VZKIW5HGNjZIz3FMkG0wRM+9fvGxcsl/cSz1L9G7j5+6a
be/2/E/o7oISd6NNVGaAUUH/Ctfnt4LbXxMggphW5w9/PzCixAxCLBJcF2LVcuKq
4Zc9gFT6km8/M7hs5x3Mn9hG8lV9FL70NZhnxcAZc1CxRS4y4BnnUma/dCA2pC/K
Iw+EyhcxaxHJmFIRGJjrAAeriS0eVJ3MGQ1OJeKv5TuhQQvDJsNHhv5s048X8g43
vzlR/Dwrro3IX+yDlcHGeRTOxCbdv3ZANv7q4piOOW8pAazjhOs4305IxiEgFw4j
dfBOZzL93nRCkZSkecbHo9cAr0VnZESPDIbdXV2ahPvf0Eb2l17gU08kHhdtHlVM
6hnWBRTa68c6p6RircQhgYTZCBsfER88BfEKo1UPVSQC0mIGVTulowMw/huyARDC
s0BtkJ/UMzg4CDMYO+SvPyOyAOdTKaN/KtbIOfanzEQy+2uU3x5eThsKBzGLY6RQ
lDkQKn921ylqkkWRXuAMa9W+VCD9Phkot5B7P7iMe/vQg/QIMcxqlTWIRMh8tpcP
ciu3fOv7hAFUVUgkDo+gAn+ztQnHInGwzqRi0Rf293yVL56DLKTbj/IdqiCyorPs
B4LyEOUMjRU0cLaUAcPh0k+49tNfeiVyCyMdlasN5MU7agBdEqIMoxFeTaUN3rcz
D7f3TMEkzQlIz/oU8yXoOeZU5FpBa4HQab4eK5MPxMXybAmLkGUsvga02bSDWW5t
ANxvHyjrx+hlx4DzpqvQ6+QHRXilOChkDV2M+Vx/hXSzcDoOtmHCZx9GHpWvKf+9
2ZBBC9gbnQT5XQH9KXI0+TPeMtObTPo5mD4Cbc8lsxFq3P98Bj32TRu0cS93olIb
mDv3/eubywYiR/OeXNWzgZoM/YK1NySbzn4G52HZ0p54kk0ehwdal6sPXTHUT6jH
VHrTDxr32oJurqWqj/C7TxRg1P5keIx1yOCC3dYVdFnugeZ+y30hL+qJBgmZ5gnI
hHy4NitmZ6b+YrTFAUoB/Fv5X+Ho69Balp+IGcDwKoJcO8ofZYSx9n3Yffia6KB2
NI2cbDW2PY6IFZZ5N+Y6y9e9YaLq7/5xsuwI3VDOFcwkaPY5Z+9U7GY2rbVAEwxo
hXYlrxixXQcKSDE5bV1ytKLejg6IjBXb4w/Ye7gcYz+AxaD5YikN/qK4y5kdBdEb
xnjK3PP+ThVVArmSImWZwN3ZZXwdgXiKDV/zjfhD/yAgKK5O4/aPkbP0KjxzKpho
fYlfqK7a6Kfjqvg+/sPkoHKwGVryLADyxyhffCF4AZy7G+KTQJ1vD2Czf/OUyc/k
wuNfK9LmnjYg04Y3iQAR++/rhHtAVkcAyyLSB6CyyH11694fnZSXKwwenM5xMwEv
/61ZGSyCMcVaiBq9v05ifXNHOy0HNiXzdWQ6F/hmpq3uOEPStxygGXlxeBkMG7qk
fASX6cjUgxgx7la07tNpSE9PdK9q0DJu57TEfzUHl8Xe8jBPlxAvHNv6xE+J6qyD
lAAuyBBSzmFUQKCzBC79g0ad7VI3dLNFznaExK8s6T/45H+N4d53S5aNUodSMTc2
3k6S6r+9ndEJjbO1WmWvd5JpwG+mY9727JaTls1siv/OSfOArtPk1Ns0RKZVB2xi
LiGly/7oPeVfgea5ot7gv0qenMbacW02mhi8A+7VJbuiF9NR5t2YqEVbSS8H9A/g
aWwbbrOfYz+a/ZtKnZWBd+jTShUKRSEmnFzN0rOLAy7g+NVcroYIqmGXk3KFWdAl
DMIUzK+Ns4GoKeJdh7B/1VNp1glrQevCOFyfV96pl8c2ggmLkGJ6CWaiLvdiJvfe
24cobGuGpCC4tVEQdxVWlJYCdbR+WYBCXhapbSGW51hotrP8xTKidlz9gSrWDjio
khWnRF08+ujYeSzt3lUcG9D4v0VpBO5RQQ4XFZ0H7n6uDF32PTbWSk1dC0VOsPHu
P38So3pl1GtJ2xBzRYsG0I73WtV4BXmDVhJjjap71DEe95evYBZjx/yC9Nlrszih
9osntHe0dSDjG/V2Z87sLEXvSNmpXO8cyKPqRfSEPDAYAM0+WHnBfqvXhF54WytS
XMbPFx8KEET0O/tEED6x2RLHFhKwokVzIhvn/Rc4ngbVj0ucyt2FE/2GnZ7PS3hb
QxmTXFm25JFBGgRyet5XopXmIpX2c5N7iH5X9yzFPyZAovEZ8i16EUYo0AexVqW2
e//aoc7HULYzeKmi2jlewaH866q6r8Jb3Y7bdTvDd03b5Z+F7IL66yuMOMOLg4og
l3iqHHEmsmIBwQDk3zMqi3KN65Yw3tHjvo/CFC4GMxD6AOwAL3+6ciKEOoZubn2v
RSbGbsa1e/jKG7Do2oXulkjS1h/aY12JMxDrzW6rzjd+ON28+CKcEva9MuLRDL1R
OEB3MZgc6JBcPb8A1b9hxXR57oLRjF8T3iQLiUTyCkImqdnV/pVSAG3cJzaxOfYs
oSLIPU/X9J4AFNL8XGbqFiRTtdDUMa5L5lh6qTc1nu3qHyJdONUt1z+CEo1g/iRd
723XRovGt5I1h3yQW6fDEEIU3slRp5B4CmKZvWCET0ViqQp+FStfSrHPtf85HW4v
whwsVLEmtlS13AILVaYutedHGXcRUWDUk0MvRhlaEmQiRX/PWcOHgKsjKLL4Ekxx
XzQt5OTX2m7HDy4mBf88Rk1xY/GAShvlT0TVmpgVSyR8oiBlzBd17uCzq2fxzSPX
9pzX74Cs7kegK3s2Ds3zk2x1hmlF//gs6EEOn5AaEY2vOi20KacaNNzbQsp6LyJ4
kkcxXk8o/SnBrdJHBdtgPyhiI53wq/71eHvZXOUsW6EJVQ4oJaNYJgIFpySlHG/A
luVxoIJFC1Ttznd3YPli+5Qqoyt7KSCAP5ZCjR5n3Fp1ilxsLF/5qjM20qm2ATGX
JoxL01BFQ8Ado4B3gIoBY0UA11bucRw/q2jjfRZheWIwffao7bJJdJd0sKocdbgy
cNg70Gj1uXXajKp0fW644H1Lo/5JIYcUWMzyrREsc82qZ4lRHTVX1nGL83gTW2n7
W+/zwgZa8kmNdY3H3CIg6p4GSSXMsPr+uE6UfPg4+SmjhepX4IkYCDChwzEUuXgI
KrzHZCTFgckbCXNvmUNk9iH/ReyXyxMJtUhtmc72KchmN01gHsTZe5h8Tk3pmksR
to2BLHwM/ikGDbj5jwgA+Zqjn9xqJ6kH8MCyLmw4Bb6Gv8anMfBjfMpaEuTdw0TG
6OGVkd5ACNfzEq+Yiq+oYnXPbfeu+G+jfAVnO48OCYpBpe2IU46HhMSx+OLO+MWg
nVz6n+xeQtYhVZDlCFrOaHXhNsfsMUr1n/kH4IcV3/dqSoeCjxXElsJsQFC1gs/5
GRw7e6dRIBAKsR5fiOFTA1INJ7DPTRPJgtuMenRPDqPhU7ymgPlHFbmfPzbhgbyO
nOV06/SunHG8V+315M3JarcLhn+lUmJfcmS37RiLuGjcT3RVN9jk6HV0FoAuzPrZ
ioq6ybCA/4QxFkrivS/2J3v+aowqU/u29dgCwseOAZsK9/vLtWm9kLl9oSpmTlBo
d4g7vuIoL7G21WCpPpmvImzdkiNii8vyN8HAWyMRg/vPt7qpnTPnbvBGDXdSXy6o
95pPp8I1Sn6oBFPe/TrzL9REpdmxtG5C2ygv70b+1B4rFC39U8+8t8/DLdh383DJ
fwNvzzQQHV3TEyyKnAMN8mqOn2yHEnvPlVg7+lgQKvV0cy8d+nos4CTuKZXNLgra
eK1a7NaBhesQmQD2lMIPg52n5xJwWKvVGi4MCIWkrwhyBQIzOdcuD2Neqd7/K1Aw
b9P8dnjy3tLOR5UdgGujDpyVQQzICq8/vO6hLocaaqFoO541gI+3JjDxZuMVuTOH
oxtj5sYj3VjOXRabDC3IDGwVlTxhM3evdILn25s2vKs1PiQECOqmo+Mw9yE3p4ew
i2IrR6l1kzbCXCFxhMJcFel/xEzr1XJvNr1DsPlfG1iDxH6o6Fh9JXYc6Y+Y6OBV
4QmYofkC/kyL+bltT1B8/TTnpi/MJTABcIPR7cw+84zOrFVQU+vwg70aF/g0du2a
rI3BuXXhgDmhEy6NG8hPXc4NeWZU/PXV/jQ+vZCgcj1N5HnRRyVU8IJbs15JVgZU
Li0eRJU2nvL66xnbZ87f3oNIltgUajvy8uj0O0MzEuGmZQk0T1X29TzQFTuSN/wq
xtwI4H8T6j5wdiHfVmt56V0CvLKHvxIczgBv1ac2DvgaLjfBUBU4QslinITE2wVn
9TKGhKx0lb0ZJqlEHtlaQm237FaYtIOp2C0RymxuuQZ7bZ+Qn0Ku1qi40dBG7R1g
XhWN5gn5/JFy1836K7uTR/raV1I6i3LJQkDrFcTdurIFpokGfpt+kolCoEQtZRur
TbLXBhbfM66YUjpIorERwS8EL70ErFl16GGlKdNKFfG0y1ojI2Fblra0kiMHLp7y
D5HJmOsqH2aZ5c0f7RAWkPvkuplcjaG/j7tNlxXr6IejEdYc8mYyYVqq8pu2MBzb
abFasNNLrp3HH475Nfh+OaXQSAo9Jb3Jy9eewMCQnMYoAO0cB1dFJ0zQmrwfTpDy
IFsEAI3Whr7XUyD+rsxmIn3Q0ZT6EaiH0BQMn2G2YNhRbZOsmEnp7wYMxKe2jY59
hmppKS/0Oc6Rsm9Y6iohz5oC/GoHYKMF+pACpz2cQ8/tXEekzeThPozE69Lcv6SQ
6Ixurh46xRGldQeYZAHQmcyNxXx2TRvDyOjEDIFdPLKpdWNIeHjIKmNHFY12wtAN
Jlov5xiRUKeoVqEd/QI0Ux/q3iI425xPfOnnX2kEbCu2+SXxsX9XksNtNwngcT+1
0DUEZU32/kngT5i+Hl3jKCE4TyGgdfJfE5C/fos4tbismTAOumyESYvKH+dR5Cxb
wyBCDpUvBy/S+HFu14U/psKQYy+zOQcO/uf8zh3SyzODPXSGBLwqRcSLSN0cGDcm
yg+MI/+91Eun1A8G1+0ahRc8eDWjWMF9UrjyQ+FHx+zAXUbGFMeO12n2a0BWkj+G
hsMfW5Sph0tXXGnZRvJDXD377LHF7RNhWuKhJrtevXJlCPNwAe5Kqk1KZpzC/kO2
ldECWkHLh0oMQUOx5wVGGh3YXbhG6BrZUgKYSt3XaermiwYA13elagbZrwO23uEl
T3/sX3ly3301wKVtVey0RT7fcRWYw57OgmqoHNXxA6kaiY3mfaL1C/0ox5kbUqsd
Qb7YPVIxI1cuFIUx4fh0uqv2gnJrUn/tf4GITvPpoFLzllHxMCnkZAvBk4WnfWkw
Aw0NbDNPN/XBK2HJQ0Kg1PnBtbWEsfKPOtHWfj9pVSvtYY65nTfyT4cNAw5Z0Nyb
8Jf/vRplK0zhS/TIttk7WnECBKw4YtjeWQSoLt44+fZu8c2MXHRVVQ2+JwrEyI5G
WKCj6ZRfyt7KdHHfIOtKMP+bB0tCANcGd2/VArSxr3HGlosPqzo6y5Gsz5LSiS1f
4MesOcwjxVMgg/Ci7Dm+eSx/LYGZpnrKD91J28TMBrs2nDD6T4svGYuBLRpNzCuY
w7MyWHUQsg4Czwk5BQnxbzXgZlAr/sccf8z4zZCnCsRkkzBz0dHn7gruTcoEIV9+
MDBHkVYWhSmbwl8wwiY698qD5ZayxMeEak9j/3dapvynlgkyBMD85/xLYqJOFmPH
T0MiddIaBwNmWL/L10J1LTb2XvOKuzWrWEFpfYRGuJ7ZKeWLH3fzWMSkNuIg7K09
DIxYffds12N9tjkY8I3PHW0gXOuByLrTJsvuCU+GVdjgc8pluXROGRKOj8AaJ6wq
qhxbLR3526pn5POCFHCfK08MF4D43MEnL8RmgtMzGN/9Cu4hjeNSYxSXCDpvDsjt
BejC2Rt15nD5JSE9+0o/QVRlws4zjH6Y8aIoizZiYI9N1k6tz1sOvcMfu3HmQ4qX
+apcOj9Jp00L61wqnPLD73PPpx5wC1F4Cnd/hXpFBFJ4nsaEptTDnP5f49COicDN
T5ixYUB0q2YUu9HGFpUjonG5c/oQ/Ic1lrjV1eMUG3neN3qSgYlZeTO3DCIeyAGV
KvKs3U9Wei0U607QA5svlaOXpPTyile8SkJwtKzpb/3mYUAMwZAXXWDfY5A9rUCt
xFkhAMH1l05WMz5ukUF/k6zxeRHs+4Dq34MKY7SU+g6Rw14gg6aB5hJsrTMKYwdb
D/JYZJw6nqo+CIp3ogx/jg7PTyDwTldsRv7q6QLWZoqYCc6WARVwxoGKEknXimJw
/nB8Dq/LU2wjp1gydx/hj7FQuZLOsz2C0cmNnFvoGWF36FpfNuHOCpHe0FwTSGrj
AvSXRlJW8PCPh/Vcj+1vGy861or5wlVnEhRGlMvVzzyUjo3Nqe9beGAYPmNrDioe
DS+DCe/JAtUS1gHaRXowLqvh3p5Y//HHUMuhYEnmxx1sia4ai0NQnA/p5gu79OQZ
w8/dqu8Uxc1WLhCnikiHoHMSuIa3I1IM1f19s3PRRq9XVghsg0Dq4KyyV8KP+s79
Yf/nDXvDksxv+NQAgXEFgH0Bzdk5CpfFVbKRPJNu7Q/T2kvRFqFlF9boKHHlVZgH
UpWlikLY+KhLO27zuJG7REzcZ+m53pd+5PM5PZ5jvTGoyBEshmWhC77X6yCs8WWS
Vp5nEvWWcb3G892WKnaC1PZ4aiyPX0vaXUSvJkSuVAIaJ+w/RJySED+r+QGpDSgz
clu+RzqzJoP9SvbL6qh/xcyYH03JnOJQUtWgFlsFz8v0vuuHU7b5tOKUff+ucFeq
s7CBNWGWZflvy4VzQok4SwmFqZ7BjG80NlAKZnpJwYKis2stHtPP9rpEjKLZ16sG
ON3jmgG9yTHQrt5LZjyp0UaKAN9r0Fypp8DnyCYUONzTRoeL/aISGTeVw6opKASP
U/hCfRBtjNzM2OHTtGDxFpABHDoBzmL3yJyQ3jXfWlRA2pupqEDP1a5Vck4IelU0
NSDuUHfM+sVlertLqweYhIBd1Pamv8D//KoY1xdQ5LgVQAXjo9u9LmV4NlFH8X2w
5TBLYS8CYHtvwcxr1U0M6WbH69v76RmCgPxwG44YDD4A8JXyFcxMqv0xogqlASm/
vnhf7GDhQU1Bq+n+C+B2+sV3IGJnMzdXa3eXRA09ahvIwuvt1WBNmKN5+NfPHwOJ
Ryy+x75zoDF9MTm+xVYYzCRUftfHZLPpeEOwN0EiQ3T70wJq9QIYmRfNnvSBm++v
xJA6yLW7UfTRaAYZqwpmOMnP/MccI6axSJVelTxyYhnrmtVyfaimXNVYZi+r9Wwx
GTT4nWHkTZJWBvVPgFvnIuUKizwmKVD5VaCEJRi5RdnzR0T2754f7fOdH0lXIKuI
CnKZbO+pcvWr/Sq077aTTtOKktDWIHmqNXpW+d74odRBIwbPFaHQ3FO+YwmfxvhN
Ay3nnXbmUMqBiux5s5ngxkAxF4OBwoJWCFc29ciqxNxsVx2hOjdyC0IU2QUT+ow7
UhtxRJ6w3vvv6Vn+XntZq9PcFAHcje6Z/fYjCosEm0P17COrKA0QAWtUcJuf7+BS
U3onAjb4gSxxUcH0bNBm0g0DqzVBGxkXsXdaMfFLWhqLbIxCT/VH7kMDIgSGc/cg
J53wCpVxIg/RyH1JgRkk34spcXZJGQpfz1izR8pFGDlvXEHKvbQKAeJQLLFFhv7X
SY9ohU7BTspxZmLcNMRuJ2zS/Z/i4HF3YSx8odE9nLmw1BGFp7uMakaatsHZYKV3
FZ1cozAGB08eJSk+ZKRj/IqIcP4t1YLBgyEn+QIsQ4YJECuR1P20bhkKmvWK0j8W
F4iWTcKUmE8EA3o6AtbZ7A1S1JMgfUcgM0Qrqc+Q3AhIMVYNrozYvmSOptzUlq/o
AOhdcq7GJUY5yt4MnmLfulOYVy3I9wE/0eCTYyigd5a5DtQeju7zVzIE+xPZoCko
vwe1uPyd+oI3jFfzAN8YADI6+kFRIum3cbonY+wJyfDTsE5hQy533Q3pIbOuDDK0
+H0B5eSZMQcJm8E5wtSDLPnRQcG94lkN6G8kQYSqQHeoalwXt0heLJa/rU6ZSaxm
VS31JtsvXwbO/OW5v0TfmGFSz7NZmOH98n1RNNRE54F+rN6m7XcaR/9YgUPlxmDI
DotI+vlLwx4xDHgOF4neKm/tHRjUnYopII/HEn9kA7TtsOtAcipKfQNWoxFU5sRe
8aaUXrJXmJ3hZ5EajBYVonZvyG13xQKK2pw15GFXlJ4HQUc2z6z8JDcnq8V1a3rU
nOwBmdNDYa95XYCKLB6VqU9omDYwpLlvyVbbIll0Yd1Wi8BlF0J049lR6LsSHPGb
jHgH7zIbl7QZ32f2VaqtsdFhHe8wbzBDNN04yq+/lMIaAUY4pqisByYJlvWGV6Nv
gUW5MAgZhdhjpTtHu5vCppFRENgMcspzZggDGa0S7kLeRfJ/+Q1Oph6iQa77E/fT
8UiOVGyylY2u86hjg0Dq4i1jvh7hgltYD9ui4qg5w/H/XdXDLCyGXgL2zn9nnYb7
ddZyGjnk78Hr2BcbTT9CAuLW+/UBPQS7Y1Z9ILTb9CC2ita3jHgqxDA00IIlglie
EJCRSlI2S+Z0bttj7N1AxhowpWwsDs0kpVR9AQQiNJ10elEeOVZ5j/p1TaQid2Lj
is8QM7cC4rEeXBheDUvEL7L5uDcb37O32SZDThQd2NPuk6UtLG/ngASAdpolfZL7
CnPgn5Xz4SxVFhSkeAFXnSqKBdPcvW1eVwVKN6jDVwMdsGsocoVg7QUHRYoi6W+S
m+JRo7xhlaZ7T+nT8A6S1EBgiKME8b6q2b5mhWRwFYmgRtB31nMpQF3EJPU7fxDZ
yvLjKMqp9P3IIbOiiZp5V8smfwDUUmjzCw/i0lqTx9Pn4iV3RvWAKHme2MbNY6bs
z1WLub1yNSF1/lDaKYFKn9lCn77Z0lAWY0MWN2jwaBJbgX3x7qpD9vUsQX4k03BS
xu1MJ64Q1JPDQ2kQb1oy//JgBWz8f1nsrVi7kJL87lOD4yo/FEpXMnfyJYyIjB8H
2IDgh/Bvl0zHzZ90Z+93HbaZC+arvezvfD06Wl/nPogqLmLErTyAr7H7//y0AoTZ
zFozn9fbLfS65I3kEjTurggaBw1E3b57wYSqZ695u1cY1ZQpWRh4oclgRCggPxb5
vehvpGCMUdsgjzU2Z4DOvtwMuXdMZ3DE4/ucVe33FPpcpJQ+U/4iFe6rgtqbMZRK
+TwqoCOk2RiCMOzM2sROnlyiFbgPXmaAKldBHC05WBtzu2RteD4KBqkgFKo674wc
CquMUFWdWM50zdzMf5SAhOB6QSbnCCgcKgz7C6nhircafaQT6beZ9pQWksTL8aSh
1mVW0AtLFx/ahMYFK6sY1Wk+uGU2xLdkeJ3we2DGnJULbylBVqU4WNQy3Et2VLv0
TdD4g62bYTyZRFszS2ADJrhpeUuLopGQeFIVWRZWFKrwZ3mXe4LoxtNOY9+RukRX
lZ2TJOItAlO8lJU0COt3Qbp/upeoby2npIemZmWwb2+xjvy9M/QRNXX7hF6NHFyL
6tML3C/R/rXBgMKFvcvhvWeg/9YVfAAdsXxVh/zHOLpjgpqEzVa5TqATcnjgUbyz
ezlo5OpzMWLS07W3QD44tq7Potr0OQxaKdAGmb80aPOA1wtENzSnDf/W3Z2g2dB3
uPktZ9zLQ+dT1LLxqPx75LR5CwGfMVfkB6ATJM8aPkRSqpuUnfTXGWcnA/hJ8duc
MNAS2vTXUle6seZegz3aC9GRS+Rsoc7gJDclz1a/k7/q2xCGn4sLcuBgij57ahzQ
bWu8cM1OEdG4Sttz65QA6BFErA1TxsGdXU5ezaQo+GarY0kQpp9EY5aOWQyAHCvv
/EiNRw/VZVbjqRUSyyuiHad+gRx0vSIPgzzSQO89R/kwA6hsc/rlA7jrSXlABU7e
ZZgiGs7Z9/8bCWDy0RkoWU4gD+DeOX5mOIkd/FYdChW2ltvHiEACStmhLmdFn4aF
Mb4RBpGHBIFuZ+SDhDoKzkFyjlqVagto2lZHmlShE6w6XZt7VaWSt0Vk0xkRl9Xs
WQKivChSplf3tGHBRrqacdEsim9GSiZNxxzUairU3WagJ3Y9QTFg2ZB1g/c1EI/h
P/nuStHcGNYYtgfP2/jrNQg7QUdkNDlRUDvjKq3QCUDLrVK66h9k/UlAjz8ljLu1
WJR19ZfIyYrQo20qh1xDDqgCYkrSTrt+jFzLMHPVMXNqOe8X0zrj+TrF5V4RlWyM
92ypDTjr9drzW9cwLm973XZIbig3To5mYk4QkNNgOBc6V9+mfR8hUVz+p6Ifaa6B
7rY/N7jvEzHq0kuYvrwys2Npu8Picd9WVqrgdxFoOzjNSWb/PNmBFmv9ueo7Oz6I
eckchvheOGxWQYCB8buRITCy/4U+CONNyM20uNXMjQY2OSoegF0Xqjv8pSVHqPHg
DLBMpDsymwGlTTyiD08OFZYX8goRTECTBtI0/+mILV7QDUe5FsdhIHb9Ftz665LB
LqighmBZ4yN7cMBFuKoYoAYzA/uUyJXDVzeF5mpDsbEvH1a236gCXyPScwpGPsi5
uLysv66twAUNjc2JpqgnektNu80dahEh+9R70RcLJk/RJZbF25Znt++rSCzoL37F
hf3pzoal/EgmzHHYH6QaPch4aiSK0PI1vY3J4aTUJxCeACJ+CZSsi3dDzaD09iHh
oClNduGLxYku77av84XCVYN7vqIqfnL15KOCI2bVGcqNB5vP6KlXQFiZVLHoWADD
mEOpkf4PppbcyKD7JsYrsnWof76g4qjP7XUefbB7C7fVsMX7WDKVTNa1X0nyL86M
Cq8miMMXKDAPkEQehysYMCGWtBaSUWAOsPfH94cK0hYCSk4h4ImEXBBWes3tHM5S
Jkw2b+ecQa+yGzW/Atg2j/qOfO9cd+FsOuKmOcKKSd0nqpQ/8jiaXN2/LoudoyPS
/hDnqWT7V/TQTz85j9HcoW7/mWZ2S2TOBR/tuTv5NUQ59h28qqPinWyZ3VFA0/8A
sYPM3M13QFLMp1He4gBK9GEPuOkatYHyOajlu4mlqjSpnCNghbtPQzL9oe+w5FH3
d0imOf/tUx2yVgJ+w/RR7U36BRLdCtPm+tXVYgQG+2OC8oW0Q7hl42LsugFQwdlu
tOh2CuLI61QrQmrNJvg3/b3Q9YnkwFP7BQD4QvdLxTil1oz97W+cYKrjIucU64pV
LinLAgjIMSbtKT9RM/W9x+6c2YT0vOhBCqkSRkpRM2DHWen2bik5Gv/foevsYxLF
kDPy05sUvBL94nDOLBNjS9MyEmLbn+qMsb8ivOi7KBBPubmiQtjC01v9xdR8RbJs
bf9xqIV7YA7WgyvWZswbJGLci4nVmeqxN0d4XV2jfcNtvPAlhF+mQ2Xp4xa7Ukce
7UwPFVk8GTXv8vDCzbJhus2qGZHUSQ0T6iyxCyxsGTrZW0g5pQR+0JDdg3gXMgUJ
FjwzIn6VW3OFzgXCCHU41PVBDve27YETnHhsQtbTQTojhDiZgkzIOGypW3mw/A2/
309lvvZHAOF9IuRgMEHqov0E4dX3ELr4sr9c5jL7/U/SFh1Nvo/l7adql5hnPe97
g/TLHYkIE05TzdcxT2MhXAyNniPQHO5w7VQlfcyF/Sg2Sv1ykACY3i0ALVx+zoJS
jbGX4fWLaLBap9TlN1k1mHKb9INp6n9UFGOOYN6HNAs2+8HC/hHBKq106HCVA1wP
oJzZ349qf2kl3v3KuIiXOmNnqZgJU9LDKNawho1wjuu0ee8hKiJEyCBDKHMO1y+S
+R6C7wyX/AFQmKkP/kERGWSMmwEmz6QuuL6/z2QwYRzU6F7MdsK+yQuxCzDFAF9Q
Hsui6Va7SX7awspFuduINh85BhxgfO1XY9ynRxPo+MC4OWwQ3v/bcxgvkfJAfFQ3
xMDTLk9YRmDtN+qNcjddC2iP2ldGEhgpUDGK1XtcC1qNgpDIUr2PXt1swDuvRZbf
Tn9o9ueew228uRbRTbVSEUZx6zSgITlYprYCdaaN/cbvygsOwSfIZPo2Rjn/+eP7
QAkCAqIZB3wmJAaqs9o/WTZj3c5t+GDdQxsLcvce033heqnnVNUreKMN+ifDicEG
iP0cjAjEXcd4uz38otJpk2IoHjanPteIfmbuNvRTtQRmLH3zmvnYw3WWc7D2rvx3
kgEzuSJIW6iD55ozA7yzQ7ZLT1elKRIBEr/np1f/x9katciUssPEjNGoARtAEbJ3
81XQYm2wCXBm5MtcyDO0zuORn45gNkfgoc3HhBq7RM8jGOOtBJZMM66ilo69l/sR
+90juJWAXE+4aYTWborEjqTjCZDE+ZJmc9cVmakaG8ZobFgnj/DsOGA4g5FMPTRe
vL8oD9lsjFQ7mYRk0pXCKk5czVxDwdYhTiJyb68hV+U7cp12sd0p3wLcMXlal1Ml
A9V1ndW9Wh4/+vi8z9iLrzriVJXdVkwXYh0h43y5cACyuZBP/FstQEPN1Te1vVlx
srPbmmHpqZGja34b3zSbzQ1oL7VZJkcxcAtAYOHnmBcogbtZ4gGDFv2RmEf/26cK
eK4InWHK4HKIAd+/9HDdpZ4gSx3blo48QsufLc+Ww0htUOeEjyqg1C1rxYkcouzf
r/3Qm3mWeemUpxck1KAHFYgqYzoDXOls273acuYowNos5JAK9UifqjPrQXAS0Jet
7qBoKFmSic8+I14u2l6WgnGVzFntL73Bi68asLti8XdBdFicxMeXXZrgHi6KEgdX
lg1Tifk20DXH3Rq72fSbB38XtCG5qvOMC1el0aB3IyFes0FOAIn88EQuPLiaf/zC
z6AYxeJlLO3PgprMjpaoY7uLQraJi6b34iqp544XGrFV/7voEvWFxvNM6OW6a3jR
FQlQOqMTRcBFlJgQBbYOOlpKYwYz3/g8sR1aLkoNPbzuDg/+pd8TjiOV25aRy/za
LZIttfDDunastvj6UkznUWOhCmzfS9GZlclhFofUoJWzJ6xBq/m6zep4qzFGA9Mp
TZxcAUWS32JXqX2VsUpaChzWGVgCFBkZ97IWrf34NweCZJ56qQ2wsvaZILkvOz7I
h4WUSquTjSXvTsj5gK2O8jjMkZusOiHAWx/xhPokH+woTv6UYBDRImvRccWtFRmf
2Frqdc1UFhSru9nS398YIa4HAAwVRrcpp07nj/TiBy6Hj1fGcG27apsPGtyXsADo
+JrK6RQi/nCABHH7ANXcwmWURRIi+sUWqwDHWLRhLTlrfKhXDn8UuUAmENVgIWia
Nwp6tWVQhO2R1AOv8FKrR1aCZP7zQlFt83laqrHfjMXWk9F8pjLk2q+HfJrfJzwr
3fPUVb6BIJ9I2oxYVWb5dGaMJGEFTvjB1w5acsQ8PxICFyQ+WoloQdh/8Idx7c0i
WwxZerD68Mkt7k6z9sy9IX+CuFcn9bKkMVZpLxq1F0NqTaM/OhqTqHBusRh/fz17
UGZ5i8JKLUA+D5IJ9gRUUISe1UWjQMGPb9HH26MQnMusk0sM22q3Kg3AXoz13BJJ
vV5T2d7q4oWKMx4jZ11MjB/jL05+ScWIK2SqAl1vmNJLZFj80ggWiIzQBstDiHa1
BRtHSTXDayCONylo2+Vkn2WF9xPMfguL++zCjcyNlV8f2TjOdyoDJZzTBtm1ENGI
LELfpvB+hCozor0nU8aKWTBompM9R1VAxUFbpogBXxLlkSboVOoIOviw7BkA5i7c
9In+yYsUefEzf6trHLK/KZfcKtR9cujwy5v0Cuc2pdMu6OfTx2WD2eJsOtB6sbW7
8Ioa6PYqIafVNOkQe+p7/GmSLSBFkLfnKghEnynj+OmfTQQg9arsEmFnUDfzl09c
mfWFhzj0dqp91doRORERhemGDIRKLWNGN3VQQwWzc7XnBWT0YhEOobsJsK06K3qV
eGwjcByTwbcizgnuK1Q4/U9ijra2trcMfy2k+bQK4NLTXSkA1z3gKtxm6AU6Ccwu
N7j7hQ8gCwxFN1TJEBzJEVCE8YFFw5ik76432wqgPxccubZJAi4FZ1xuJeouMNL4
NBV0/y5pxAiEycER0VimOTSXxqF0r04QmUSE19r0MT+GbcETYls3DmnrlgqYFz+p
C4yoMUQdfN/vA5r6GRTfgRgzs1VSOlDl/XipHfCDMmD3mW1E+BEY9j0QvxPy0d3+
FyrV+uje+u3ktzQGeMxZL+fTvFD9TzS0FOOXYwfCo971JfkLe/B1qlqNY8VvaUDW
FDNmfqOmrMfmisi87Y7jbT9ty461ZosAiypE56lJXM28ntmNZdS7Ckt6KSBa0nzx
6ZFVD4YKIqP6LsP+vIQT/FN4MWJNyRzmxG6nF0xJYe/oddm/aB9YXxhaRpaEh1xA
1f2bXUF58JUEMiT0DZ3oFowyDSTiolxIlv5MKG47bfT0/zC6/W23OuWCmO+PH4PW
SAmZK/SMNkEna2TVIDpuIYDo+lfHcB/ZXvxcIl3pjkn8K4QqZO588R9xEXiBC1U1
tiz68zO5ogtqW4r7Piy5cRJ/HLPFHVrqe0YgOszccJlaqdt8vFTZ0KBXHvpu11SI
A09V+2gmtkk3ipcgjZa5cTmsp3S6t5l0sX3/Z7dFksbzpzC6SDkqBQUe584xQHwq
fea7ixvHvl90nHzp5rnev/tra5TIlDHC8X3/foSzuls1N8tkG+IOZrMehsxumc6W
YzKDmnurLe1WkLtii3zRC3CN9RZdHT9hLCc2XE0dDl5pvn1fVEU6WIB4lyTW4sFN
tU/GYIpQtCznqdiYhEtqlR4TUVHpLpyl8DblVAckm7h8ohQUkqhvALJKztYc+ZIu
CVLZ13nAWvkpUCEO+M0GKGl/voQq6YYGBVlgLt44u9aLTRn5pgdEjNw/WY8N/+Zy
olCKGyJnH5A7dBI6ArBQfX4OiTlVuDG5yoc0KqcBVzMyTjDBowgxBHShzPqU6Kep
nP2Ib2iV38a6VuoafMS/CuF+6j1iB4b7LMgoqoVaQOZC+zKWiIQ3I3xOqQ3gE5bR
7z98CXPKyOkcUysBtPWF/DEW9GC+3QJXpXOhscfIeNhDqPygJSDNKVVR8T7V39u7
yqVUGRTGtxq06O11apFv/zgC6/G9QO9d5fe+BZbmbDCtW5XSac3010VeWkhr2MSJ
oKiW4Ev2n5cipEpRsfNpmYqrf9u0SWMuq1yx07taokoYfc0/PfgE21BHEOL8w9ci
azBHnSwbS0fu0WULN4HxxqLOV7WUjxsk1+HEjyrchBsj/nuDBrTUhrTdoSmDS8EQ
rHcl6jFL76Ls7ZwcyeqQ9yga9LB/ls1aljeHeTygfxF/HVhL8E8YtnfWiyJosZ6i
iLYMTP+gp540Xnn1ShWI+ZQlQ+Y1VpZ2VMwBihshr5VRS+e82t+NppkJ6JKQuWp6
Iktop4//ZdKm/DyyZ6HmNBllmcIBKGIb3Bt6QyTFQZ8VNyEBaF22i1fCGKyaoy7Z
jUE2ppzX/nBnWaEGQDOBOJvXDgawNU5CRhMj5AtorrDAtl8P+NL5I7mON6y2ZdN/
zCzHOvlzUTO17p6zg2k4/IIOiAAX9bu8KdCt/1/6nYPTs1eEqRcVXwYT1JQM3XrX
Q+BHaCS5St2vfdN6DuyIXGf+Vno+z3D14FKvhq2xBuorn16cnJAtyG2TjO6U3uwX
pCODKD4ETgzMJIbNrpPHJtJvYyGew+jTldkquDQ+xQ2Py2pKpLwtdgcyaj0Uxy/d
TQ0ZJz4cOBdNchwr3AOTaI8Tl+QPAygBlf5PtmA+Yy0RAfsE81S/9C0bi8Mdwhm3
i/8tELl2hEqwEC1Qm2apYgm+Bhgu743c/xRihJWWgSLUyUqzuD7kuCR3CjQonNl7
SqcJ3RMVyfRKdhlJVY+EaWU3SXhfTPUEEwST4Q0KLnaLnApNSUJM9Q+Z/yL6ilz/
WsdAg1MBtk75cuszH18OIiiKIDkV8G3RtLbdKNk1jqUnh/QKuZr98wrdqXKrlNHN
bfBDmu4oXVbWbt9cA9A+vDIR4GWIMiqWqJC/scasB0FNcAoigjNqLnHzsK1hLAKa
5ChC3Q8m2k0BSd3NgFapDg2rBE/PqFAEnRS9UbEISRCWSkgjhItmW2O17OacwzkC
y8AnOPHEUUG2VCU4V39gTGV/YQJhAn7p0+hT6v21FEzI0/5Dtox5LEJRTkTxWG9I
OPGcAqB0g+OmCHmsbxNU8iCChZneuhL9K75f6DPG2J0XpCzrlXRwwl85jcxo/qG1
W16Nx05wMr4MER3kN5/e2zpivSJFf8u4ep8Hu++neTvGkTAChuoTu8GN2CChn46q
xbHAEAFst/uygj1esV6RjriHSbt1ifB0p2HG/CyhfIYHRbNqC4uZbth8uGXSPjgH
vtdZS4vHG1WWmt7khZfCrAEMn86wm+i/XuADm4pFzRWKtMWl12Jfg24ilseRqXHc
kuFtQD1OFGLZgzbOoLUXmuvUX2Gtigqj4D4HaZRJJUnCoInLxskG472i3xxQfOYM
bFgSijAGn9ym+E41EGZ5wQy35t2jwxcAJLOj/Eh1xsfd/04cca3XRpaoOlV09MEb
8lcHcvr3o5XcWsEsk5fBA7qxN5qN6opuA+KtPDETaKAQKv2ktDoEPbN9nShrI0sq
vMgfSFzEJ2tGpT/2tlNlr62pjPkCQN1JMM5gi/jZ3rtQcxoyerp2EByBKFVT+FKy
ZHTfGZUnx44UgaFRU2O+fLCeomsAE9vrkmvtZCXjU4204rqrCllWAmedfdxJro8U
0CGVAdh2WsBoSibh4XVizdJYkZPQDrDt+gprLMYSdu1pL/BsdCxWv6tS3NeEXfVp
MORl5x0i2TfhDETEPDjeVA/gmXl6U9MemZ4NZStnalEJ+29s+CiB7uePrpHtBuW1
NRdjfUHgJbbz7MaOD1A4zw3wURUS7ex2DowvQYgTt7oRgojMrQyNBbIIiZOBKLen
l/YbGtyIWKDTfw0iLmYY7EhzFT//lXI4XKxsOWMiAQyl9sfHffw/YxYAHxbqtzXy
SK4FuvC6i60zzQsC6nLqGASfi78veV5UsVA44CLDIC6lhKxcitdDbQ5o+ydLbmiL
QCaC4wfScbejJtoPmo2gw+kxBUtGBQmYK5+banJLjzQMY1qIWyBwx8w0dhFrYVni
Q3X6uae8nWJ+NghR4sT8/kcoi2xmNVqXJnCb3e1PafUnWPRf1i0Oj0WYiIrous25
UX1Lw2AuVMSaOlSVXrbObtawng41nS8hj1NAwDYk253ioN2Ojw0Ru/VRRWXC97xs
bbfsNIRrUC1cCEXWBIsTwj+eJp1TQVMn+HabNl9+WptE+bwwrOlOcolWmD+oLe+1
/WIJiuqHTvEykwqSktkLCNl0C08uB+Eke0d7lMtMrZKBn01y/2lDvj2Y3Fbx8/B7
QpQ0ujn7kyA0UvHkXN0/Kli5L4IvTDR3IyqEK/DF5YtiOAJ3Xx6NCxj9GPLecVF1
Rwm164AGcytCw1qD+LXfOanPA/MCFqcbqe5mOAgOdNyM9rOYWW+CGE9Jcms4lW91
WBrPZw/uiNU6TPmy1/RnYtFu18S7tXDqdzKZqjKrp5QT89f9dTubZk+bxjkziNph
3qCRC7piBHQPWo/5EdxzvrW+aIkCg9tpiNHdMpf6SMtnpnFK8fDQpckNT1INnnFe
zSXqfdeQohzmKr0/gmp5KCvmmTs3n12y/mtRBK/kONlR4F1Iloi4h83t68dH20iy
HPrL/vUbcdctSYPoXiTuM/amd1f1CEAD1pc0nRkN0hOa4YjJZsYzS3T6IwhRqYb3
J2HpIqfvEv86M3uHqgZ3qzjNXLcNITHykY5muQeXDHermsF/yB0pUv9DtuTy8j7g
TOzBBznBy9emnujZI9PdChoUCSr1wc+BksKBZIrfpkdHhgAZuMSNanVpbgRdi22E
GNdX0h1UngwZeko8QikHsjoRF4OoRTQujrzOuXa8v/aGN/mxmLFauriwoJiGU+F8
cOK5AaXCvuNnmUVU9kZnXCtCridHueIXDT0ani2V1UBKjWojdmGmST97UidrUYeS
+5IH37BRi4ZC1dnxK9xf4BYlch0nJEuEw6Bbcg2KskkkaKQ1NkPouAJvRjNhttXw
hn9q4mcLdEftBuShkXHuOk3yEIqGXCRJpfyh8c/4Hx9QoZwDjbsVaQ0MYNumJQ8n
HCxnz7U81lWevui6WMddcc0RxmrosHhOB+dj+/Sp91e3bXL+71QzOnZzB+27dDcb
cTyqMtZaTwHLIoweC1PF8Vhr9DUQuy8Y4hmCmVpqO4PUjghypdPvip0IGh3emn86
Yhj8qm2bq98x3cD0CNN5uKZR/ZmrgVogfk8xBLqJZpWy9NfABN0EOsXpmywHrmKB
B2eXfp0M1OqSDue0YndMrruAWsAyPyZvPgbWmT3Y8w81hZpOry7bJm6fB2QDQtHg
hLIleOqn4oCmbEI39rf1k3Xx8WsPI+Y96x+zno4jYz12Jng196H5dJ57vuRNU1fx
SRK8ZqJzd7W+hcXmnlor1iWXdJQGOJ7vZA+ToQBCF9jI5XpNjd3Mfoy7Iln0kId2
KLMe4rmXZWc2DYO857Jr4sTs+uvLwf5KaR3AACUv9zNxZ/WQOEqojiyWKSwjXvYu
M+D/xD91GT0cLVvFnLnQ43YphTB6DvvU9tDqHO1M0qs080tKHYiVRXRiprTep6wf
9siCz18qFH71+fClAPf6688ulDwo3hklpesqikZdOQgSJrrncwr8cVgewi53QWlC
UnLtGKG3iBrlsPdTIFCdyexPNCKEi2KNfDqRbSOi1FhkwC5ZPmiLiSEcggA6pu6k
AHYu0wUEqxYXY1JCuSfNiNhYDo15nCMqzFN0/M7ucs6ADyhIm74tRN0dnC8FvZ83
s/PdJChDsVfCAxi/FuAtf4CWnYabXsEp0JrzRm9OrrTuYq0BMutBh0NDKsmNZx+C
bdN8S1bzuPae+nYoC6v6psgUF9ayiMN7dCoYOaJe7pnSIp+Y4Ztt/UlSgxYtTOFz
m7ZADz4lD2Kffws3s0kRB49F3cZEm+D+p++f+dnFDne5aDOkauPZhCJRAMJjwnMq
YhjotQy6KjV/kRHaG0uHMLZrTjn4T83qOn4R74gLpTJyhQGBisDJQylwCLNfmaYm
9Glc1S3bNajUhNFR4PVdM7ifcwJ6VDmdiqv6i/kgmAn3r2LCohrz7UAItN8ZlyGh
K58eLQVNg+NPUb8Ft9gQRbdwTCjc2k0Uaa5j+B9f0pdZMclvtU2HtQGwQI3jhoVq
OI5I3dj4YmAHTUNplARItNUtazCuj/scPVqwQ3YPwhixoMTY+u0z2dD4AdZ8o1le
xuYT1MvzuAPdJTlvnFcIV7ADKOENIeLKzV9dhTjIPt5IO7yXEEv2HWG5vIJ+sgNG
Ws9tQu1O5g8eBxSGaM1D2uDeYxu7ZjEMgFVcgyGh+g6rlfY4VD4FpqwWHGT+SMFy
ylgffFybSES2WqwuBqhH3U1cizJgzezYbp/K4ZrC3fNSQonQUcSpalQaeBUo/8E2
m2D0wyqzzH5ZYADnWZmAa6I/noATj3i/2mE3Ljx8d2hCRBcSLn/lTOX4+GKzFzEq
Y3xQjyC0kRysVtLt0Xc0o7A79CUl+tl0iZR4VhgzQhRvuwH4cMSxhpQq7Ddw3wmX
TIgPORRoQZlsuvCXXmKYDRZdvVfRZ9ggWvRXZVHP5vjqSkk8EPY4WFIc76aNvqg5
tjzCqJuxbo5X11sryKF8Xt5VgXk5L5f3OKIztybmMdZK99BiKR8JICYCUUP2wPyF
jxfMC7ujjKbiKSOEHHGYVqElPWJ+vFJbpg6r4eQQUrljwFyq+deeJKqxbWHtlf4c
arA8Ip5FQYY8mauXRx2fwovSnH/SUeNXIQnvNj/Femh+gBY4zIIiB306HNPcn9db
8UykU/wleLZZUD3bY6lZ8TPuPXTLgPfhpZtomtNjqxLv/vHAfDebOe0Rw0MImTlv
LXJORi7NsG0ahTgsMvwh6gupo20nxhqjdj9RcPUmS3HZHLU0zmkB5CZqf898ymN0
xKdn/VuKmzWXBhqsZlv18jc+Ko2l6gd4hkmfDh/G+glDzWzdhgNbQGoZK+9VkEq0
ZHoDrlFpZHM7q5SuitPzXRpNDXL+mWcK74AmlhKSqjUCSO22jaIp4AWXsSq76T23
PIsuYK3RsGxcT4lvUQPKTC6AFsqJZuDZ/ODt6tVOUhzyQpg1C83a9L2BZTmHOOte
eUo2Ss1jKmi+bO0G/hvd3POEt4atqevJQgHhKYoyH8lfMSQpKvm3/W1TexatFkDh
pNz8teGJS0ybUTb3NHqTGYpJPnucL+yMuZmZImykpoCnBG8QndEs0Vm361G/frh6
8wNdjsv8AZ7ZzQ/SE4wv0PpU/JzxNdPWeSoVandNLOz4jVdAENmPrMs6CGgQeD7f
vncNi2lWlyoes8tdWVQPl21YvryT9bGARv3HkHeF7cYOPF7N51ucsHk528LE3G+x
M2oR8FbAcpFvYSXexAT6sj4n9cD482ae+gRhFzaP3HzUqOIQ3dL/vucRUctIxD5K
AgM8ocKHxPtjS61A2S90EuD9Q1ejnTB3Fwlr2cSXtGKdDZsnitcsBMl2+U8z7utC
1dALk2lrjuiCzDZmtjaDktMahKp1e/px6NdqEBEYc0J/q0kkKYox8MLfKvCf/LVb
DuaAZ0vpVuZmqJM8sxWXHZ3viLd6yTQ+aeHwdEDQijSy34361j1rWtLuDbH8431N
KeGSaNCAl1hrK7xrFmOwLR6wDfl1WafmT+BZ8hMbdXFDtRWeCaTdPDrBXKjxNBBY
rCyczMm+YqruSDbyfd/9sl9pEQKJFl50C1zOuxZAKpdLfy2qW4MzyE48Id1svy5u
Wpga4lfRMsJpvu1oDzghA4GUfwRjeoLkhdk3mWfx+f8eGyw8TmGjP3mu3Uua40ee
spJ1ZYPyIa2SCZHHi945xasbvv40/erpxBXvxecMCoJBvieZDkAbPIPt9JYt63BS
eZT/y/0Uf7oqT9LHYndMRoIUdTwDy6U/BTCJf1D7ZWnmAntpqK8yKisZMBqEJcUn
zBUkNigh/twQ/alaNwc46P7onrBoLkWYFupnAZceo8zPi0+mtJ2fhu7N8JhYL+Y7
kmzUiBzUCuKKrfqKfv094/T3DxF43gLwPFZ9jkVn2USy4bKOY3/UaHpWKHAkC9qL
1aCOsoyDqr+dl0i8ujDWgKoNasojS79+Y8/j6/gCaRUPPBEZAKSC9ERcCQSrbp2r
XOpb+raDIzDJ4TeQHEb1WrrJguDlBGbcrtwzeXAekg9n2fWni57m3lPlephojZ9C
fV1k8ofc8ziYxSUKetCPzWhPPpf4YiufqoQmrpuq9G/HXjcbRUmQdliKvzzhpaIL
Mkt6e6KCjh2VetkL5F5A6MYhi4eN+7CTWKPYwmY6UxQGCDtAxKTsESDrNU0o/Y9q
GdOedOFOJ9MeOKaV8zmJXOH816W6NavVe9PxzzxW9IsS3Lv+qxgLppfKJEz08CvH
lNBnfUk2By0S66l0xxKlyutps61xrxRARLYYceLmrsimastuMF4s4BHFcVa3utOE
ByrpU2//Jd5t0SGOdNuSATU+OFECdMPXgxrmTwqgM4gflELI2gLNRNGxaW+r/D9I
0ViHNO5vix098dWiwFi+IwC+lCfHN+BxHwXGuaAkFUa+0uH4zHGbuhvuOB6qWZx5
z+tX+eYV0nbKpfReG0B1muCTtgvDMvCp+u1sHjznkjjboVYIR0lNnZcLCWEIlYBZ
ijxXgslmuhgfTwO4DGC4RhRd/3wtQGWEOYUtTp0hrnmf/bJ2cdgfpqPerN1gwU1p
FWOkRsnOrxNzDzCDwW/2Jw3BQJu0C02oxL2UdMx1GU3a60zcXtFrRRieOxB6yAXV
rR/NwNJZL5dsYGxaKdNBYQCEaxE/wDcx78rqh2Od0Ts0bxQ4bo5BnXN8HEutdvbH
xgGFCu62vUu/JshvoboUeim93vRaH2eI7j6B5Uc998N51V+Ec6WFTTVSuWUJQzfE
N2Y3CfgAzogYi3UydCobJtkBkhgmIBb3lNI5Q4JQPKuWwNf+QKPb8qeb7bDCefPP
9eCaWdAUStbaWRuQ+8lBt4nlmebT8mNMDqi3HZ7MEJzmaoa/h+Uo10CWtwqI7hIg
zKM9ZFTKwc+mBV3aiZs73ek7+bEIJ0z1Gvqnec4wVAQABMF8mY3AWNKCg9RPHy3f
kb2KgFQMWlFhlQ1lCNxPe4shdyqa4Ne6i/XIEZAYUkJGfewhciy5/EZ96ZDHOeJT
0r7X+f+fvQ6JsGlGjmo0nH/F9WuF2Punvmm3A9I+zx/yFmWAJtg5z8Uqs2jyiKPH
FhI5mc3GtUEEdhAEvrl7kr94GsI3ttXgcmOIagQJZna+98JGqJxPo4Di/Jef/KeT
+KVWCHnmSQ9mEqdsfKUAopROy+e1ADvBJFMJh097CBcnpo7YcKF8PTgcxJFtSTgy
0GSuGy209iYtU5/vDhhLsvzeMARzUWS3P+r5GgBJD4NSozJq5uwG6zwXP3XW8XkL
RvrlWF+QZH5GwBKUQmYZ6jjge7b6Be1lJPZx37gTgc0jEu1qBth/HOM+3IWCBOH2
avq8JVKwAoXu6+Uj448REdRAHOwQHBwTZMmqYzsQqneK7mJs1Bg+klj7Zd5QsMvv
IlKlwYqblK+DEnJeAvKKRQojXsE6Y3s0Yu38IMrFVctHNhVE8hBMf8kSh9buyByk
KmyrRq4u+A8bsU6roZIiM7oZ3bzDeT6FGuSR8DFFM1LFyMeCL6MbyEAyxxNnqnEU
aL7GihVZ3gInoTBmGpGdqzH/gU8GU7ZC8v6rJsFnctPp4Cq7NwOdIgIwmuDYD5eL
w+e+jhhGdcVquQ7otyy5ixXr0SjVYBCV4oU0QTfvwS9enl9tNCheiDwPo47qs0tQ
vP4Z6UB1xTnsWn5SWuwvPimoFdkkbl54Z/zxhMvd2+Pa9mpMDisKmWDE8Oh+3CZ2
sMlySe1JdJKpLXUYewyJajAnVptROiufxmskexGDVMTNCVRK9RAWqf6YJsjksHns
0F/QEqOwuS2FQ8YTJIwOXChGlogFFb9e05U3v0SkCYPPrumL3mWCdy3Uu59FgHU5
/ej/evtbtPqT7dIZlEUg7tt99eRZ/ACCsrI3xdMJ24nSvULyqiRxXtx7eBBfV6HJ
fM5aWGUjQRKG6mfxI+sb1L6p50LVl7E9CKH3458Ta7AILHpWRqKjApSDiFwtM0si
JdvuojBlNSHQkQlHdglvwc7A+n/oDJlJ8bd2zYiGmnCaiZC0DISRKls9tTI91XaI
ak5KN1GOjTl3F4hFV1uQRkSWpilfgRHqDv6weOhlkbiNMxWUhqXzYQjbs1K/FcGi
/dhjpl0WEdNMq8ko17dJ7t+zx4Ts4DVFP3rkFesxO8NxRp8VslGLtII5qqT2ibRT
wrRpZSQDS8G18fZFGbdnkki8i+W4S+FbjXB52fpB8mB/nvJF2/9dZ6zXSqzAhTtt
8t+E0wIKynyIolR1rfNxTF9BkVkLT9MdfcSxmmqgcI9a1pec2OERbzCutcdBqMV3
lQ/EQqJZNkgprC5+i6qnzFgspxG7ZzwDCjjsEuV7OmBhyFPuQmw5w8ISwuP7nWKt
`protect END_PROTECTED
