`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R1BUtaaWxxUWjacRF+bVeyHkzqWqzFOJSLl15pFmMSPWceIpwE86lIxkY2Ieb75l
lkFS1mtI21gtf1ujiOrRrGfcKDBB6KoJ3RgNpk9qbEMpvlt+waCVaGytUiS2ull8
b23sbKGWCXW76jtGUDIKGxcNyscanlLpU8HcrwPi2CPtQJOL1E4waDwy7Ep0ajUa
XYcUpmkkDQkzYZoBXgekK2At5OJY9ynbF/bT3iUCoOBBHAyYtXEYojh5MTbhWPwl
JN6bhjGFQo7I889W+bzoFlqrdTb+7XEKnx1MwP0WeSlyUByCM87FCezz1cz/yB2J
Pxl1yvVqRtV0NM0FZU/g+mbhwxVOkIihodP30ex4MgSslsY7DTsGElY2R+CKcnh2
AlYRog6IGXayxd6im+5Fph2vAb9MKXbBRYyVPYbFVJhGcN9Al18cZwze3vJGPXGK
nFGY2tfK3hcsi/2l3mrqO+TYxXPm/FXUGwbhe1SqbYuKaYqca0OoOVNID0QrQ343
PWXn2396bwgWLKzgrVQc45xUUMWuv9RQLIxcR2RJjdY2TjlDIJgLBw69AbuVMYLu
SExydek3YVig6BKlMIutgJxJLo5AkAX9eY98uXSLikH7zmtpc/RNaafa+NQwsoEy
wpnWix8Dd5RHoXOf+/SXtsrlZI6at8XXCKTeigCseAXLsIpHXToBVhBqtCEGBRi/
1SL1Msh5nG3g3RChCJ/gC1GVX6gzu7y7HjyGHzinq2PMQ2sPHbScefiV2WErMYBe
xEzBQevrmVXIvhLodXzgZqcMMRihMmOpvCOAKIF/IgoczhMl1rQuTO9PGnW8vqS1
HfwkI46qAJA9UgcaO2J7Ubt8WQvTCBSRwdhkIJ3eSYpc3BsJxjDqYzyQxJ92dJu4
NDYlKgWR8U8gCjKi281kVUYrYJn6IycewvLtPZvXE3ydgrfFpyDsnhNajESat5N7
77/hnBGNOeUFB59JyixkbwsExVDuDycFEIh+qj7l2FViClcN5zE8j3gOaOuJE65P
3qnlJJIHpX2CdO6imHGYxprIzMQHeaJEjtBbEww6wshe4lfCRZDBARzQ5xEJSPpy
RM7PciI5B67wfp5bqFAUVKhGSwH4vkf+hldMHugSGWYvaomfTuVEc7PPwwO1/kdo
vx3NCsnW47aOqxxkLY86swiinN3Pp49MDFyPMEXIaLXW47geO9gi7M3Fkp2MwtCs
gZ+GgNPn7OYhplGmh7VYGnI46Zc0O0Jtr3UXpbTRd56KDnbGJbgZK1m2C6m0wV1g
`protect END_PROTECTED
