`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AnR4QswWHiFzxPHD6Soi7qtGX3tQP7VDB4OpOztHl5cRxWOfnMtezWW9zR0YSd01
5ImchDFixN20wyyeN/xVycyA2FTj/Uo6rNzW8ixuch6GKwaSfDq8TX+S5+nISBwY
gIQeVvPsRjfsH0YAtAlteG7cjBTuK7q/GoSSY697qhYfR8ypu8oBWa10hCQITgyr
xlUGLDGo9Fk29kvzMEguga3Y8Ld1gLsA8F9XvRIYqALZsMM3hl8aY5o3Pyk8T7O/
Bv51AivSJTkAY9Tq/sypC5QA6pYQddlPpfjb20BAj4QKgtzsQ3D9Gvr/uV/3Ld3/
aP9NKfAsrdJWlXYQzRqkep72tp1IA8jFzCgubuDHskG8ffXFXxWG+QQGH1A3Surg
TrtIxuZeEcQaOCDouzW1zS6e/aioeSclR7wsj3BAHi1qrTO00v1Rj0c3UXCWQJNN
E/lttxnY+lm/63ojJr0QCr6eJkZB0lx5n6cp3dva644donLa5m+PdByIQ6ro/fyL
LdUlryQbD5YhmBSksm1ApyxHriI7Qh/omxECZ4w9y7GzRDDIm2ObPX2XwJq0dbBO
O2FTsb0oVpI+Ta6KCf/heMj9pBgdeC17+C6wnHKiJQDFr57zM4DMLlrJAetMO6yu
u/TWnvsGdGqbLccyIoDiZz/4wdQ3CKEMX3zuH94zymAASeVF3DvLrRn1Khi4nCmz
N4lmr4rcS5VVGNDx9v8XYayBNddyXYKgsNMHp7RfC4ygNdAUilPncB7VBgpiD+Kx
/61RpH8b7N/iZCcsqTJSRyKyLL9TQD97eWqFNgCNFPCWiM5feTvis4k+EAw9JUeW
FUams/8JXZaoVhLr5+XJcgV2yL2nYO3gonl/zksB1Wo=
`protect END_PROTECTED
