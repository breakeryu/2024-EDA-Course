`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bHyThLqLsD/jZokImQzVRUN0VuCwRt+IhZLqoPYARKEP2+Pao7Er2Gs3b4i3btm
b2RfjuIXKhOEpTkuMgWRQjyhBaPn5syO5MjhgACTOC1UBjvvdKSZK/PGVklO/uvK
8YOdiyIqxu02vOx3fqdEPDf2O9xB9olhmgqJHbcJ0CCNcPwaVyDJRZNiPHrPmG1g
Psaz1s1ONwuT8BfkqAw6TZEWGxsNZE5NFIa0qoRqeWqWFpJrLPh2OG+aFmShKymq
oXpA7fLFG6Z9DWC//1Xl70tXbdydWUXF2qZdyG34nnlYwzCOJGsbi0WqhsQSlhY8
w9xHFI1eK4lPf3rW3gtQ+kSzyAbTQ7pPJOsk7GZ5XhkPTjn4sQ9xIXCTfinWzaWD
cka9ftmMz5jjMfJndNXNuJfDHrc+doPmX3pKkIdxB4fiBHEUNrInH4AZQ15cb/qL
0LNkOpF7WHb0oC15FYdKpbnWOHR51c3gM4nsbY7wxLuZa2kNPtUk6Ud6hiRHaxwt
KRY76cPilwnQH/smYBGCQEGVgV9nJ5UjWNCF1XIB0CRfuLSmtGhasluV9F0NdS68
I2Dbx2EtYKl/qd0LbM30A4/9e/J3braabCDCJ0dwraaFzTDA3xInMIcRNNf3GlLV
f+gYzvl3TzKu7r+iMa+5z/ctrwDWfgMiJ+kJzs2/qMNcu8eGW2ifGAJQ6cWMAemG
iT1VLfRmYI42+nzB4Fc1a0+2AyBzi4eCYHtIexJKAFneaBETwfo0HPuiem68XZU9
npBmkqBKteMaZiIofMrQuJU49BjrdV8Vuu6caRasX2LewykAkf8PDsjDnSQTGR+X
U4heS5slnBPh+kAM3noYDZQufg2+CXo3rnD7/rffyuYdovIFlqnGmA3V7dd1Gdef
AuZ/xlquhc9ToJuvxCMwldQ4S7jEecP/e2L+IY4XiSA82MEMhyMwxjrzF5E/XLKL
bCeOBUL91bcdJP4GfOTQct9cQH3s8ElYaONya3T1al0W9Jc9ujXJGBjWZ7aoW2Yd
JzbXO4kxf62P5+Bfl48TvYvDK5V6M6J6TbXZXzy1AawnIKp0MWjHqLn3UZmbbk+o
d8Chokqbnewfivk0ZmUnl78sHd0pJT0mnM7NDCIc8srMjzexokBLy0INEhkK5HHQ
yqXr4qDfzB3uTKoaxKJlMw6uRc0nJ8+r+LBaoiOE90BOZKt5CR+8W2G/rcxLHeJq
E2Ymwl2xxWHDcu3UEhegfr2wiPNRRIaCh+i8GwOE2rcUml+YB5nWA79OAGlakqdi
FRMJBLKD+2zYnn1v4XES7ZhanJI4sbLWJV6yqZtoOf7lnD5Fvp8v8XMTxYKJ4mQr
ugGtpp8jyiAwU++1N9kaokuJuumDxRyNbDDms8wj9vhIqYFsIoPH+tDQJB/oea0X
zYOimq0UpkScXkfKCqOG7REEMltuMJM5MbA/oxN8hAkCHOxfKpRhJvsQ3TVxSEtu
+dE4v3ZXQp1n9GbRGSRuwR5N4hYYCt+8oS5OOlEm7yxmMxxOlx8xxMBOgyAfdXGo
ZOx2Q/HSDGN0uBQMXgWgYGWLK3M39oZi/Apw8DonWMWknyw4G9IYn9z2p22HabqM
7Q5oI6AAdFHjEkGHAIECbff0NUWmfmCZWLTVhAdTWKRN7Gcze0Abht+aR1aUg91t
KagsYZRxrCdinJYSvwdY9Tv5c/33rrEt908t2a0ybMJp7iCeCh8eD2suoJgI8O8x
uHSDJVlhvXecjfFZm9oZ3YGxLjsPpekgbol5XbgezBlOJ+vpKV+JBIANx3zKe9yr
QNe6XiKwtM3c5oP85lTJz2AbdDOsmxV6++nooV1kcwMwf6sTnrI/Q328Hv7KZd+N
+vFV1dBjmRiSNmI4dbE7cdzLhON8MeUfsu+ndWpO2kfTFoMhIlvb4YXKB8Kbq2AT
fHJyL1K8xP3GbLZQ+RBk5A6Kr/EOhGYxQAvQCU7gJBBjQ1m+fBfZgFpB1xE7d0XO
u87gUamkMSk8vjH9k2jvsaCg9ASGpuB0lbRWVxAanPxGpTpnPPjqugGYbUva3rFJ
k+OM4bmJJBX2aWvYpaEysKE0xkH86AtGm9Enn8DF7s106IxSV1vuVVWlLC7ssZU6
9HBzjPRXXs8PY4BhVs0OENWvzeFX2X7SKvnI5Usflt6BiuUCkINlJ39XPihpCxID
EPgcFYIZgshroiAF0ld2uQmhB8/irUzDHd5cshxBYujIkUa7lA4wdviVr7vfVFFd
4k7K3E6cj2UWIrdHA6QQ5NjnqdtDcpHNuPxqg2KOq8AKZL9k7xO8UDg2l0/nuAqA
O0QjFZdY+lGsYOzaK/4C+c2R9AFGAvC7yyOsZUab3qGJzAymAK7TBw0MGT+7bNoh
8t0Qq5pakMFPcNqO+9UYWUHY05E3RTTlLIxlzHeuv5jMnn+J/Y+nPt5ZEzjKxC0A
PnW34BFQ6glkyjC9ZkLRXv1kHjYMSu74b9nTuGA8udzbG0ddQTuPeVbEdBvFi3YJ
DH5Dz+ZaCOdOr3pMuRrFnYg+7GB3Z7XfCGUNgPP1INbqKOVrw7fXAV0+P1THR/Ue
Kz1IcD3uc8ojMeU0RREZjj7EGrU3iikYlUieTCJbgJ58HdAbYUwvL4JQTNzDEsTJ
R/g9T1jx1k2InDRlojfUESR+TGEkZD+l1Gu5xh/fcM4mTIMIPHYzHlEA5W35pecP
MLjfqRUVE38Pe4ad8S7DKlG0E6EtchPMDbZ/NWUrre97IBGQIvOEmYaJGq45BJ4m
2lQ3ATAHX+/1WufSE4180f/7O/i14rlwYZqdwof4kqDIxbQmLjUo9vcThyXhMoxj
2LwHcTAScRoqqWDsVB3e6yS/0qXRlYVaC3USCc6uXy/cJ1TP04ZOWjG1AsJuB7GJ
R4kpqcSSxHJWgKcYUXwCfA0G4NDmzVbPdYKsOF2ogO2VICaOX3ktZjrtx9HLBQF3
IVKIFM1WIMRY9RbROs+VVlvhK+OvR3wm2OOQsrfp20FkYrIUduNQrQrEJbG19ie+
jz21Ptj+39pNPs04Mcy65pFJixdO9fPLLH7AyA5+lnUu8+ET1QeuM4RywVbF29NK
8Ws2o7im6Xf0rrHNvLNZHBlA5iDuea8+iQxG1XqMC4LcX35LiIQzeGdQFx1y3Ajl
SOW4iUiYHQoASFhswXsMy9Z/R8YvkhJyPrZXQ8QGlfpcM7m2GO30tb2qsR8cb5RQ
1Qacj7fq+txqG2uw1AfzDdy5i74sIp4ymHr3jaq0WuPkxHK4D9vAwvBjge8BTk8a
k9bWbL9gP4zs/FiMNBvN+G5+7/6wJN6ZIHFB+S3pruV1F/0pv30Z85r8o56xy+P2
UjpE2Y9QlJhFwXSEGs7K4DsoECHwHmBUFrCx4kKnyohpleXDdhP9gf5aZWlD0kp/
5pkvqlBz9xcNZC0FWK36T2PAw7LjBVN7UIeCHBIh6ZLSABHmwJmaZpFaj9GyZS/M
8lcrWBDWCdi5Xv49kO24F6ytIEr9Hfsta0ovpov0NJOvedhRrQ3g6f76bGGOjbzj
eCqbN91u9OAoU7i5+RZdQzvHNHg7geNGWa98eFO8H5661j146E6JvJ8QY4ac8oJs
/C+rkaMdySxIXq7JwWWWATNCyOaAOBNLMgvUuowXlxszR8KgkL9qI8u4QuzzJpUZ
CjhLvpK0nBx1W8U8w73o7ZJke3EFDmCofr1wQrDQ6tqwO+mMWAX2R36BMg5d0nTT
g7ukRzcledOzo07Hif1cBePKqIBVe+UPD1yg4sIak0DnvPHMWSl6QlphDPMFB1jM
7gnYXvZ+JlGmfAKiUJJSHTACwTwvqZgiHjQPohfDZ9PY3OBSayAEgxjCi/IXm3Pa
cDLkNnCb42+22x5jbcfjsgJvmR+6N1irIOK8GO6sOHcRyYuXPmmbb+vrmSn5m2US
Jxz/v+FEb/C1B4j4SL8gqBlriH7WHHKV98IPZldQQNOY58s0FfHrGWr1WUapauZ4
zgRsBJXJcBAaj+b8/+H9LLJ+NOJb6WiViev7eyiLtgFNUtoTSrglR4cjTdQka5NK
4vGVvYWAdN4HBtyFJhsbbTgrJvAu4DB1WuIlXGCvhT8T8tF7TRTHbmXOmSFgfBqk
vPd7NPsQEMu2kP6MlT0VYuSOtr8S5hy1g/ifqjlBrNB6+UTYMdq9LTjOCAqWl5TN
Ih5XvclvBpMhaN5yHGl0tl5w8vBqM8HYt2mvWlbh0xLvd5drm/O+YIzPUlj5d55e
epFQf+NJf378jQzSIMGNjzs9pyxfa8bQNTGZK5f9vYcn0Jxyq4BXJn6bJSqOmmFH
IrR0pGY3Bq9EAqWQAB0DTVg2IruQuOi3atDYIQRkoXx42UGnSi9NDjtO27W0QJQ2
ft4u9yRrNu0rXoTaegJpw29ELA0tCOXv4gK+/ZlRPi9IhhY/YRaLKBRY67tXISWL
jFhVc+a1frQwd/VCURlma1t2JUuSMetbbHD7y1b9AnNzMYre35JosF+IOcdYiTrQ
9Nxn+WWoAtEW0IOdMGO2+o2dYR/PajJmRSI3uelqfp523Wt+V6QiUjASkLD+M7Xk
gRz3GgONDyCQzYrAltKb5ml8yooQoQPg0zoz+flF1Am1nEjezLCufSVYWPhPLt/G
Yq89NwcbXGhKcemnRLqEi1FwlkgJpwbVX5bg0Wl2EMcB4f+4yUhHSSheX6TjG3Zd
FdT1tfeC4hWIvWTCgrOzNizAHL+qtIH/kiWg4r3cNyvdDhvkKz0CndwDFSnEt6MW
c8KxM0o1ZGyNilue80slFn3/ov8alacK+wLrTdoL5z2VTg72aAu4HQBPr+NlH6YW
zAcjUsfMH3NkQbwRDMCheFg2ps4RAcCD5ozzsJ8vMplnDESe2d0TXuuhi/ECSGLI
U2HdVKYrBkjfoWIwyxSYepa0DIsLFed3U475HgsMj5qet0xuzpe+sDfftOeqNXIT
BOKVjFLMbkrO0uvTMSUH0pYfQhtrnsqPMKihHKUB//XiJv+OPR9I0hvjGwrKpW9n
3khwpNx4SUrTZ1Gr9b1hYx77s4u9GimEy5ajTjIKr4+K9kLox4C3hX+/3ZEtFt94
vg5/xBrmOS+Epb+dNO8NgcUxEKiWuW5jPsZIIHb+/f9KD+o7DRLqtgw16qmEYgI1
pcXuT38KHLgYwGvLyf7nOK8yleanYEUMUGbnl2rzXh7e5b/My4OCDLSiK8B4lL5/
SnfVl2uCUQHuWrHExf8IKhEuImzauGPdm/yADhjgij4Zeog/8lWWEWzJzZYJxE1K
bBMf/m/slsb8PWyHep0QNvJS3eqFamDI9ZTVgiS2Gct1vy7QttfuWLZVIsP3+1pn
zE4cb4Jhn4ocQtsj4dah+ovvaxNluba2t9fATXOQ6hoXLf7oKnXjOw8y6TOB1gPZ
BfN4O/oAjQKH4cIBWCnDtbqnmCeLjgsEqqQaVqSN+rNTVIaN8/4Dc7erAhKzsWa7
W6CX6fWkv0l7H6f7X8oiQSDMxs8jHTUzUVtjsylPjWshzw0FP5j2c+YTDuQheUbQ
lgnfsThe6q3hzgJWoRNV+MIbyz2b9qt/eo1+wjm71x8HvayH/PDcwn0TrLb8xYLk
9regMyCvraLscN/YsqSVGRuOs+xX6n2psHdz+93rFfOEUeDOmQQY9OA2RCpvfsdS
ILJAU8drFOtRudeAoydRs6TQl6Yj+NLtsFeTTXSCESSwSwoo7a3l7prywsdoUq4q
8ozFEHdqGwsxTp/zsEEQWw56pK5HTk5YwVnIy5zh58WIPHFd0xjo814pvZFjKX0E
KQo3uKuqSaM/wEABMuUSWkIoJUyD455O1NYlOpxzCmNxEVpmfeOhCBPFk3EBpVuD
SU7PZRY///zV+iEcNU3O6z3+DXFC23/nocu7QYi9FBqNSVYp6/SmsPt3B+sgtDc2
3HKVrQ7IsJUElEliaet7dcZRnoSpI4CzVPkf7TT2NUI/YqvJRvy/qrVk/Zk4SGGj
C4VChUQTUvWk2Avtr30rA7aENfscABWgs7t/3fnwTvImvv5FTlq7CxsltWvHTLxV
8M1GEVOT4GnooozmpYIateB/3xWyNIGimqNXv7fIBeCY+fxVMaovPhk7mQPwjuWO
2HGPq/xhu38ape/0/Vyai4LDNwKNocle4l/7zio/ImCYzp1vAUJ22lNMB1qmKEdX
qw6ajUEYxRUS1zq76LNuwZ9ovU7O3yngEW4Ix6L+JYdyQW6WMFUtF7h0uCJWxUPu
P/emWpZZkCnBqazHiClDpQ0sQJRoQU0O9+XyRNVQflbBO7p6sS9azvsNfv2e3AvS
nKNv5vXmDkd0Qp0E6ucd1EdazaBvbR+3JGNoSyETcPuAkiPeKFz17On0cVruwvRI
Amo1x1Ko0IZSrgta9MrEAWFdW3xP+//9T0ugKFD0upgiv7cRCUyGQmyYxRW5x2tK
v1tQ3xYXzdzVlklc34qQsVumiKieFgKLgQ1XN0M6TaP8Jo4RKjljpsBP971F4E6I
EHZLKQzbvkW5dvJYxplhLpoabT5W39Tny9Ge//iqWV9l9jOr+e6zDdJFVduiqNEh
Uod2nU5oaXnSZMRDHKMpmeiGDVFgmxB9/FgAiUd2qUaOUxInNUWjAAvpVUlQTSpv
RY29X0BwhWSoPIygyKdzDpqakDbJty0Sf2KE2JqAObfw2C+SLc4OZX228P4mweX6
KcUXYQwS70LV/fE1r1gKNJwicPKw+jpeVad+PykqzFfgtw7Ay1hnbeM41mmQ+Dw+
A6nqdZKeTPIpRsjklJo7Cnbqw0x6W5G+G6IHJ8Kl+G+sEmHu7r634754SCsuf909
gCPURgwCX5D562NdiAIPuy/y6/SiQbAhYOeDq0DzJJJGGEIQcGynWKEw63sWUCAG
0AluZDHBrjx8ydC8UyA+8133Kd/a+sgswiM5OuqOae+CaLMPPhYhFtCp/40wOyZ5
ArOyJiNOAqFgSDcyIqlJST3+mUYAu+APwZoYGfKoX5UG84Btf3hSieUiZq4I3pag
D+AMCJBXS5GPyYw04G9yxmVzC6WDMicSbwPHGCsoMi9A1gqSaW5aTa+tMUYf52CW
3Vb7gwVfwTi1VlhbP2woqFuLKnDKx51HTC04DLSOy2BTPJiES1hlMxFdWlN5me1l
cWWRzb2fNNBjBhPM4M3zjJX/LWx54fFAkOo9kz5XQhuFsaOP+3xc9iGCAXWxjPNP
B7fZ/FNM81GIGf789nCUCk/jrd1uD31I+uJ9Nv7GRblKSsV0NEi7fBYU4m9Y+m+C
yv/fk4t5SAUflaeUQ1+Yvbc1Ww9LAWIe7pD7vZj7H2WgEJ1RrPYHTMVpIJJSiczl
YYReK1wiV8opUEjty9Vx+pfuluWB0GeH1M1eynjCz3u+/m16uzQQuBblR0IiSKmF
oFU2fL4yM7qSVFzt715uxcXF8EgkfSfUYVNwrEcNhNuZsOrKPmqlhXHL3WBOV/6O
tQ8dyfffpJcWGneuH7fopl/b4HlZlNUCF6gMYnVnSLX7xiYZTdPKz141st0Cm6Hu
Nh+r/TnC4qEJXeq9+rWt9F9WpoZZtrxxArJo4euAZoFQyUF94KqIiZcDDGo4McE2
kgVDBBmxoPkKeH2Qbigri7UNSz9TjgV4e36Y1ycatZrBSjZPMYWVdOGiQt8DE1zj
dYtLjQvVrWIp3n//aWn7QeMHU6UKNoDp6Uy0O9sxJwV2c5dWjlgTiVPUIqY98um/
1OYMEnnFhtLjMCA6PVKMG427eWtWin7H1151dIMz2VmeVSm841qcVyiwOsPeu9ka
sPFFTII+GotivxClLySIybr8tboprbelv6eNMkMBKkuhsOLqkX7ghp4RRXnL9GhL
LH1fF7QpO6LY951xgDPOWes/cD+8ODI9ZBfu38SQVx308Gj2OTjFRERmEu08VWvD
WBVQYLuDc2oxHaw0nals6q6bw7o6W/kENrbTFq239cefjxS/+r6clvsR5NhSKr4o
pIOAi7JWy9KdZt13U6mYAcgcHYAUQI9cNZNSMf2T9YzE3RHCqWXqGUWYllTCC6M8
WrlKrYeoZuMA/omSI+UxFaYb2uXQA9LGnnJzKmoEjheZ8ZV0W2wYlW8l9tpvQQep
WI/Fr3LwyU5ni17FuSnR6HtaOj0QujeU4t1zVvKooEcUSg7layNn1GRdFYuBKAbS
IglPLmZpOthRoBaTf5I+fPOZs5G93Vnh1GNuHteiCVQKSl6ot9KqiwHt4aoOAouX
7ogeM4zXmAxAFrpUkvXHe94f3+oGYktu6G3oyWs0zolyvrtTqrAiZfhxWcdKX/4f
kmG/ijb78QGhFEJkRw7p675fuhbYUNlOLQyF2B5Fw/ZbiPSMa9SLRzQlZ+8nGW75
aoXCHQSSx1b9LaPnUe9O15+wFARUwS7N79JbM/K/UlMRz/VwDVuObsiOjSPLToou
kSWEVjCZBUMW/lLN2wKAXodiEBQw4yd6kK+dDtvmV4UKhEISX8OWNY3shk9AJlGS
WIYRSXkPcdj0BkAalrf7xbwcWhZr1Zf5UeW6NoertoLDkHHfX1T6DYKPN/XhltpU
WOuz7SsazASgsOKFEoYC8fTI1PhUrvoLDr9d0Wka0XH0DWq1aUN9zYJCVpkPSr6y
ngCSvHPDOUPV5Y1Xg28Lw8ruy+7xpAcYg7BGYfpYwpTR8o2OtKr0qoIS/rJelnW4
sECo+7i5R6ql5WKJ1Aph5TlydjS7hwbo6f1TLn5ZAylQkqFgTXMw/ftSDdQ7uPaR
8nRG8Z08u9PY5XjCAZAGEAOBMj9Ftd4GvH0xyt6v9JlA35WiZoLP2pwR+y9W2K6d
RnhEjFOZDIyvZzcLPyRy61nQLj+8VBqCdCUizF135y6xR7H4nHHjP1F9/5yUHq3R
IUGgkgaAbXhJr4CBhADZUCt4UdaoWyB29ogVCJ5GO20rIKCc6IfevS2VCkcQg8o4
IVF/EJ+PUNdj/WO7AFeTvZkrTR0PyA/cEG2sK3ue8ESKu/8kNLJ+/8wf6yDnhgHW
xObJSFOkp44MnOmNWAmUVdudazDz/UvwWl/T53sDUFnUfovGsrf9Nm1CvqGKcyuW
7lUVFnUzzqx+q+ui/lB7DVaXU9X+ew6OoQUwqq0za6Gg2lLs/cNQUI+YBgy2Jjyf
QThCOqnnF6+pZqHti2Sy3SrHRyXAP7aNNsv9+oj37MUibwjiNALyHrfQ9xOUX7H6
Wr1rgygCu8cBntrtMXTnKuc5mFyuCkUDi/ipVYxtrvk+Bkqoi3+RyqkCgX7QQFxm
DYyHH26tv+AfEd0qQvW6k2IE+oMtDd66G61FcqD7gTd61UBiddBgEnKWpFh51eGW
XDz7bfRuZ49PLRnokgxEPz/Ium2tZWfV/zfJo5h7XNoqgLdm26JUEIOSFsmOmJG4
cNnZPi9NEzSw7tDtN5XBct4TYINiRcB1fQq5kLOIFK1yPgHtctGFJJLX15fPNdk0
TbEzKK2ACsv78ue67ABb1zlNmzlXFq7X5PpD/JRTi3KjWaeVvsbSa7il46L8XWsh
T95dIQO4CgfkUI1Yw9vadOPNSks5hV9Mf8HQXBprEnJhXn5u2NfNcHVCSn9/v4He
e74prjOSG/3vOyEGvmWK4QPIKk7WFGvuJBGaL6UPVuq0DuoN6g8Ji34jsb5PLzcR
O/PzlVK2GdE22DFGc9vO+RPTZyh3VpkF0TgOgJwOSlUR//Q7bF5s7IGj+ilp+pRg
LPN27WQk56Lfnvrnyo15jWYb0NlkyFeYhxSLbaI8hYu1s5BLcTiHYhqe8Uqh1efP
BoDSkSRr1GTvk3K87MiDpJMITqYIbDJm+e5D7zQb2Bjlv/QPxlp04DsriHyGcSTl
8GIeg8nNs715daTGxXnuzHzUz2WRnxI8cvpcWCid1VL3Y0uS1O/dkMMd1l6prmmA
25MxWFyQucBYYBfaiTT3klBaLKqFQIT3V20QL09G3gGyw51dNRnCQQ5B/SmAGNUz
0ko4k0i2GwcvdWavoUpNxUTjcQ2wt4I/Tr6jZYR/g4jWZ+lFO8Ia7TaX4EoPwuFj
svsmMyA5ZiRXpG/Ot0ktqG2XGy/fAbAQ2z9a1ad+H6qiQb7aaqBZfcqUG28bdeyw
WSaBnJr6LGGaA2LzvcwQ5kae+35bFX8pnpMnjVsYN0C2ciwXasFpgNJgiG4GXMyB
aYAQ+woJDXYe/kvTRwl5nd1+TtKZcbNuu0OIENSum3uJsT2uD2Xz/plP0nMYuZWh
z98o9bhBgmDjGXN3VTkgRID8hsMCLjZk29JocxnCfr4BBfHHW8h/V53Fl/jwcCx2
mGiMi39speCIf4LbqQHUOOPUoVNMj8Lbpj1r7Pd+uC1nRcB8xhoquYUCAXFbQt1S
FY+JlKnOqhL+s7XwWhJZNvwUAn0D2nLMcUCYCchGMNs8uzXgYlT91YhyaLE4Zl5/
twb+LvCIWVVmqKYWewQ3M47RvKbxISW7vQZTlzIjUyASH5Cfk1byp/VyPxRMCX5K
VsMjT65kz1WwIaSUFsPRDcq2cHnckYqNTAVrmzh3aiZmeMfo8i24BdFnJ9tiCwiT
V9eOnFw4Jik6Zd/pDrD9gicyAEB19XhQsv8xJC4I5R1SQf+ex/RUKfuqtPhIH4Qa
nDoK1ZmjMMm9j9ss6astFZgg7uiP7H89P8SjD0jPUYplRo/6grMk3joxCWvddj4l
lpVA5Ycgu8Jjd06VF6+i7VePL+U9fcm/JkI6bGVlBd4Ckt+jqhF+K1F0LV+t82zM
zKbJ0Bbxc+TV6eV9zPd3qfT8CJRy+dA2AJh2AsGssPm45QKxXdky3LhSzyvXyFQO
WHXaHSRPDWXS7s5ZVGpT9yUHCG++UquGTX4ElPXh6ryArnT4WVfUL1v3wrlj/WwO
fpmWTxVCpUa5eEn1DBis4I1DwI5CSxYEZTjVse+xTfHNxAdmG8KURUUYkVTIEDvN
Z35lgRnah0WA+XaZb06+0kHJS7vUwd5cZE+hhQucIfiRjpZzstZKd3R92GS4z1Fe
6bRtIh66VwakcD7JJNJm7u0dwoIbZxnZ6uP8noyBtT+QYlvbmw3GgcgDGgeUVADn
RS9igs3l/lMmEHnsHEGf0iNYe3i68EMS6JjZUWA+L4Vsn6nWx6YxTNBeSlT5p0ke
QVNvC4WDMtWLg52X0DUcEmu3ot3ABkvNInQ0ZTheNL7COUH3Z1cHbEWexBJYa1NG
wXbUwPfs6pOcrKdiO8hqOb6PesxmXKS4KKGm0u3syGU6CvvQyadVi+2ZT1+OP7Yn
xCp3KiRL2aQtXypvWNjOCYQmrj1BLBHKg1XLhWr5y+/jBpkjZRrVN559qgF8O9oD
186ArwQ6HxGfRB32Cu5ewuwpC476Y1I8eRh6mHB/Wad7T/s02qgPxmWbVUUT32LS
pSj5KHx04LLyilaZ00E+fcGTWp8++a3E3Og/fZZtDGKRfibfPLgtiUf6icWtK8rI
ToRW/oUC+lgZEqJI/2F/tIr4objoeB+qu82o3qOKds6sf53k+7MHk75k+3dmo6ta
g+pmZgg/q6eVku3vJVVq6p1c/4KoDc1g5j8HBLvfiPW/r8dYa7DuG2sXkEC6ECX1
M9T2ZIyDGeydKdiOz5lXijEJeqAI6wy5jm/LipcUob6ZSDrVPfamaewLbtiePjKw
dbwnnr2LTV8MYKI43htpTuAUtHq3akRb7/wWrU89Vii8NuykVxBzXcNlF+CcDYdB
nsb6qiD9sFvfj79kA0qUvGFpkRSNtATGZSxQqXWzGFw4A5f8r8aaGkYDqA1hH+2B
q2HRRy8fb1YYz5+6LupRGvmewwKmY2AeIeZmyxnY5/nkGzJsLx/1l3qGttZWpcUh
9vyhykLH0GtgiVqOzTBntaaTfhqPmRpi0Ijoz7t1zjvvkTWuVr1Qb9JlmIND96Oy
P+WSSyBEwwSIOQ3eDfbsHyYgbIdnlYTBURYdd2jY7er9YBBSnsiQB4DlyHK5Qj1y
ycyx399GRZURZA8KjICvaI/CH1ttOl3/tqRfpq33fdliCxiy8YB+vFRI/IiyiFHn
L04/oA2Yxd+r2eG9OasiDKBoWVosjyU8RoHdjVcqvWe5u2kPWlybCzvoLFZbiGQl
curX2K8GcQ00Wp5Vx9+xiJhR0BVh/RxpLIgC1sUkbJZbz7pz04m2Buhy9szYoYXz
Kn8Npa81pgkE7RTdJuo4aZ4NaD73QFhdZZfLf1n7ApU+/P1uJ/3Wd4Sf2f5JWPVg
LzPBJdkTQTnLc5X/FjFOdob38XkkO26yB4+Snt0dG5hlm8uUGkVyFiBQZMYniW+0
YaixZlztNKRuE94H33ML7jqDOCQCgZyncFCM0sujyKG/ebffK/v5KiXBbgff1UTC
yfPjJDlkE87zONbZ/ckd57TqDeIHJjQBSgQXB2qvwUMaWD68Xw0Jkw08EYyFIWzS
1NGmMMvLsdony3VfkIHMcWT+DBjeWOFxEz/gHY2mpiXzbjlx7dqTsMd7IrNOh9ub
I30096FCZ/0VFp0z4QBaoH5Tl0ZIFV6Nu+KIGZ1bHIjl0ivfUqU3446sObbLXWIx
MO7CNgvbJP9JIsQxvEpiwCt7JCNQiZ/ipfdNC7a3j80R/PAl5f+gfccPPGydTlsX
wQS5nof+gEQabcfYmTsc9VplzF2vhZLX+/ScMDAb2A2Z3NsViv6r1B1cfUaWKxXp
XOnirjbFvG6/BvVSMxfhC72Qr6BZ4b0shxZ8sGhvneIZTwXhvV3IuAKy7VpbKlkD
POhjlTQHhWUuIf/QrOAVLwKrU5QRBp+I2XnyW6IIgU2AVit8Q5PoECMMNk+uKNRd
7ZY8BdTxqEU2YaM/PgYB5LVGiyDiSHq4oCoPsTjGNAdAeO2mTznxpyn9TSGB6Eto
I7orSYRAq6tsCVrFQEm2Wp7lDDmENO7Wm0Ra9seoOt9VyVQLw/ic/F9g47WfmOJG
GuPgfXaHOrGq4K/bGBFrS1vXduakorGJ3i9/SmM4UIO2lk7rLE7LV7IKWqtQ7TrH
sKH9LMUsVswwMRk239r4BUU7JLS+TEnXR2b2SKQOOOlX7LuP6HaVnhz7pgIQA5mS
CHa3dnkY3dHVCBghbMc/geASobLtJ4u2UYJuJIiaQZocmUJHABNcAQ8BREAqoE+R
gc4/xx3oNJzpR0/uH6Ho6UpPsTP7rqUgEr2kaoHc6YeW7299FclrIPBSfJa2AJDK
LM9cnqRihFYvIWAFnA+Q4edF2Uh+D96wgu53Aas4ne/+PVVFv+VT0raL9RNneMKZ
3VhftGtmIe9e3tUwzaOeAoAnk4rbdV5Y/UPX6/syhoaHJHVgLjgOioL+aDJXb8Mx
X37nxwRzRAiCEfr8+5w1ViLe5pIZ70xZVuFQVVCSLqkzTcYbpspI3PdtNnflrsGV
CgvHlkV5XKH1GTeUEsyqMA5UWGID7tDwjYIDLEJT42Q47jpdwR8w8JwMm6dRec8x
4/eNIaqwiYtA5F5EHV9aK3UUFxB8KyXfPVbdYPmtAKCdxb6G/oS7o0DGTnfHjLUl
wIXRJXTXChINXdhfOaBLZm7bKJs1IRK2zL8A+t9Hx7Bhq/Qq05IYSlMXfDySbz+M
lKJE1tbE/A6xZ7XzCNztlvsJLveRb8LYS4Hk9Z9c0JrUI0SU51hHsxkKEtDLy2/r
Jt70HLWfCAZaLZUNMiuTuBthk/+e2sC2sNZiWVFMzBAeGKal1bOzlstXe/Lb/riy
NS3Pr5CIHDpG7IKhzLNX0lOO+6ZHlKl4QVsDack5sJrX5qWINISn5+EDJs0jbgs8
gkBM81B2ZMAIVqmnOHa4ePPZDGz4ZTSklzp4cTJlE5jwGURayf5ahl8cdIUQLTt9
VO1QzRyA1SjwDkOsOmAUDBUjpV8gsCjGE0p+l7VuaiaaPGKXbYzjAshC6CyGmlzH
7Sjhx4nxl1MRrdFeyEwbMcG6RpoRsKraCmymCJk82AGcPYQ6fEAqweZW8h0qFfym
lzMV5XQHRftXvmMe9LlmqnTUBPMCIEgRaOMFnjYzKWKsO8JBjNsS6QK2SpM7Hv1m
z80oO/v+/2RLBwmvinUVa5In3SN2ZwhCpYWIUwZV2aYOTiLfTlieWNChdqns2QMx
kgRh88VHZOQYFUlGEMyrh3T/zyKuThvCv6wOkqNj+lbUQPC7fNGrrbom0qFjWHji
Zf7NrNctvtqDTrXB1mpwFn12VDYtZmXwIN8olGJfMyTmZxh4Hjx+Az5KEh5JDFhW
UDICkcP5vs94RR/mKXSWFrq9bW6YtCqoPTI8OQFSrYbbleEJKyyeMvNgoS8P3My6
UmLqD2WpiH9YbpctHJsoiT4WZyw4Zeshu3zoZm52rxg1g6Ca38cmXZLEIKh0STtV
IYDQ6fo6s77Y4HsZC/ByCqKCMlQzXdhSL4QurTMD84e7PPbgpJPNUFBAt4C7WWZs
3oURk2VV1VBNNgFLf7smOAfrpCs49w0kBrKyN4PCm874NH+xgT5DFd/NPRdFlNDT
63Bp2UvZgdlPr1kUNpC78nOPczLF7B25c97wDAT64vvWXcq/za+pfXqtFyljVL8+
G4LNh/IJz1vsAWz05yYSmrfU1nbkeH/NG65/IRZPwxGfTlT8Tk/yl6E3Pu/JnWEv
gDW+zkB9fKW6KsXDO5EDyJXC+Ys9NGgp+6T/lSDA0F+vUnqkWRXZNmX2UbIsksW1
2oIgxGWgAYgdmqtoKLy1ZykhPGyBP8ApO4I0DoyXuJPZulwl8LDL8s3VIP0427pz
TrFHg7f2hIQr3xoh0hKD+1FWrLOdkoLgZBz9uG/9b4IggE5XXbdtwC4LFDC/gNUi
+N3eFg0UJief5wYBx3QruJ0MnKZTXI6AkZcDT1l/CFvfB9M/q3uV+sXDu7efj/B7
wH+4SttJsUfNy5dRIkCircPIQ7jnaBK5WnaFpb7tHFFDGoNf5XChj6gjfUMl+v6u
S2eJmxxZ5cvKJD5vKBAu2Hks1o6aLzvueZzvhpdDjcpkQQuflh+AMNN4tJ3yOtDw
FxDcSFbL8l9zRsPVuhTx2SJtr0lZ4c51LL7EaAwidRfww0QrqcESBBn8qtc1CHEf
YueLlXW2yV/10Dbf2+Z0NsbX7ngvNEJg5dNn2xsESBBriy3H9Kt0dlwFosj9L8sX
YxZ5+UM8Zvubv8xraRYQI6GkYTd4byX9Xiwdzt2EVxEiOgsTU2jRN7j2ocJJH2Wf
AEag6vXd+q7W+IaoafoX1ug9/rFGzB8oORjXlB2WaKygMzsfGCohTtQSd6oX0k89
IO5MqxapqUo8Hur/Q/e72wNi1pCzZVSOz2g4rMjfFfuydBsyUG9ucAC7+a4QeYHH
V+iViUyyLPrI2mC/f/LicbStX3Njn1SIF3xqnC/QD9DsjGhZJ29oFefUdD7M6tXz
WAeU23s2en4YHpMTtMbr3xSDxpO7DizYK6Z1XKB23mIG3wqAGTIZoczWno6hVO6z
yIsbQSTqD9/PX/0TgcjYgSXA/3ndHX6MFfJ43dhaPLo5sYO1Teod5lHqAbdzFjYN
0azraZFy3G17r4/128NcK8eb6Y6YATabPan7O25dKJ77Z9EoBqBghOAg6Yrd8jH9
0zqvLTqlhQ+58xat80e1hmfBsJ6XG5iagF229eyR5adKy797jgK5aop7Zf5vZe0C
fWgNriiEcgyufxWFys1NTRY8E7lQJ7+F8oyx5q0cPHt2Hr72O89oWEKLTRImKuIh
ACgQyrxQFivW8/VzmMXboPy0FWvO15lGVAsvNP2YiUZxW3pwTGzb3sTmfAT1Utdp
ycBGIKwO20b8LgaGxKmhZFA2q+OmIl73JxB2ZYSDaVp6TSJDN1pi+LDE9EQd1+uk
WVuPcE0KYBNXFyNCfOrheLVBe15uoXDog+jts7cBQduDItoP5gVr0q8Sqy0pGsjK
72Ftl3rIrtn8jyKxg4l/TWcCxDi3+HgTKaLFsXX+aRhj3jN1x/q46lQxANoQhtSX
XjLbJjOTtx/x0yzCvSRYbewZjNh2IbetL9CjTt6wDzzQmjDb6g1Imk77VnTU8GT3
39aTLNtQllprYk4cDV3WqzcHjai1Hwz+prVKQ8G0mX31+t2fU5kWzr1G9JQ4DcRA
qZDj8kCuhTkDrAIVUwXFOoYyCcp+7XJ2cdp34Ph8nE0ZqixnCgT8YYj6KGnD2FOo
it4Jf0kOTvh73IuE0i8DKCNT1EOpzu3mvW8gCiCnPMc94B/UPHGz00fiKv9jOT5h
yo38z/O/tFvGZRU5wYA7fFb/mR5vE8F9L9B+eblTMJhrHHHzXNnY4tQTqwV9/kf0
sJksc5Ng6t1nKN1JbHf8waaJkhOkW2l0q6sEtOV3vpF9B8/Hk8JJDo6kuXLu7UJD
mdu3YpAYhiQchW/6uypccRJYuEEZ6T0O3s0LCPjRHArW+0V72qKdpQ189gC7gsGR
qTYOcYOR2Cs8vWRYLHUP+IEOiWPIqEqMIs3P+KL93IRPBomxpUuPFmEvccKIUy1u
aMU3tRBRm4NtsBjslWJIxnVeXF0+wqGxT7NoGXV5cCQpZ66JZ0iQQGTqQOquI1Gp
lhL/pJ6iDQHtBLyuKkPL45/szpY7RZ5cbeVQB1Qsjuink/5WaOtVYDqSboaGzWDQ
QqkW0z1yobdmTSHspVYhJkKSrxPL/K9AiHZPiBah+GZZ7Df1zMX0k6q9IDfKzp45
xbF+1eJBjDcq2S2qWpubiK3mV2uXqs7UPEF5bslgBfVMqFgJQ6r5aoXF7ZD5loue
iN6QfJy9Q5cw4PzMG8vFgR/MSwSJFFlsNazCLqkRwpUltwPE9Pz6gJZuAJWnZ51k
lji4+eHKE+yo8XAwotNxcXJQweBOBEy1k0YKVS9UbbSG7imv7IsxMgfTYoc4xIdh
ZtV0Bsi41bb7KR25oHbx09LtdgzgpZYwIGpGXXZNduRWVA7aD2SjhUg4W1zu2gfA
EX4jqOvzOvIZKWYBce9koyQrlwfhjBV/OxrZVZ5oCPXgYqyQ/CCMN7LlAxbaec3C
yksHZO90nzfHRWc4J/KTXkAw0YU83jh9Og+8tol1TUX7VjTBO/NPc5d7lYxNiZKU
DMQAzKo4cRHm1gZi6H6b08Z7jO/9aONM+hqHJ8Llx3x9RRG5FiZq4Idg/CvHBZHU
5eiLpptPjNVjruyDHLVfxTKOYK3pkdZIVw0uXz9CbUeYHsZhiV5qwXvnq8nqEWBo
6zbPOTB6hdkKD4f5EML66kSbdCbnNPhKT6/26xdENVfVp6kpvAXDEsfiC2riQRAc
UNsfkssKHh75tLsQpaP96wUeYkdR+oJKbZvXltIrOv257jIPmvdMQGoNOrAAdJlE
LJ0PoWtlwxfgIrDCmdhtxh+CRqJeb5hsmghpeJqNHsQDU9RkzDpuwWXopyD1hh5x
ZgRs0DvYd22R3k3G2GrAXJ69rq0ytfr7mQdcn5M9M12x2kfZzIvQmft8+Nugkrvg
M7JV9ihHmqYUftXi/sbLnZIN6KT4iESm2duHzLzFjwpMDl5/k98nKDAEAqrojca7
lpX0KJOgsJC5bIMhzhRQ63kkIbkpuD0eXQ519xllZfQhyKQ6A39goK60kGCDWM0l
m9Q7bwbCWbPJdl5rNVQwcjw1ePQ3QhPA2hHcX7Y8qfI6IlLMf7UIO1q4cjSTEbx0
lNZVHwrL41VJXtek1b58J+eOLisCGeIuF8Ob1sM1TF16d5Zvko71xPu8bym+qXPI
H+lPIKSuoLCHfQXmRWz3kWLp93aehY2wUujPZF7PiTi2pvIahWmtGpg9vNPDRe/0
QaW4eSFkvdtPRLDdpae4p3b/DHMF+DmEat2XW4R04cYUyj1Wahzx+MDs/HVHph2H
38AtSjTn8aP4EJNwcOE8XcYGbKOGezrhKsme6ugVZ23Cp/Do5rrXKyFLNsA6ccA3
axVawrUHhy/33PbMdJq03T3/bG/4rmLHh7p+fVZuYR5n00H4C13dXSYo/NFXChP4
3fTQcmXAVtyRKS+NidWDvZmHmtl9614mdilj3aUPiklrdmp64ZSMEP34v2tOV2/D
dC3bkcOMIBYDSehenKqKDBhIIFZLDskOw2ohe3TbjBIs7Eji7q/6MPo4iJPvGESN
6HZW+9lUea74gTJcOl59egKgbllO4+DGdCPeZpFmtKX9xfqBh4983Sk6D4LtPL6Q
YF9dHk/ttjBM++OSjxg4gJ17kZKyAwQTcSPWR5v7XQhqE3Ny2YlILSUV1bMfsELU
NZOdoFgESqGWcfjyaFIveNR9CnMMrTmXU4VY7fPUzpDtf2EhVOInG0sb8EcODcER
Z6CwIC56d+rxw+OLGwTU+qdQ4C4cUXKRQzcmel0ilrgbBguL2n3/wixG7hTtW2Bw
2d6bWbnkz+/rRi/1+sy4VUOry3ZT6Kj5i9eAhSkHMW0BHBkLTdDDilVO8b1QpyWj
0DU6Vc8SYcLsNQ/PqbVfilwaeAevmDATvPh9nS8V6Amvb1Hww8yOdEqyKdTfmrin
D+K0G7tiw4xQVZ4bE/sgiq8kvNlYziCw42xdHD0LHPR34cOziD0RKPArXd84w1lF
mSAtZRVdcnP4UM1/ztwtzkuopBHBhg6KI9vqeW/kx2BNOl7xSlDy1nugq470LN4o
z1DHnQBkCQ3WsxWQTqWE11VHrnqKjFTbELbJI+flM5z7n71pd+QHfKFupfsno1yw
uSsJr28sYeyYOCcya7PLCZIqRTTvm60OA4yhWF8eGdn4s03Os6N1xhX7wGF5uxFU
hIYJDvpaMgK43iU+9g3RRqQ/Wo8VFyx8GO7aCNpPbAhogQHDqmoU88ICv9Xvrc1t
ci5IfFtvpALDf50MUo2Wxz1V1CK5smogx/YkS/XRPu/2BMBnq7dARwaPhTh1231o
oPYM0Kf56ZfKPjs/L2mCGvn2s/0E6tv/kybWJzEVPxo1TMTAhi5WsNU6rwCQvK52
rDA1FxKx9ktRoIljHx3AMjp+C+iSS/ljdrBuVxVcShb5BXBTeg8XbtDkBDprX4wY
16FrWtuPc151xqGQ3wOQgo5p2cqXflvRRXodu73SbjtF5JgOqcSnGXzC9nCg4etY
2b9tAMMOztNWCLzPAI2Qs5nRgkAk5ylrTyoWxUdb/lOujwQRcCqY9o2onTq9yvAJ
mJhGQNvN7JqEKUh1HpZkV9g1q2wPKhBd1ILUV8WIwUrgixsXeDywhNXAZju7o3jl
lTQFoPD/b4iCOLwTGuykZUYG1mPDS47Dcd0qNUSrI/WCItMSsboemcyDR5gGeAS6
Ub8VOuKl4WnTaJXyY0sVKuo5qTVbshC4pJVFsOVCM/dXeqLTub/9hv+6xsreZ8UW
VkcgyZTuIITSQATHOO/T5K1hVUq+DYB532NkhFNuKsp8xjPDGKtgmReEfGQtY3el
V48J+baswb8oTyEOdEPqfevDNiUmH0HF4Dwa3eIdD1dGhuMO/28J5U1ygJXnsG0Q
Hy82MKcvSEousd9DUJPjx5USm6g+ziCdh27bgqzGGse91t6r038MiaQxR0fnmTkV
pTGQUCEjpZ66+zLgNCZCIUipxVIEO6Di7+2KHKktE6u5XUD4264NH1dMaFZiytEY
pyD33arlqwrJbPMwfMUiZJL1xlHNXV6g3qJeBpdv9+KLZcDss1S1OJd+VrcepZOw
PU+qRZFxK/IJMlYm4QgCIkdKz3GSq36jp9xr4yIUwjFy+x75OwwNFICKtC1pgcxA
Lm4B5O5eJuQ84WHlfKXvmzbLSwOQIcOz4mpwoDAJ6oWTBrgVgJMPvRzdureCC9K4
Y08HQD9QndvomKhCKQBO+HoAHLPlgc1m1aOBXHx4wOI7nVEHVYoZLuPoo8BJcniP
ZQ1RIaVVWJ4bygAj0FEd9XMjKS/LyNUMVTMzC7OgiGQJr/V+TcXTU7Cg9Qh6nOdI
wDhsMeNAW5uPWe0A41soHo28VuMvlZub5CISh1vQ/9kNpJGkeDO4Gcg194tGxlBG
Dtk+/986v85YBQWwtcfeVaRIdvHSjat0A62R2ZTJNQGArCVucYtWDcRnR4cc4zIB
uMdc/UaA7PF+JCO9J8AmaUvy9x3Ezw08IfZU0unSPiYiiT44A/7Vgd2xIiRJ9wcr
7AYHD3vuLiU1J431snJv5Bjlmy+E+4Nqee+APLH4Njm9GtYFHTapB66pFWf3h6jd
T7M4bE9RF0rcVdkXwLHHmHyYxzrVYwONaaWhhWFNczAsvOBRj7I928++VdRHfkmy
0Axa5cvVOjvlPOVo9XO1DtHBwGzQsLuDEj84ZoGFEhO3amtn4bo6x8SRSV6BI7Bi
8h4d4rlfjFSVBRX9V5Of80ukO77vzqp1e2m8L1vQF8NQgLlmc3GYBK4V4HGR48a/
FtTBFu7B+mCQDepk+vgHHrCyswZMfjaE72DE27j4H1IkuTmHn9mcl9Pj6vb1ZjFR
JbYxaJbve3bKDhr13JG3B1MIaQAiv/YN14fR0uy1YIkmMJwgpYy+scHxdlUn1c7V
DUHHIvN+Y2PL7sbiCbtEOHwJ2sZhCcUh/Qpm1Q1AobRb3Wh84mSE5klEYzvngnXq
nLqKYqDdXFhuQGZLixgySBjsrO77vOFMMj2cd5bnCbGCJeGd+D1bHSRdkWFEc6Ta
zaoNXJ0Zf8KoZF5XgT5gkvzrLRtcYpscaWVfS3+L2/GkRZSjK0CFI2QKoc20LZCu
t5l2po5Oe0e6wD3d0xjxcSVYN2TNQUEUL6Cyrd5yzAbeckLPVHSVLS1DCKyC7qvn
E+1shnLM+BvWrgk5V5/SBWGbxwkjXaE6TAk10YiNhcu8Sv9XEVEkfcoUPwA5zTyf
wnAJmS+gDeHEyiiujFoyzKkJxeNusLa8SEmgEmqEyY0FxMks4pbO/ExBcpGVyuAv
5d4v7EJgz7A33ME0X+K49Q0ADceJd3vw6l5NcleyXuZBKuJdSdaJp6y7SNgnbcI4
ltIsBqv0FbtOYLYpIzC79U7x1yInL4lJ5wHe1OR9Y7R9Qek0CM4sxmkpL7QUj9Xr
XbKyn1X5rvZVf8gunlxWbVOKL1R9+sOQt6bT3hgaZWcMZpnAKo2VgA+5PuReX7ts
jBAGwLvttdpFRwV+gSpIeq1OJn7yIbC7XQg3Ot1K1UhaIeRtRNeXSUsgk6zeBJjl
htXFfV9fudKI66yJqBQgmBgbdhbFmLSDwIgffb0KJZeiTmE9GvR5wmbeFMNiU4HE
EZHWQrVnkM3NELNE5FBszHdjnxVRKV9+z8j7qz1gW1aB2SGJkM1odRQgsAS2VjwA
zIpZLExvk4/oT8Y3kA5LbEjiKsckeBJDV2IIZyJM66ralaYYDHnCld+7dGVq7Sbt
icLKK0RihrB9WsIKo2BdcjyfOr4g4C4nDkA80EOW08BnnQmyoXfoo5O0Dm1pbukO
BuIecjdD/krWeXNa7wEbXxMVh+12vnV/mAnmViruR8r6OkdwdAWun4OuOhcm0omG
EryQUfrlIJ3WYAi1ky2M2Ri6QHOnVvmizgbSXN4qIEryR8Ax6NqxruClXrK9hL98
UY7DViMcKzWHw2oH7Ck6OhlzCHJXPuugPrvtwgqzNEMTe/fbxGoHCofO5Bvvag/P
fNlUknP7kY41jIolI/+AxHLuZeifufNGQQDDyPaCr+N4C3HbrrTC8MadIg0G3zqe
LpEjIpf5VdPFadNPndnsWQL+9qaNlDptPI3i6jvlZX6GnNBwlc4+j1rQ7HZSZEps
7i/ZHax+KpY78CpMXU/q3VvmoYvDA4VYH7nCrm8jg+4n1vwtzwfxSRbslwqLzWIB
EIeht4xxFa2btR2swXotQgLm+mAycGtNIkllfyF7PF/EWRIVikxJHiwFmOeUDJDC
vk8hUdoZQQbG+8qM0GWW/sRSinezZG0MsFLbFDv2nRSMw3aBJtGML2X7RP/TlUQE
jxCTMHBBhcZMVPUHDagT+eDXjfS/BV4X/SfSKk2MI+5C/Sx/Tr9tREinFNyPnwwn
QdHXL5iRvMkqVNnTdjPy1RmFXjxCAykSsUKyE+BoA7lVeog5nv5fd0OjTiVqYNsW
mfybmf8gZA73VsDb3iMOjfWSnt/CTupBkJCzSERyCKNby20ZXpVKYkUkfMJX6zxr
IbYuyf145/hAk3cprtg66CRnAqwGaBUj8Olv+N1B4VC4LV3gZ+IbpYCHh1TQenq/
8kiVBjh9zB5HyZ9lcXHASGl5J7upenYXe88BxC8X/DILDm+O9AXl4i/j1dYppVBq
o8Ay3FZHOAYh/izZNOB3umDrD84QthttIuH95AUXg3qp4kcy+UAyuRTzVNUdm0sA
zl4TrT9DV6mLgsGvccRC3hICeWXBHTOqvVYrAaC8vOu4BlvHCMXFjetFQtTGWT12
cYuJPDRsuOFveVypvurCyyLa4MJkyqTfsNiNMYzsAupkI71A9Nt4r+HmT83d4QdU
kEyeBDOzbHWTZrZSN8xM3Vr3vVhYl0vaG2cMTYy9BmLu68MiM1hKYJ9g8ATjZCQs
cJEEBeIxbaDS3aHQLzLaZcAE4LBAYHyUqfqXiYqNheLscSPKnTxWXGTRmkW3IX2Z
JyUHMwDZsd09UQSfTwYufblde5zKN3mvAY/hxEWbAVvyQAOaQY9W2lAXwSLfQDGN
BsYO0dbe8uJ3vqtHYTX7x9oO5aaumLhDx6jSmKuc9cQONlCBdWU17LtXOz6co01B
uc3sVCSPF4+Oz959HIyAe5tZ3GHaUGfGiphrIEaUI+4CaI3uJ7rP6tL2rNCAlq4C
pm+wUvRGwd/qSfaeeTjpqGzJ7xF0gB0ZDn75E1Y0Uq68Wd9ZedEcJ6RdG0MnMJTJ
mZhptX34W5jWi9+8HLfSTIubD7yWqNAJPsnVqNKJZ7w29lU45vd4k81nzGHck7xC
IYLsL2izrIH/M32f5ywjSQjlWOko0WgsXLkfxt4kxzAD4qIqKQcabk2bIIOUJiIQ
fHH4D3BUG2WX2t2HwOYxEUHhhK2j8ZL0ba7cDl/vFsJ76KGuZENV7zNHYBm0GRNX
MwTBdiStjgbtJBMxEmv1AA//XAx+QDPFQp03iFkAVd6yjixXDWJb/1iLcV7ITZ8D
yEoBUILN/JuA0OjeN/f9bvNv8L+hJsWwJ3HmptnUqnUhtuHJINPsN16/cwUnOPq8
4wJGZebuTrGHVM4ktmR9kNiO0efdlOUFmfaG5SPxZbFwjpUL2iuPRRYNZdx1kNSl
PcqIwZ9+IoOYV7nQx8bBRMZ9dj7WjNsRp4+pZlAjKLmaeARtl/bZy5Tj2jIG0lBG
94dSef8zGAaG0P+rplYkn2gi54UZ2g/j8JEUbcuKyNW+LP6CSlDzrIIR+7rP4Whj
2vL3Je49QSWc/KgVBTxMf/fvQt8qq+hKIIIPdN/fbZ4FqtMJTtZKlhsdc6k7iVnJ
L5bcaqJkq1STu4Cv+ad5gCrZqLv1LNT5VuwFJ4UXEfUd+BgOyx8dN66ccLHWGht/
G94Rwp1HQUD3KNzB8cwzXKtNvZFW0pTtIROQzZdLidOEDfUcbXwTnSCck2FNpBur
2LXUrzbtI+k2k8eibLAJ1Dawp8XFkwrOdg6XJJ+2Zn02UgBs9cih4dw3EqcdgWei
+HPJYr6kGmV+4p0FiRbtBKjMxw/eBiQWXjruV8h1XAmp89tLHlXJKiCtCC/GxSsb
FA9g8lsjABb4XhLIaSdBgZmp4qpI8jWPQirTL8IsSPfYI9W4uIergnPPezkgNsne
wkempwoslOMOMM2YWYd8BOva0eKdO2dcqCSDvBonxJ+iFIRTv+fFHiQIzK04qVUN
xe2w/kwG56Uuzug1gtqQ+ycgU+umOVCSVelU298wqQNjr+0cH5yHn8n71XTkQLF7
JKsmRntwT6M0GOrFR5jOCd6mRSbUb7R8w6baCiJfmhbWIM2TPI1WkZYAIDUDaPs4
aN7XrFa2j5DYeWh2MUa63L26jU4aVBqJCZfjtjiKh9GlrD1W4YMWfkixqUm+AyEN
NNgDMPtbaZ2DsrJdTvPthsJl7tgR1BzN5+oO2RL7/lOJ1YK7R6oTJ66xHlfXbi4Q
gbiH4bqcL/TMbXYvSv5Q7lF8A4oPq3wL+9WFpyGfBbnXtby1YcMde2+OwVgmcbp1
L9qZd06XF1EfQfA8YJbNCXLBY+SUqeraW+2COjvrEznM6EO3zCaRERKGFGsfsfcI
fdH+fMQ3mXD6GzBkgdRY6F0Vskeg1slZxvJyhOgJx+LS07FQjEDXLsd7StKGM27l
v1RQTy5jcYHpNvhiSrrGfh/htv+t7smdb48Z6f+5dPDjl7TnRsZtDcafHs4BSlrl
FmpwrYUMGNM6ki5KGDdbwbtJ1ONkc5qeTFqohqlqG9d09AlONCvKsZr3c7wIer2z
Ahp151GZcVW47FK3BDbVdsqCkoLA4zAXqUvkOXRFJTTK/pG7Pw9a69q4YE8SEckw
zuV3ng4L7v//MygyIAxD9WyxRfQNf5XWoDbpLHC2RnrXicQN9GvL/d5EX/xo9aTs
3q85c9dTxDdJ3oh+M5tq+it725nTBao6FBe9TAn6EpVjlKNnZ+j5h8xy7jCaie/A
GhQPiPDVXAGLPlm8Wrx5/t/2UXf7JESNc6uM9xC5bOOjUukyAyiysgaVEgvfhlyJ
PlTc/y9YTH92BsdLe128gfPH4GAGUIggknKj86TVl0i2ZIyzXpxiCusxuEIQiGPG
CD+bLd4j6zE0jbxKzAIp17xMwDoyHPWHqzKtogl4UoQ=
`protect END_PROTECTED
