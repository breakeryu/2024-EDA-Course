`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+iI6dZKOSCNe6td+2qBY+zalnaabslIIVndcoWbR4Ovl2DTnPpnPhksbcHfdrFe
6g1PGp3xeLctKJUY9jawuEYgazpQPAA+HFnw4yJ83IjyTlvkGWWWtSJfvROmfV7E
WAHprd3LDDpb7Jw+6Nf9IDrf9IWwGd4ypbo70K6RgJ/gyDhqw6sue6V3Zm83xI1t
xpajcUgitxPWLiIJrrI3Ng2yJuZjcDTnBOVl8/EuXnwn/QRTPxtimwLTeRjcGuWh
Wg91A35A6/k29zbw3SjK6cAxfl5YLszYwH9vX0jVL/Os6D7qlutR6QfBCXYV3PQl
HHRz4NurWgIVyv7PmJW8ncCSWQ3TXv4dqkJViEJy5wFsDlxSgCBaaoi6eNswOT11
z9Mecj8wvrtPh2TLGMpZGmVBPKDjoPMlp0tv7xwtOvjBJIDFAWn7zVZTAakpFjXP
xvESFK5OwRoEHQbsCyPLeDMK+mPLXgDbX9Dk+ZyQfOzgiQ1POMQYmD3/GPFRh0NE
zpnsyWERUJwX6RJcI4yONR2QazD5XIrA67MDhKHvAGRnkg8lFPmkIEoZQImBhtVS
3a8edm+wK225e30bZIJH9Qxs3ujTOonv1tgqhVxtWSQhlk/xfruKge3KmIXy7HVg
NqbiafT5qfpu5qN43FGcgSJ7kf2BDB7l/3weINe7vEaRnES2nASUvSu6k1EZh+Sx
58bhwYhIVfRYhANoAy6qmyxR2ea7opA2TRvokBWvFrPzPasa/X4enSFg6OxuLIK9
JMUCh4EqoS9JL/VCSnlTWL8RP0bWM0bKC5VyySyxuvvmE4/miHpJvQh4NcaTmT0e
DQxYDnhZrTroN19zUn5WLu3fGFubcuwNkNwNYJfTtGleE2s6QDpufP1nmcir+938
oqIyGydMtCIFvGJBPDgmJgshDZf2JFs1T806ZJdS1puWsp77BkW+ZNeYDcdiNTWM
JshnPIG7uWgW7vLydgU3A8y+FO1VkjfTcSEoJdWEHmrFD2yKx1L2Ww16TUwjhb1v
D5KwsNN5CR34xuHIuIT7UKRK+UQMIcDT4qZcD1s2fnFxE8ul+C4rn8j/RDPLRnUn
J8gyvflPtfNg5zsCEwYynBOLZFdN9efzx+Oa0fKTtWyVg8LxfmGgdBeMQAdtkcID
dQvRrCC5NH0hCWw01brpq9YOHxYjVmQrfkulrnwY1xkodlNWUixH+Fx69TMT2Q/R
DH40C5CG9w4vcc0tQW/8ngz8NZswsjpP6prxYn0qtoayr6oo1P99uBIAzupso+dZ
en9AvwV70AGZYv2fpqzXK6r+xixieZZlubcBWH9ckXVfhqezAyP2YatuXsQ0Tg2j
LwT+9mycsCiq36HXsk4Jrj/awGvErFhgPEvi6AJ7YPByEgZX8UmWQROtIr64yNYm
ck+J08wN2A3j+5S9BAAn4UVuOhniYF0XON9PssVLSY1rgTO5uwyUomkgyF3s67bb
xmtx5F44W2E3BQBkk+rp3XpaRidW67+7GutcOpIPzJkVOMOPBzGGy+xZ7xvL619u
W5mDFK+RrrMQUMX10XosxQBwyJE+LocT/sF3VBKiYDQvleGkYIEHv196o+P/SiMM
GlJljLc25NJ7fho2RHv/2Nt4QuuM+jhd+rIgBcz0DgF6/S42ffOU4hvHrEKb2RkZ
PBAco7wlqnHzg8PpcmwlnTLJMvicJZVF2O9i5bWjo2tm8Pbm0g08GuKG9S6kVwia
wvKayo0ccx0yZ1pyCwSjjWZOR2uTtJHGt9EXTfY9/whObuJ+cuan+Bb2dA6OSmVk
BiQNfCapl+KQVVMki1eqJiQKn1BOZSnz3RPbiLltR+2Qa3z6e7F6ImukP0GoS5HY
ieRDZAt7//nrSA/Tv/BY2nCNo200TctjJgHlexn+jqZT8OaNI812q8MY3RWv6fuj
Q5AWGsWSN+KHwmEFNYQcmt5ntN+dgH2BtBckUW1uyiIQdaQD8BXUx3HEMlmhEqWT
OMQE3etsvlQhRwSDYXzDukrwUOLy6D9aYdWvpc7wAykJ7RKQVcbIEeRiApGMcjCc
aPKOgcmHoRnSx9YxHzIfPCGLKQ+gsRJsd3XvrCeHPhphzs9AWLkGA0dxd8Aen3ly
43xKtJra9EBftrCmrTIOhn1eU8aOEV2JB+ZekbUitjMV1xTijF/oGTFTia1bdjuT
1JvncJlBCyP5i5M02TfdTp55WHOs1/bFQb7yuqxUnmXvmiEPIv3hs6siE02pEBUQ
nTzetsrBzkcQloLZQjHeLJPg7TGMUuxN2EKfOaJlKUhwPSAHdKUCi4UNccJR4AHv
TuaI4ww8AQ3GYdvKUfKLp9mblI3xQ505WN9p2HtwtZ/ZtbZWcY3YdY6zVCID24GY
2wK7CkThbNWdTMW1VD4ZCXoDUs6rmzCJ28sclaS5Z8GctT/l7ttd6dTkAfg0QpGc
0ICq57ZPaix9AAzt2gd6eHvoVleSxiteYPy9W+NNjT0VovBYeCIIdFaMXnEyR99K
ecfS4y0u+sXfbp7M2l/+1hGzzUXF9UUIdPmJrXLhWlmOlQO9nyd9LadO8GPGHzJo
yNbk5OvDZQ073Ry2MERteR6ZfSN9Hjj4YYfc4F2QysieApgi2vfZHqFfJK+jK7sT
3bABzTlH42gAaJLZ91u4DW/F0Z5ljtWO3Np2Zhwy6dxKGBLX0JO6eEdeybZTwiQ4
LnTgucAE2Ec/tu/yQlhykiohvZAI0/a35Qbf1fWzSMZpjgSXJQwO321Cj8heBQpv
eEMupjx/QjbF7j2bDyXIXVxt8V1onZT2Kze8WX0bGq/yEWz6lbqOf11iCzQmMqci
xw2b7BZFNbZAxRWFt1KCbg0ZuiJBtw/XFX+JqWsbfEQaAFSOnM3DuGVjPjVVg82s
j+dvjd357i+oBYstzvKW0uWwqnbDU12nIzxESvC9r4q1N2SXrYazZj1dpXuYM6Mw
vkL7tf6z4VOzuaQUZRPx8akooXfAIfntVlPFuXIOWOcVQsE269o8dSMYz1nIsG6z
9tA3SOa0lhrgovie3gcewtieHr/JyL8V2zCB3+d/er3BAJrO54+AYWXaE5CZcQ7t
Z2SK16OGr+6bkMkUYCpj3cV2ODGmsCIAXP8lTW4aBeTDHGoQ1gd0bNiAqKDthE1w
IwKT/WUInMuTT/aGW0m5n5vUBv9P4tB+ZCDcDK/rI1/MiiW1DBPXma0lwVBNSS2h
9jTHyHGrJRNo/l15RmsxKOf/eBMJeLxPxdGZsQ3i5R+h8V4UeDqT6hMqh5Xb2ty5
HRj1zkKIbyYK0heIgM+sFk8M4hnhrM8uXRPUFTivBeCysvLL0pJN9Cj0xjcwlkCI
rGtA+QrZM81ALv+Ggzgeqs47heMLOvdj2OOsGQJTsu11mwlsHFpjXXnvcwonkNIh
RPAh937UHkxsRoQkqiV3mrvbrKTGzjTjM53PFk4phsmnZX8PcIT9liGvLpZYPSlG
ceph97jC6x4EHFSgd56AxtMTHN7DvAKUGmBatDi4KgKeXTJJ2hZp1eNILljeT+oG
6YlixrN/KnBrJayIetnn/HnWnKGZUesk8J/XEnB47SV9an2+nNjAPDnUY+dGEmOg
TATRZW+KU5KDwqK2vN5hB3AR/bZQCwkFf8q7JpN8WzenWvp8NVpcFFr82TngnknS
pnd6tMmH7DyVTn8FsEmrMMUCKXjhNLZ6p3AZcTmi0mKSVfVYuUZTcGKKsrrx+mCh
rK7gPdEAk6xG6U9FhCeTflCBF/OOrG/kYG3/EHBSBzweFLDumzm1hgewsOKZaXgl
Uy9MXXKfpdqakBDyz65F1FyWmWzcsTXHLDcavy5gsDmiBn+ZOplpc1tCfmr6GFkV
faWcB9/HrBgYdF2OroZxxhj/qLqO/jM61W82FLo0AUN3WNrDgdMVlVjpz+2gVYzH
SM08MHcUu7wuFF4W7GC0ZZtefhKI2bMyd/1tSUWjhzAIsJiuh77C0+75eloJQIMu
bSdLcfCfCfqgj8ojkqAur105tDPfrmDDPbA7XKIYgu5GXRaKum7sW/M3YrZqE+2o
b5k64TI5hb0Ku9LKowhg12Ul0Z0gIuS/oxHT+TOwgssWSfYG2sWb25mo178WX2Vz
StXGJUKNrJIA7J5R7BJIN1KjkfpjVQHBZKMQNoOB5FTQVNOpmtcEpORY7bCt2cAF
og1aLDaF18IWyZEJ5WTsmvA6REeQPucwZ7kBoKGaYd6vKrM8MTFJU/4PSZqZG2tj
Oz89C7avYE+TTJaET44PiITLbTlXhwKYlRS5VKTojGY7nVcr8iIZEQQ/AOi29exm
bemrECt9R22D4LiO1rsigs4P1YSOk1LUlkfaQuYR4X6W5bF9eAm30wAq3YWz0D1X
cFO66Gu92roSxBd/slXH1jmBCXvRsawN8354UWHzStN96U35/eJlsrObYyL87i5Q
wJr5n4NGNoGNhPRI1go6v4KtDoO80RA9kHsb0FL6UjJCdqr7qgbU9GygL2wUziEf
ZdstCxnqtBoLRQc/zEgDdkRHeR+Wfgo1fxHwPcvL7pbZ0fhy2eA7doIQ0+xTRVKK
mEoxy0cFwBbQtzFh3/nyJewXrwQiEBrX4cokhcUjXwhgzz7mrMwaGOmTSL3jH02R
kko+3a3MhlZ7Qv0gXrX7+ZIMBvjpYqs5+PC4TrJIPVqiEJzW8aHolGjAxWTjbWOg
mG0CHGWjxWCy1cuT5SF+7xRAE3jPrZ5g83OQPXqxbeemM1nHmhD44JnFR0MkJV4C
NUtHL7ZBcGI94bI920zaJ2ZrnqA2JCQ9RiCV7EgSOPk7iZY+dCbXt82zPReBuWn8
ptH5x6iImEzJyMHOpZZXahrNtuT8+qzqU7e0pVTUB8Ty3lfyBYMKv7l0FSY44zaQ
3Hc4sWdGTnl1zdaff3Mvf5Beb1GpuqDDUAmtFbHSFLqWTyHK/2zfUBGABRXwc0jZ
cCgmiOnAAN+PL9kqXIGZf/4Do9ARZoU55h/mse+D4JBBUBpC/dSSoH9Xxk1upK4M
ScBd4ptlK+QPHEb+UQe8uA+m6VmGvNU7bMXh4A4Zoyc5eTFV7KaMcJ88V6qnP79r
gzB+35qXnyyQ6XNIglLN0B9fjO/gLoO7qEFX90IAEJzhsHA2vTeZQVMCtKUPLWZ2
kcHB46537js4r/w+WWyYBqAaUv+3fWN0ondDlddR9yIe1OjSv1i01qhl8nmsgiqv
sCWU6Y7kWHsMlr72UoBC3I/XBiYrtRtiSZHocvYLG4oNAd7q6W0fmbu/AZ81V+9z
98EmUflFhtJJzHf9qIkq7/k2IlAtaShPhz7dNvBxzynYwHI5gEcayAwc6iYQu8qG
fLmZNJ+DcvPkmEgNjnUwRODBHbn9gjIx2WkWmXt7HnefdK6q8nnr5FMbH6Pfg2YG
9q4rjCTAt+4cUKk5WK2tKZ6/nCwimSdNM0Xo1o1HLIlAA81g6nnimrld8p0xTXwL
OoEi8XLP5naXL1rr83AAiww/Ys7ZtkrwtjCkuxl4XIsuef5HNkaus3TK6bVXlavo
lzEN+bmOr+Adx1Q+gEfOI0JzEXABzBFf5w5imzupPfyy0PbjWcMuM9m5gciQLtYD
PQReku6gH7DggK+i+hpMK/GfMG/iKUt3/4X+559T1I4DHfJ4fO8ho8nrvTh61gHJ
rFMadXR/afq4mNZvX4CsJ3vr6vIJ6xBGT6lUeHdCOzdI/YLX5dRu3aHYNSndvL77
0zspbtguqMi614JeBMyIrgNyITFIDJRtM+tNzigYVMHQKiagT2HcBXlSxH0xuZD/
YU9BH5XbZw+N2gbOubmt3ju+ZbM65BB8GT3TV4hXXSDBtDTgqkfMpdcsyXNvyaA5
ToW7aFfYX7BqcCgAJgYEqGxoiZJSeRWUUJ0/AbSsoVEsH707TroxqyTkhRzh5UAQ
4mIh3FhYNHuhWNC8wxrzjlhmkqeFTXlkTonChXrRNeb2Xhcs+1npFU28DK6dsuNW
E9DxhQJhCNBjdh1FP+NBkMCdm1Py3x8smOeHGCAFq1aWuLBGpYKWKRYoq8ZvB3E0
FvBBEFJsCMjuvwb2dd1SsJbkzQONqBHRkBVX4+ZSgn+m30kNmzHyMiVA6/lVX/sr
zjQA6FW+lpXR4dgVzKVFuiZtkMfXfobPOIpVi6lvmwX2eju/+Z4EwJ7XHfqgqubN
4gMMr0gY/gen/GLUevGo3GgXW9B74+dkyXi2hn/stFoaaM2QNB+Hg/0hwK11edL3
zUS32v0SQcfOIdh/P3N8dorqOA6CO9hW52U//r0Gl+1PmnoNw9HxXy1d+7niNMXN
E37j7LWeNhVN+GFZ2eIMe4ThMq3Hn1qHDjhEcAsZL/iYvjhkjMX66HXsQmHU8Blp
TcAd7SpAPqPlo/+wVgFhpaeoFUir4UkTnjGZtf+/xxCtwSbVUTzsBb9EaH0fDNtm
opuxl6TwxF1FuadjR68QdfuwwG5h3SbJmxPW3pGSlwZOo/AoX6lnr5Zy88Gw/mBu
LKZjy5UJw32eSTv+Ug44gN1UZQn0AeZyyXSa9haor8TlCrTQ3G/YPDHOhC577YbY
EVDXr92Rhy2pQO4b8YYKyB+2zNaCOlLOVFTGc6VUoDilgI/yhsRReXUqyyk8O8y6
mqHNWFbioVSC6w3IX1p7boorTDrPEay5LA8En1KNWaNg52JwxSGXwR+pN41/VpLj
QpkFdx7jt1WPVEvgPYAkFisl2j4H+5opLKH56S8ukOkQz/uhjFsrOzSzOOcAcazr
/o+SktaBpTqjOyD0lhuzyj/+kk3Fc0fS9NuR3MK11sOu4+Qr3NvLgloltaDrLjcz
7Jfp406EQl92Dofg2g+eXDlldCRImJYTVESXv7YBjUW7zsCGF9MpSFXnDWE88qLV
lhvRV6skCASuq5qFbNctDrTlV61j6aV9rkEyX9r8/OdOeAb+CeAOGe/WSQBr4Myg
kVtDUBdztoEQDXkiUUv0M6v9z3ctGCmjOohSCvuHaXlyf1whdzBiyGrSOfr0xFy2
IDmPl6iEuz8POG7w+ycaENy4ypftUMsMY5TfX86fLmsyclBWe24BvW53owIBkuhs
3tLigaPqLKTCZxuCVoWRh/Ocz6Xlmjd2wq1hzrlWJhxtJFU9JHozm0yZqoujozp6
57PL3gqWBU7Qrm7EKCpHt8qkMy/+aeIiakcMHiD7OiaT7QnZSLyqAf0qwk7xawgo
tbSbCLgJ9SCzOVpCqYDK1QXmDvP0KdZl6CD8kTWXjWXHhbEc0xra7kwITtJUrB40
Us3gRroUfX835fI1ZkNNpqpIr4gjlL3TYv1pvgDtnwq7CAZkU8CV3vZY5oy5suhe
ZtcBEuTfiKJc0dMtP6DxkbTkA1+1UEgytTISPYT2sQxzeASUdLVKrP2zmEKFmrXY
V3b4jXsSpbWO0PPd3i6V7YhdEQVfJpkho9xZNpglNEuZtFi2H7v+080PyXoYV3Bb
DE5Ty5l6Vy860s4Ga7vEX73thk64EAUQW0XnT+33fvPL15O+RPSCM4nc3VDkIJHf
qwmz6caDRzbYNn9e9TTVQH5jlrePqiAYk2RHSjp/bv/s6MbaxDxGJSbSfZEiXLoq
azxhWX1jMv2k+uXi247p6D1ntkV3C6SclEL7M+h+PW4K3skAgs/HxMw41gblWTMv
Z4f3SsYuHj1IY4t0W4aQhTqc0EKOPj0sKphyljM2WuThl3rENKyv05zFzRn2UAAz
eeB5H0XyhWJsPM0AnxWxlMhtNsJPEHseBh2pwnjRe6hEd6g2UkPXtaWFhUlAGcm/
oDvsAaL50QEWvnZPES4yvakcf7C9HyxDoLOzhfDq4Ox1RGywPJ2Wn0eQLhj+ABAf
cPKQ6QXkp/ssbjKDUGL6St/3xPS1Tjfv82Y8YHAVXTHAlxj2r4xC4jjMFFv8k4NL
WikZ+753Zh4UWJdt82Fka4Dl4MMHEHdaTLOfNCcIluDV936ShUywI3b3kmxreumH
Pkcw53Ix5lNpncZVO3uGvJAxy/IbA2semOvjw+EdnmxINSu48keKG+Fx+MKy0dG2
0FuqJrx8a7XmLc0CM6ZCMZFuZh3m7+huhhkZN7XKsDVYiGCRQjGBDI5gx4edx/tM
7Xx3LAW+PRofk4RQ8oPKS6YdHiW+xBDZwLSKMR6PnEYrJYacmuoi0mJG9x9PqBl0
tlcPcZCBEIsJPBBBHokY2TFQnY7SnZ6d3PNdJqb17ItpFbgTisZMBUft94wpld1K
yZhCmBUtlGlzBUSauk3SULc4YxY+wOfK6cIUcvCjUPZnyz9mpQxjWy6IDL2mrrec
pCAk1BxABy01HRW+MSn/b6sAG4Ej8wVFRy5enBK+x9AGwBlBBAXmG831Ejo9BC4F
rfCy8PaEJuZv8m2broEqRfXHPcfqQWbCkgqb1falWhoHHbn5F5SYXW5OGQkWmvfr
Omk5EoT5PD/yvl8EenMRuo8UnvLX4WtX4hvW0XQ3LM5RR7rgfToA0E0oGlH7xZ20
Wl2DwW6YkpRp9X38kx+4x7HscPy+wt7513odPzT8FREMZ1D3aa7ZubcMCXD67S7K
pD4xhVoHCFtjCrpe42OLqIAb7XHcPM9zfNv+zSezkELNkBGHhOXwYCnFIkivvSdZ
HYvomsDx0tR7Rb15owQ/0zUHqn2etz2SQWHzDd4C6aOCA2vNXiOpyhTNWvOxLFZB
VwJ6KahqQ+GhwnLkzJC6/qWpq3oPB0yYX8BjmFYuvECBkFELr3qPEeCiAO0wzNlo
9cQ1LmpSa6QfFwf9akFIsLvM5lQMcQee7yjqTss4pyZYWLDsCH0UvrOS7/Joe3MC
7qBIGh0lH0PMS7FDrCDLVKbkMAhuKmKus91BFtiKLVywQSEMtGBSzg7iXqTlwbMa
JExCH4Zb5EoPOwf72s1jMohK/++Vcz2W07Efj6+GMoZbAmflI/Qmy05DaE1TSiru
T2p69CMYFJhvjG6BYpqyBVmQI8vHhU1x41KGy+HaeqAfKbNlKDTHJJEfSnK7pBxa
1UTJRBNl1roLfxnWNM03e3rEsruv1wWxSBjR2sojFRz2tCoUfa5oIJE7A2/6Dj+s
A1bJCImEEOgaSqherfEvcmgWe20XD3qBEmxN58YJaqyi9/mx0qIhjy9Wb4AQQ0JI
6bgDfzNi1k86M2F1K30rf+RO8XyXq18zO7v0HSfSyvgwxghei7aslpnIPe6XCV6n
0RjNmKTi0g1pqkBsRd3FNADmxSbUCJ28c2SNF0JE6L0i+k2NjRCZJODcKt5J8zfk
r7WdwMGHxDms9KBRHY9qGceCJtl1SMoS6ECtCkjMsULfH0aGZCJ44/l0zREywxHT
0D3LDUf559jHCabTDHRnOQLWpJswz9kpuuq1gL/daKw6Onrtt482ks24DVb7Ifdh
C1V3bA7AZrQG/drkDaROSohrWp3PIutMMLKcEDLVhgS0HwLxnzDO1UEgbAxsTd8A
1dLc8EHXmOqNCx3dteaur6GA8JGU8/hqozD37DYA26jatUwsTAsK4ISRcqyL2HR+
/7rUZadyJjMmkaqV5vIILBntPGrRN7OGhXLrKz/A+JKFK36s4PFMrsI1FSPc3tbL
0zq5PuAui/PCx15cqGHOxZbAobwqL00VqfuIxG3jGWoDDjHj91pmg1/c9d1HsRvV
ai6Ugahu52jYBk2dYvqEziFYQLDfblyWbtipeAJIFJ1EF3+ACL5XePqehrFsqAmL
pxO14eW+2DIT28cSEI6YFk8iRcR1TaG9St5xMxAfLGzOm9e80t4RTtWiz33wUKpe
RB8DhUdKigVKtzX5WWnY2dlVWWIAYLZxKG4F6x7fMvrNa6PzJjWFmAPNAHvFoWJZ
/7g9hRJfH1xo960vWkJo+2pF4oZKMpkbBz1zW7R2QKNIeaWVT2OfB61g9cIBgqcU
ujSamjKsHHrd/BIbqmSH2OE2wM14QjJ6ElCkmVqvI6FWye0aNOxIz//8pYNPa40G
apciK8OqgcykaUeocKq4ZmBULhDjn064dwq8X2BRN1ZA1fjXNJPqChR9E2pdV9+w
SPiDFJiIQAezOXOltlGnSuj9jX2WNFj1apd0c39E8s2hquIxFAXEdmtPSMsbjj9L
3GRlXkWuBqW/MjKciJb3aAdQqcODscBJu0J50g8ONejTlUt5/XoMailBN5zMFo86
HP4Ne1fbCEw5QetdeJqrf2rMILW8ZNM6nqdqHoIdKNFOOzCJtQrySdfhPnsdcef2
tpYf4Mgmm4k2F+8YkbzoHOOC8Q3JcJ2GAL0CnFH3AI2zK2oxIxoEjTbzOlFo5rO2
jBcysiE1UoPVKHrJuFYZHgvUjoJax2hHgqFsMjt1PfZkQzYrbL2nyxUV2ythkraT
VzRJPXDnco1foBps7ty4RHGRtmOd4TN1gFj+FfgeL6053TB32ecrNeyEqJquwQnN
BGK2wC1YX87LODvN1vAjCSYrfbKNrXd9w/5c5SrJ28m1RBs39sJ2VS6AQyaLInKc
ji/5meY6U8KU4tWcdEoDs3Y1eidBBFeuNQtNEe/kIpvF1UC4sY4gPBUaLAeDlpeN
Fo+hd5++t2RQv3cgZE7ZdrDkw+92RQnJ+f5CJBdAyJrIvLIGY/BsoeqkWuTdAA3L
LCNoK5Q+e45qgnNpb+hHuC1heA8vAnStaZkPJ1w1GL36aS4Gf1jLnI4v0qi/bNcL
Z4VJA6JhPWjO1x8bir/BpcG9hNLXXz1+HmVhA5RL7ZaRsM8irXZRFpqFbGloH2Uz
uOYB1+9IWRANHNKq4E5wRNB6qUAsEF817aQqdyz/w6KTs8Uq7HWzqa4ZcDGqnfcx
1dy2RX0ZXrQ8EZMjuqntISkTswwIN0GF3QdQ85m16A2ZuEpXuNfbk9kwtZReoUOk
xdV19+Ogc8ssJPGmsqobDPZ+tOT5AMr0Wb17pK7kIcRVN4AKF0DADbRaGLoT9YKj
/DRRWNAQP0o0lor+yWG6QJf3o9t2XgF20LdY+pX2xkq5WvYfywqQI6ONgSqrIBnq
sYVk4bzBJ8EuNUaneWDuEXoUzfEj12qKt1sgBStH0dEL8FzMiSIaAGnmhDzNTiKN
rgJMD7YwYA2KhsJs4kB8GdtBURyjh5zjFqlWxwlfOkdDqQvWvR1XPCeCD3riyWKp
F8levsdKOWI23NPKhbpxv4BPjREdvXpB6sECD8Uv4tcaBRkZAprOPm6Qpr4y4cAG
YNI9qnyaY0J8R4XYZFjMfAm6gxJEp+omZi7rgzhXL9hskppKsLua57Vibccv7lRh
fQBg1/97VCi/5vUEIEZ4xORAwKDZ19H5FZTcAsUfo0cSBV5dyekeczY7Mw6OdSGj
97Bh5HBi81gYv9umGddoild1GWxnV1BYbm31CFvFinK/Z/cqBHyqMNiWiDH842Pi
fABhYy2n3790rGRtJPqw9rKs9OYfab/aiGn25ZyYXGlP7R3efaX2QgXJnUU/0JRq
9zp6lBdRxsmhiiRMWIQMpcCtsCch6+7/gOgEUBDrtYfyv5rHf483I4cxTNmwrO7M
K7b3ZOeJ7z2BPVWf8+G2fFSNKSvP3vGe2duisbUBEKiabJgBf7tECCJH+setCzuB
9k8U0T6igA4Fr92fMb6RIsKcUrgDqr7yhE41dfHMhgl1GZgY97bnGq2uRLEeZzQJ
qMwFa2whVJGwPTC7yAovwYP/yl6qTI2SHYO2cjIWY6fAipIDwYVNpTITClmTgNxX
bruPhD3I92oG4SFj5h0PWgeF13Vi+tQjYA+hFVKDuOhf0kEjpzFAIBrr88DE4Epw
bNp1BQURu9ipMD93NFsY+uUknQEkSCzbQCEboDuAqCkVARdRqXcWm7eD9AfiMhEE
2znixhlZP+hyUxgRPJ5r7JBlf2KPEX93BmFF1OzyGnxKrak2tS0g2t95htBttbNs
tNb88Q3aos4nJv/d1/Uy3iKHznQxanycO+l1w/9Z697Iq2vXAqU5JJD7DJNtFGwS
ptjZu2iIr05s6WM0lQcXY6sG2EYDf+kfLer2hJ+iLWYb6t/6hFsPkM+yEWZ+N+XM
LebbO0IzGU3iLL0NFVpV0PpRIVYfmkoui6S39EMRhKfjykBoZETHg6uGGme1n0Zh
o24Edymq4hHEE5vnCXQhZLhvvozEPdcnI/DJUOmU6QPbnYmoRDB6wXFznFw1u1Ws
zAYTjC4HxgWxu6/HWCSKqn3pzG8sGVfsRPwMgNxRzkYeGX3griNI6a1zIozTFb3p
1TWsSs4CrfIHrlHc5cz6cnCFWAezkePQvlmIHk/FjjqLeZfMpZk8mEP1NhDcjBls
IoWURqHQK61GwudMlq6XTGxE+xm0TUWVGR/PSXX8dLJpDeEBURlNfmchE9RSa+nE
mupyzwomfAXlXOtbsie6GgTUB72dvdQOYU3MmadYpXq1gIMCKQqvJeHgIxM/pTfH
1k9aeAU388zsptmTMbdmrpPx56A4NjHffjbPhS58CQJKwkoi3Hn6rcELxQNrPSrY
+mLIsRBy5nMAjzatJWqKOSh4rAMANWDYl2Bqn8+zgZ1clp/NAdoG/1UGpqSlCOH2
iIdIaivnYRymGbyacSxZZ2u0sLaTGwhqeOYw7gxZd7oQRORVRnTIujVQ0s6w9H7n
m7MoRR/z04bgT/E/ypurGT1J172SkP1FjrGnJM/ZuFf/zgItAzOffDpfLNYKCs0K
qTVuZPfsCSNONlhF0w1SFYJ+VO+uK4xuRqgOENYpkdrnHekjChuoPqRu0cLwQFsi
JMNvNVtIjG86n8toYRNIeU0D+7QWQUreuGCWzSRyGZqE+jq0CJOzgWfTWgsoInh0
g3U734byBxxsui+1ozbsczU+ns4nqmpS5gP+w/mSQHkvvvRowmOkzwvg769tQfIg
LEWJ5eN3i6inUjy+W199xUcNlMq9+jVNAdADi/h+M9W7NQGaFNjckXZtJNsE1oHZ
d7M9G6A6H/rcojKDG/i3lrWibbU2HthqA/s1pUBrkfrEqn0l5++R6M0g0WorVI+x
JUwnU5iZgwahphdRtArxkcxLZR1rkenI5fnwVFoBbqXcG2gi8C0YGJ15GaD80nhy
s/sbtLU/8AYCi6pABjwbOHI23vOnkGJy2nZ7ScmDIfxbbmDbnmEexZEy0uWJLs4R
RrTFVXI8NnDD+xqgxyjlLKezNWGnQfX3cxmGLz9RroizIO2HoaJcaoVevnWQaM7J
Li6vA410II0u84CUCiQI/idEXG6s4zpmCbMAZj0EX9747VsGY4JPOilYmrjRMjmb
tyZKauDblnBvdmDxaEEgS4gbUkfoo+KZl5wTq2aTW/b+c4qWTdRexhdFW35yvGov
KvGeiBv6PFVtCB4l43qg40JoWuBsovAcUBptATK97i19nX5nubZflPa7UiU0NeXT
KYhBgcdGzy2gaIKP2mZlTxn3QnFasX07HYxoCw7BQ1rkeXOenjRfSlCidahbdg7m
/cvLIgz41SFMocmwoUpAQp0EhGnSOChAbiH9xEEh9UL5reAj9RD9n6IUKUnF3y1J
HKgvWxlCVpQMsaF1fhgxpX0E3huqgCp3btaQV/L8mDuQENLSV6BPzamch/Scma8s
Q6JnuyITXZR0X47PeRc0UOv5J0k2xHe9RNXJiPlaECR/vuY4fk300VSlk68D2W1Q
aIt1kN3cpIeUk9ET9L2yB00dUE0X+yW4GDgo3U451EAk9v46IUBsy3ysw7G6HRp3
He6ERm3+7v+L0gnLQODGGEhu/7aIRqZgSckmpPNfU2Ub9gl+3N4dNfmlny/i4Xwi
BaoThYIdYIUZNVFgTNyHznZW991WESDz20ThQ+oH/tLhI1yAx2eWFnVqXoLC3CAk
yALFVDcqxhsJ9gnXi3gpyORdos2QAMdpcd7GWNY8TMRIjuA7g5+cs3dh2kKKuQld
wF0V1dN77efxYsVodQBae6/2pD+q/DyjTlXYooDhXWUbjyxUJy1krnLt1Z3oablx
/3TJ6QJfiYrj34If1CH0DdQlEGTfqH5XBS1sLJJG3GQqAWl0Y7jhCuIALwqyaDiQ
qp0XB6aPX2x0KR3ABUMpJxx5s0R4VBW4uICwqm0ephQbsu3spifu9UYYhqoWavJQ
2MDpC8hUvrw5hwixmWpsACqySNP4IJ1mA2v0kpNkCtjNSwd27EBK0utxnVvvlcNj
Q18uyQxUDI+iKxuFFu+8OG9UZCR166EFMzj/nzgcN/o7/RkdUz1Rn/YzfhOMm+vb
7X7HQS94UztoUH6J0f8HTDv2yASnTCv0MpGMTb1gLNpQaEkApxsXkNC0ji0PPCue
56hJ+DXeXj+0oHJ3uWsNxmTC+dh9M3rOLL1drtqYVWCieZnwHIzGO0Y4cZkSktRu
0i9ZPL2GaQm5S7HNwToNR+176OI08cSYdwO5zcPcNB5nPRISxE9pa16F2W+WEe3C
6ezFoqHmyclRFcQNRoXqC6NQ5sD2Ee2OT3g4x6bTg/TVy1SN7L3vsWCbTW1LLpXi
pYFvnILAiv7vmZw4T/r2/LdO/mQwsax8itH1SwX5/aR2B/7XhAxV0L5/hhTgn1+N
1QqJC9w88uJfAAoHCgNArllqOPH6hN37t2mzk/dq6oDSYOa96FLeclQ+yVobSkaS
0EdJwwNCT4fkIZdwX59tgQruW6Rx3trjam1foWxOLfqavn17LxMYxRwm4B8YMC1+
4zCDyppMvJF46tDjEGYcJlgcm1IYaSfBS+4zXAS/5oz/t6XjjITQUi/xR5UFbDru
mQkRbARHmxWucp29cw317dWDEQIM5Bk9TqzVnIesbnAaxtQ/1xkngBes2kn2LNes
9FoWqwZvtOsVe0FumYy2XNIQZHcDoOLgezCZCh6cUiEBI3WAhXeI9yasH132C4uI
fSWE2HE4ExCUbOwZuIB/NEavxfh6XmsTg6KYTxy3fmwzk1v6inS9jPSGVgtZQ7+P
4aUVO0cbivIFpMQHrLcS/9odLD7F8/cC3vYWqzJIFi9liu//sbrUHPg823gIGc2n
eRgRYxLRbbMYREAm8lD5TAMp6pyps5ILs3D04aNMtVnnwMQ+dh7dCxMzcWv1TpdA
43XiTFDplD3W4seduMppreo0M/5kxvob2s1/b2Rc5sEM7H2iJSpmkuTaWcOjRRHR
3S2PFc1L2knXk2uOcq1Z4/1Egw/3+He444K3ZE2XDXEheGhHIwuJfXe3crBcUKdA
HX6pUtFY0ZzFpMsauB9QWOVx92nnovEWzp2CHz7emTUNNV5+Uu8rnIUFNOMib7EC
PvHYpYZZA44BDCJ6kOGauHWBWGj31l4MTycy8zlDteBTRBzYSLZv7/uHpBe17B+l
KoiLlvzCtiWpWpH8c2xR692p0iZBP9k9lE8/LuUl3+ZHaQVw952rvQwSZFwbQJh6
8VkLsYSRleqPdC5xK0DUaA4eayQO8auumQjzI+7oOo+81nFvz6te99uFUx66WCKr
oO5J6m1ESrGli7RU4Tt8tKuJHvhthLinAIr+EHhWMASZJjeHSM4n5Ud7/qBt2AUW
ZZ2Aaem6HueblLpHLp9n0bWFwOUiVfz8WcNneRcGExuwSjgugVyp+3WmurbRTCNm
SfKEMDggUPKIUM08GnRtD4fn6GJp02zMxulpkQTtns+86rKQchQOzMzt+ado+A/R
Sye8JDnoFwrJWIOLZWwp5nY3RU2w/h/sJSpd/RBQOrJnKvUc8COdROjBo7tvgYlO
xl5SRM1NoxrmgGshM6d0xLmvIO+yzr077XRuniu0SEEF+tJHYmyDeUbL1J2cxYaV
Zw+Li4CLA+AuKe+CEsfi30SS5UyL2tcCTN3gmCg6HcuABIBZRl8kfRZnInKEfB1E
uVAVZV99QebUk7qOabJrn83EDvCtTYw4Hpoy9wiTOsGIn+gR/2RCnPHjZc6rUJpI
+ambucfSZofvUSltEPs5oMI574GYNztJATbmRQXdYHrMykSENQZ+WTDMn1EvLAt7
LJfjhQIRUgdwHLCsp+rhjo4dqxSjzz39AneUYNH6xHFjnEAtbZVw/qw0QueGJqPI
ix8HkRnMBtqeHySWWFzRshO5cu6tAtiwPOFpGEVA+mlRxuev9olNqeMD6anNkSRW
eaXjLQa9wtw8GXCHuMqMytxkl/xr1+d4i5FvNlctehNSd/y1Q2A9u4TmfDg/BxlE
QlCN8k+2bpUSo/dkpgBluDGeTR/j3kxqpZI9RzSqUNRsIGC1Iy/qTyKL4QAepKRu
3ppQf4zP2XwJQJLI/XUg3Mf5NJ0svOY67f6bN7ZyRoUF2EuUxeajikjyGkdu8BKQ
d9pN6SXQZH1ryCfcCx0XR8M+VPNtznq7eMYPJS+pafSMhQFPuOVGPkNpUnk/0m4M
IV21p09JNguJ+Y1LLB/fMC23TeAmenIFnlXpuHq9RdgIdmph6WicCIpoLqiqFw5q
3SYyOmlwpn3y5+IAeaBi+MFyLco1FFph3eKaeMyBPK1yjhET3m5ZMwKIoSEj76Yg
yZnZ2ETn9RJxmea+9W6q5QWTDpVN4ZpsPFZ+lpDKu+niZoyJJvtsl3GH9Z9ia+/r
fXD5G40dgaInBCsCIj2EaIfNj6ELiQ6wRud8a7khGG5lvFUhwbKOoQAmoCp9ICh+
4IAIt8Ow9tP1hfQAmSeP8IJqfodIxNVNjns2GNtsqTPRJCn3yN36QDWPnMsuMgw2
FZQvpVf0KA8FxQPU58CMoPLxwRw06TZWrZqhNyTmjY75eoJ56iLnhu9a0FdCST8/
KqAlyYCyFKfQFaxMJdue76lMXnEa+zSGjMh8IGE4it1/y4TEV+GKHXoEYgiTAI78
IgfArsRD3gAZsyN28T+H/WdM8cGwCiLQwTXWT6o9KNWfoMCz6goyNX+uo+4v0+i1
iGwwyCpMc5IChvKFZn4BVX40bo8qrR0215KQbuDfZf+zZiiHlFXplxX4qG1mJoEC
ty5EFBeYYWh1gesqaQYEIs93HIJkrt8suDJTVNqwPx/Jw8YkLH8SkFSBqu6u6S75
KHEpBo5FFiTo5QM4Dk+VBOBa+kZXlAGyY+jcHYqyaBWkrr4VPdxQvVKBT56rIiDn
2ajBggBpdfZwyjEE5j9Lr+DEr2wt5akBkuWwA52Iq5Bn/stvcM7rCn1PF7ujSz/d
H9mmrDWjw/lYWF9LGEbxhKZu0Z3sbOr6owQQiItADUSoNMs/NXYHTb4nWer4CQtL
b4Fo3O4vrgJJmcG0ynnUeHfGsQgfBSKKn+Jj600rYKfdY8p4KFtAZhKhjmiVcyTF
W6Igf1cBkybnW2xK+PnFYHYarb1l6cjzn+AMTZN/8hiGhDWXaesCYatk9zC5quGG
8eK67Z0CwaY0Ss65IQTfZj3S8PMxrpnzB5OdjTHKcJ4V1NvOHYKgBPbIyI3KzvOr
4+vSTHLu1VWqE3g8VuYFQdWm2Gd5SiqeVg3v06hC/VB8vljOmBRr63qQLpGg9HzG
eqO++YhgUGp3mQXlgWfNtZjSVtN9TEDCp1VhIpjSnEpnlwhaXtBuW5kbE1yohKdO
uZMrIANyGsxROFmp2zqP6lliMqH9545V+SRF2NjJsqRDW7TbEw2ItHmbDjeJdZIk
uTaBG6hJ+4ubY6J9PTw2qB7EHAghce6VgqFTzaX9zyWy6FkamDhKLqJpzH10rYnE
aF0dmshpXnp7ccT3QXyB/7+nosy6Fw2IF3ChKAb7XFyd/9/+rqvLIe5Nm4BRTrID
AqwVypx+JWdFDIhCXf6xyi/kIG2spr2TlAdRRcstTDRc80Gefzt/EiyJYyjfj7aO
KbNBKTcXcl30Qvp76vz7GVamfSVFDtqhzrebXBdzPVDYCRXHTmpj3lJifXQE7Uw9
NOFyKbq/XfenSbhBmIuaggcJTcvIlybQQSyLmrm0modOFypK/jWZSMiFbMsTjjHi
CBjHf4d4sCtxEaHKqgVprvx19pQAKjNFvC6JlyCRNwM1FprNOWezDVf+ED/Y45E3
ZamkKHFokqv5hhwdBdnj8Y5I10YRWs58JicNdhSeS9pBR+RIxy6mTWIMIASvgAsQ
aSw95PSgHk3o+ZfU0kSnaS2EhUwHm5clCfSbycE7pCUrSyKQc+MHBtYsHlfssw5U
PcHFA3aEHERflvj+YfosUTEtKvQB6+IVZZ/9ZA1fjW1F1AIkj3CfJhuQArReKEe3
sQ8Zw37snjBD8fVkl9X6m/G/TGv4Up7CQfx6ndPOQTy9RpRhwpyLc/wlrG0dHCvD
lVU6Eu40plFVXBaFTscn1cAn10xkIwbMSD7GLbAlNewUbg/ns2H2bCPvJ9AFAsHK
EefxPThSi6MBGF1rXlL6SgYQm5799tFJ7+5pTMNbPmyCIBIIrDnD3vLM+cVTV05F
dKVT+mn9/8NnI/aINPku6KnDpkoxT0qyqeKrBaKRZMDJeDtjw0nQrJk3e5xEeHWl
7ZEsdRapoZava4N2Oue9krEZQT6JhNoEahBAcjS4elCejrwZjsPLy6n3SxTXZgtl
s1jgz0lctoadDc60kEXyV5jcY9Jwlm/0ZjRtWQAofSDSj6F/niVigYbYOufnBtfV
51hqBrNNIF5/u6Jf733azF3gTFWQWHvaMPF9ynkx8tqU9wWh9ZcPBgzj6xgBCY3t
eZOKiGTnc/EfBO0RjUaziNd4ZIvTkl+5EVK79XmAAyvkNiK77ps2CuQwLv0LqU8G
crngkv950SxmQU7YKFWTQfe8CYXK4AvnG4mWiA3Vmm4jyuKVLROKRoBjZLEDcjPw
hV8GaIXdHjuJ4jhKWBM+N401G5hguDucTWCkJ//Jb9VMJB0+xUZOM9yezo0CV2h3
NA6l+8I/p1u+Mr/FAxw7fT5Nv3WFGbYJ83edGuusWkvLzl3p7mc2MUfcIgW7vnA5
4GYw493uCPJ5gLYA3e720+rYF3CSFkgYwoIDTlHBC5eLnyPPZVwNuu8wYKfBNsPl
mmKmA87SZxXBTGbCws8iVLg8cZwo9b0PV0bPA98nxLijalnToln6C/wntdUB0jEW
HNi/F8PCeElH6AAjppCgx8eY83zoBpna+97ADTLL/ldSlbRIjeB6H29hYWQ7qTo8
zwbc6PT8kfZd//J+pjRpXSb1cejw9KSS46k2forHtAFwWD9nuPfTRy4NcAU/eNCW
nLYR1Hdb1RthhSj/lNopFoWaV5OXsCSk4k0MCmjJaVBkUsBCinfET7mTGwBLJUMJ
rhPnLb326n0PLC+9eQNVVoLZDVNiGKZV4IxeaLnhZxniVEd2yEoI+Ef4n5wop5Mr
4m6NCm9EX5Ux9x+5Jk3MkLtUNQHfdcvL3L7rR8Id/QlrIBIpICMUJhzcF6vclY68
DmD9gLdI6yodPBk6iyM0pIhvBIYAtglw7dl0ndgauZgBb6en5nVmK+N8EFaq1WXw
0gVL4degvuN4+5gA3IPE6hTSnj52vYlf4vIvMZbxztbNVT0KErcAb+P9/Xhw8Awa
2wufGtA4Zu1DnNhjPm03/StExD7Ms3PSDXpaX/ez1BVClLanxYCRH/olp+ydZ68g
5JRA8MyRdqAapzBLL7FZTMkDskMTctwS4TV6hdtkUJiLL9Uuo3jgmTo0EZNUnaSb
3NAG91uOEukJ124sE0GMVu8FiX/vNJMMYmuWn3VEC0vvtlxhRvZVODSyLjJlSa9m
NoS4U7Wm3aYVhXlE1Ul+Y8+VC6tZv/CNBVpY446o1BIYpBzVWkfYbG5q3cNlqNip
6fJVj24gs9u2m2ESxa6QQ0CFoiexrvs4yhH+9nkFYu1ALcBPQ+oJuJt76pYqwHAn
VM5D/BQs+mnExVkddz+wCSwPPWNAXirqA+4tf8iTgI4hBeaXMz1OvgTjwPVVCyXL
K+75zYzqO/Sg6s9wwxdHH3OsIDfLkjrzm5Z4pQcLJb7p7BAvM/N+MnQ2Ei4MG5LL
ka1spmf1BwZbtBd69h5WEMNk01oMxwS5yh8KbHxEPnMWvjr06h1iCEmiBSXILzK+
GqmxOfW0l7T4XGummD17xfrIl8JDk3ABQ53F2I/enNig/bmOPPHZwUCQz4XUdfgQ
YHWkHqjnfc4PJKaV0EIUJie/SCfLgYlHAK+n7kAFJKXScEWD450OpkHWIy+G7PjH
0zmxLbxxT4J9GDIjeboljq1JxhN4lxmvsSkm16LE0pAcu7zzGsh9/0tHEmddGb92
VH8JlX8zR6t9CoLwwWvUwh6pDaVbOoxdkkEi/fP/R/Mo7OdbIRx6GFbjGc5dhG3m
KaELXjTF0TOdQADPxi2cY6vGfvmdbd/CYcIezsQ5jqV0dWca4hlyB3/nr7r1DVM5
fl657C1JXETMjcpzxMJVftwOc8vRubIxZbaj3uyEq8L+KAY0nFzSvuGgLkn9LpLq
ZMomcVarjpZfgKB+abNAtvPS2+YnroGgtu2JF7VOu4gwalbs3mT1Sj1PqZ3YITBG
zSYgm3Zr81XAXEGWw26BEZzfEIr7ZZwLLgi5s1a/FeexghLZuIB1XpcVdSQiUHMD
NBolnrw/eVYBONgbcwRJ2JpZkAY7CyDNbY8fACq5kqXe6Iwus12Lg8ANw0rF2kSn
qyG7NVpmXnPJ1rdl5qK7I3KTFgpSfKrghoeNQ/2L0schaLtxxks1wTiaprkoiS+t
rWsQJw4B6duNYTRcBt9Y761mT7y3WBftZqTOIfS3fS1GBdp+qpnbipDQbZtesN38
zO3GyUvpq7Zx166DmEWbA0Y4OOAXGw1toCIcWWIio1XanlyKcd6nJ10p5N9yTgH8
wwmv2AlcKd1PILnd8NV4pFfkALe2ZyYBaX98YOLrLQSGA4rqPyUfyqkqegDbyvVq
YpjME0rppymamGFTnp1YvVRWkH79FFcvTUho0BXZU19Pikh/6Jdn7gampiZa6cjY
Irhdig9mIHQ1SXBRAGhO25O1N3+Fnc3he01RRVhPR2XZLYtlRlCHNR36HXFKAz99
qnD02DrZi9+e7uOih+PBeC12e67Af1nQiA5LFRTJkWa3DljOhRmna6ZEL+QTbXtb
xv1TLMO5FoyxE3zoRylyRmkhJtGo30B0I5zjfqnE/K/HNV8ZVqGaHQoAdS0Un3Hg
ey/aWEjE49MzR5BQ7I0LiUGbNajm0J8SAFvr5LmSjYNoLKsQiwXT+bzrhqj98I5p
jxCNb8Gqx80eJN9j5met0HDCYUDDTHqDYgLd50aHLPvcTddbeu1/LS3t5+WTqAb+
fhzX98rnrTbAgxrZZiH+HYbvHsV2Tp0jW4Zl7Hr2aUOWGYpD4+DtrGkdpBe25S62
6FvWSOSyPxIhnOKaSj40IEMhM+7rRyWTAwY+qKsiQjZszdH7oRAhz1f8kWV3jR4P
LK21xdnHdBvlP3EgCJwa9RZ7pgOjC+ezYoSpGTVqP7Ekf/XRp4MGZDuRu9Zt5TfG
L5fv4NHXd53Sfxf3g3TgLHWMJdZfWMKjqTvr4B2+RZU8nvQocGqe9rgv/7pSOXPk
0WSlRlp7NZ+ip1L11KzKhXgsPIuXpZ8+Gu+nfTNKF9eaoXVEvfYs6dknTHswv832
iwlA6RaWESyZilemf1cLXpycWHA0/0YI72cAP7Aj45XZxcjJhAtnUEUtcENo2vt7
d4PoT6HjMDtkXzQHLvb0gMR53MWnmCh1TshaTVh2O5ym0V9jOrn4IAGYUS31YrRm
gIPLE63hHnmNfAXMbk5niRkNB9UYEiygsnjweu5b9LYOjn8em+6CozfZNz9ETO09
pPKjTa9xfRzwLGKqJ6j8BjUlwxCePbPy50Gz62UQLRB5Eh/SGwJ8ZhfWwtRzTQZ1
uFXBAq+v1v7gx960KrNYcgVM6Zburx9PvfIGgn0rKfKnS0IMbC02hOGMS6LXBqyy
n4UarqsZ3/NZ1yxIz+G3T5J3DOZAf2gNHBQ2+vbuSmBmkUJrFOMIgbt7FZ/9o0QG
I3ArDS5Fyh+GkFv0dVbROeKxF+umcvTegzuZySw5U2CHqlwiql1qnuD3+cdLn6sk
HVx9Yqye0w+FZoi4ViIk0fH+E3+jN/0PLKp53tVjc9fS7XyX+AUA8D0V2TVHFBo1
BH2WSHvx0MRAb4k5YgHR87C7+RQzwBtRPcYfXvk98D1tEllA7Cy3UIWMFXHBF6qA
lp1NNE/sQSHq5Besg2dlVhOY7Ua+zYJLlO91lfk15YQLcPXC/x/JCzlG2827bqR+
RwK7lZCPfpLufJvFsXjdiLK7gA4vNPcZNuILCVjA0BeCNIHwm3WV8ufkmAYFbgkp
iTVt5JZm59CsgEnIXrJWh4So1kn9+omq1e1nv1Qmx8Y8+iKNzN/dt4jfWacE6uwx
QjcwR6wO0ydyymxF6f5fViLEkgI5+84oLJ0DM/fWlzepwxSdZOmiHMt1iI3FCYBh
CblnMz1I7mjJ66r5YtvnQzpfZ7i8kYUJ4vA9eDrJciSwgPbI5bTGXp84XjECGYF1
BGSPVALyZxu7KsjYpmTKJopapuiqj1idQbBPlh2DQK4Cxrf4QYyIifXe0syNCpym
cIJaGRQxIXJyVwfcYer8BKihQFp7Vl48twW3X72L/CrI43YiV593MvSSHMDFiB4K
V7/cURs0DmDKayNSKp1P3N/gNJaf1fkQaexlXArQkDdFcyXM7g3g7N/jt9gQAoim
zrX3SbLexdNV2uQafPPTVfDDDDj3sAKmY1SNU2BNvcwLA1tRGAzAFnsSaeQeMLtP
RAsWZqbQR68/AX0hSDxTskh4HwhHiWau67ThQpPn4gXvkRzFIdXVxyXFQarx91Q3
CTxWbTGvZmoyXS2R++joW4qFpmNkdvZV+UegltZJcO1EO0LTwJDiTcwqJtLO83+q
Pv3cd82I25T4YYKXxdFAsZO/Orloij3ZThWCc04IW1JPfWKAsqdu2Zp2Zl3klBz8
lFpago78iqI6be3uj00tWTeyIv4CDvDc5Agt0UlmFXxqhkhZRFqJVH469Hhwrp8A
XSBgGJPK9ZBLgxx1ACuSvEtiPUI82+UXNPsHgshh53kK8CyAgrVEtQFd7QsOkCnS
wWpTBkJsndki+Fj5njoP+rghtgyam2KJj8E2zPWL1mb4NHCEBK2ZfuWS8nzi8OPN
e2awaJU10SOUHdEOfygdzi5cG0UxKHbDBhdEpTuuxEs2PNG1IQBim32Jpne20fkS
j6Y9r4ES/18ay3cL8a09Y4uvQ3FLkFMzqecwU2pavMYKYLAgJvmPqMRG9u7QvpC3
GjJ1elzvVn+mh+OC3x1CmmbaqQnomzbYY8HMDDsDb829DuMaY39DeVY+BThvGDxM
Sb4QcNMJImkQz4sjs+LppJlTpJhix27bMrYtnJIdm4+bmpVTCJl0vtUUN/KsjBYU
x+vPVw9Pxngzle+g0WXyCr+orgeFaXRrupMHZiSsUpuvQ0LyeAJ0PAOztchb6n+g
Ri8W8TtFAeII7ZN5tZeh6y0sCfHKm+DIuwxQTwmwsoq2aQgP+ypp54eSphRlt40+
BXMTAVYdefnGsIMRNOR91wEBL/F81d4JAEZIzbUOjadv8qtcMXQcEhp8DN9lKyFc
s7ZMZv7d3XVkqVzRZPYV4xxUQ6x/CYSMYIu+vKG8HRaFvI/SoqowOafqCoFqPTrY
US0xaKyY1HAgX20OgklRmgrQRf4dp1vBiBmEnwkoQEEs0GMebrzRwivxXhhFRIZC
sYoWhjNHRP9E2EPVfg0XX1Bh9aadcB5RGnLclMdtJCQKBHclSUwCPgfzmDTzTkJB
zVHPVM3vHUwBsYln9HowEGkD4zFf9RFBvP+G477UElT/topKHgqfeys8zrrpbz1g
kU0OYxGAB4nmYhg0X+BYiZJc5MCS0+nqlhM5AHUBm4IAvbJmyP2ioI5ftY3Ojm6G
uocKtSgxAi1gwuxUYqWIoKpOZN/uYfhsy2Z47l2vtf7v3NPCn4YqMEqimvo/GJR5
bxGMjNg7SltCEBvnRfp6BQKEsJOLHipSHPlbNWtSmUaffJb4Pp77/9H0Psop9SlV
YCLRKlgeRymDRfKy6jbkS6hcKMLYgFgftZ9kp9x7jsu1YDxXfkeOTiRICfdvXNpq
Giw+FvDb5ebFpkQppLoEPVYQHeOQG3HjazmmgNZLN52pYLbT44/UO94mI391FKSw
4YQWlRuJeWNnut8j3gskI7bc4j8Du1wGfy34ZmUj2CeFj+QlSzUY/KrVBENnnWz4
PdHixewRuhk+XPk9DvC4uYBSyK6FUp981IOhRDcMMwIqtsd7fExRLvs+XC//2UzM
wwFtpxFD88T0rZ4szT5ktSbdVWfCtRN9Lu9D59lhVQcowDInbEO4nlVEefYoBMbr
GM6fDjTmnFSvtrDvh8ychRna4NorGAIw7WAgiI3h9+ucFMQO3VcBTHnlVleOE3pl
MzL7Gd3mcaZ4Sga4wSUt3pTl0iWmgVH9m9Nq4QqN3WGyQbydsJppWI5fAB2bty+N
kqKF6qBx+iGGxs+Kjf4KbZ4gkG5x/V3NqKiFx2DCa/e6ko+qibWaIrchVRYEaK4S
+kSI21eBl4XqgSxvJFOU9AMqqO5eYAuRmekHbOWqb6A5TXvbN29M2FPWZHgFEqnv
Z9+JWKzVMflgEfM3sfVPdehRIFnKiNpHZ2DIv6XvpA3/qIXYm71t0u3tU/0m+Zlq
C5oxkrLaxICCUiVhinUCRZirvBi/fubR9IUcFQWorSj99QAE/hfJ6n3k0y4xshzn
gRwTOozE4e2lvsb8nAfHlGlbA+lQ452hnQ8lnH9p6kRCMPS+SzWPkB5O6NIffa2a
9WSblwfHRevckYxzqfoZ230HYzTmoei1b5SqkHxoG4zRQjrcQoJ9+zkwzliu9SJE
lx17qrUJClLkwx7JGG5pX+bLED2+FXWALpWVhAiIAkDEeHTczQZQpPHMbB3ZwZgn
h0NAADyadooo1lXq37+k7lSjTftQk9vgOjmQ6mTPkZEaJrY7xb+S/fmYRouNquz9
AnXiFYJCp0sIffBBmHFggQDouSCWjs3zYTDTqvAzfuRPxLpHEyTJKqiwZvjlIuEE
xUKMpUQ99O7rUsXjToTf2OU+MQpGjMIJ862TtqLYP1+cMOjfAAcD6bQIuKgmXXij
TllASa9GjA857Nxwa8Xc73Nz/tl3u9VCMr2zYYVpMwmW4z6Z09xa/7JaAQ5FnB1l
1WdtFxZ8i8AenQ8yNgv9oDmsOU+Psx44YguH+pbJviaIqLgur4ph3rad2raGROmM
bB7bGVNsLCEabrgZjOPPjjFhGFrGU33GXUw7+z1o1CBHV/5VXQDcNMMSPhWFfI7w
nS60OC+v/jsKP+sAs5R7rI9mnHLx5tFA8Zz18rHf4leqreTg8O9cfQDP8KmOwW3h
/7NEa3YQ9Ybg2N8RiEvsLr6EN2nfjZU/5UP4a2xa5DwimTPaRzGAKqvFNQBV7Y0A
frnmUVb2/XxWDgJl8X/Xq9T4Cj67Mw53LPfvTns7mwVAh3lexZEUHWq4oWyoswn/
wkJ4PheZf9GDqNfPCn5Peuh09s4smlqlaW1hqxESzWUpwGtYMyRmgq+hyEwblico
KLGaROeG7nkOU86TQ7yfYnQQmdtf2tV5YGW48ofCzobZdz+OFDtmL68WrV8CjAw5
SMhFfjGZyiPXCCfs3U+OP6h5HHzYnpO+Y2M60SU0C4cdi5X6vnjUgGCmWGGHM4yu
1zkwqSSagSB/G6xHfTSjBUOXjY90MRgbxl7N544qV9ci6wiqWC+MWQDV0Jo/fs9r
heXfEWDWSObX4B4fd1EUi6KDTDCzWzCg0utAMAJv+prUUtp4qGtV8JfZr1Y+5CvJ
xMGguPT7dRh0z6+OmHaqyH8t1jCbjfIamCUDolveg/ZSv1seVmogrsGTMXe4fxch
KT0ZwNQpU2kbZEnwfyyNgR1TRDbox3+w6xUhqGtbDdI4Tg/JgCEIBL7tx0O4QvBC
m8i5weAXlER3vN8Jc2dAujWtgZ8v0Qc0gSTf9h3v4BYTIeT0hAfEceQ27FY5rTR9
u9tkcDt4qpWzpAw4TY3DJvmYuJqCiWT+Z3XfyObnx9d9fmzAnSc9U0k6J0favjWd
UXyvM5Q5X/pdL8tQY4GHWEl5oWDqTwwx0rC6eqjC23egSe1g/U8Q4Gyrjoqdt3m1
3di8jCMfWAC94x4ki20+RIr78lvRLeUqzO/ThzG2h87WjIWbXd0DkKoPkqeAUQbM
zkHYA/yx0BFNMKjS3g/bHDuypucJ6sbZK4SdQt4FEnTOOrko4JgCc4AyKQLfpJL1
4jvZSBHBSxiPyP8J4eCqLGtRRkLtN2IdBvl/KbN/PWZyc0ErD7Yb5Odwf9VSvbC0
bwXnzwpKNj/Dsu+HweDyJX2DrunLNeXdbVjSl0jG/EWriZD5K/WJhx3iIVas9Vpz
bvX/mIv+JIfU9tFlCwAqZmjVSNJF3CcM3mXkSi11sY265sGy9uJBAuDVNp5HK/43
VTGy15eXopc1Wv7uDHmL0K/j6uh2iKYIh3RbKtw4Fs3j+qNx1/M6C1+rplG57j5i
f1w5QdhbiDDOwHBxo4ztxtYL0N3cXdnfFfkedCn5DrK1EZcomLV5HHAlnclV2EcO
qIpq1VWKQf6xfIUB/e6eWwQBnjVRLQle+RmrH1dLvZJMM4cKcGqSi0MKer6na3an
R56pYtCIQJb2QdU2tx3hFd5Rds6OmxZSo4DW4APLSnIix1cU/nUTR1Q+NupSlrWF
jzU7U2+tWlDVUdvKoTP9FsbVsVWVbUAx7kSpmw+0W7Yf9CEBDpvOLxBWZ+YFbHh2
wmzD47FBGNQFC5ogHG0Zf5u8PdsBBqQKdOLn5oad2SrT/aYZ7k4V9ar3kOOXKuH8
6cnlW6QjrY+u8ebGC/N4Rdk6fByKfNRxCxyvNZIuvKBLM1RDnDZ+7z+D+UvXAhtq
Weq7gTliylFdK/J4HYLDuo0xwaG00kUmf0xCSEDKKJIlGFgxUdaUYgxH85zl1OCe
WKLlec21EEZw6Bf8okoF9Lx5m7zg2z/l6GUQO+fzIfU7mdWs7alnKhyBuAoa/dCy
gHDtcAygWDMUR06lh3hkZYhRGOUDbg3xTRI798wJZ5iyxDfR+o2DFOl1a/7A5Blg
6Gnp2uRZXoy3lPM21/iMFKaf2ZVgQmRmXzhUDpNtXcuaJ35bxGMBVwMnMdnzeazW
MjhlivwlL6CiYHawOfjBGvJVhf49kilq1OS87nFzoBi5SdXqBJakew41Y5+ckw9q
TaVIFhFBzzUyzwMZHNO07EKXhzvfw+JrV7LNA2ua3jl5uQuvejKkfgJKEw5nDg61
11PWXywcu5ZWhA4aFhPnC35YAHNo4NXLRiB/uiRVoPTRxSytlRMapVtp6RzHk7uX
J08eONI7x9efqA0SiyZHnGz3FM78SsjCENfWsn0a1Q6MBQkrrPM7FlM2SYR4Yj+e
oz9TW7FnGaZqpZz6is7Y/Q/H9BW0THt9Zf1UueW8tkjLshyU7/iiXCC8jjWKrrTj
D6TuZwv9Zs8whF2ddc0VlYvNXa+s3FCh14LFWX/Jg453/Bfk7iileC4CEQW6l0JV
LQkN/C7X44DF79ux5V+3K8WTszImXDwoYO5UMN2kmDDnC073KFBjywpC8yK+BLq4
73wKyBpfw6LgBUdYp6jcp3R0Vdb12nTHEKSabjm9vgZu5qckGUUF6xOg4WhBAO4C
JAL/cnTFdOtjY7ruJT6xIwN+56ZcLwAWrK/Q6sAEKvD7Nk4jKDXEAQ1j2R9O3MZ/
4/6IdPpsgriY9PIdQ92CTNkWR7kDXEMbtI3qX40Uotx/LZrgbIdn5Zne90lAoi7G
MJDjKremKMmuVvDREE8XkAAaES6JBztUqzAlF6b9FhrEKU/a7/9xvYHHWBCrT2eO
WnFgQEbL/waRZwVlUYQkVU/5y35axWYaKSLzs32STOOu+EX0lGP7DVfs4F30c5zT
b9cU+EllQP9WrU5eEZScPFdWk8eIJ23hToNJiOs+PaHr0ZnDhG9R3UJ3SG0wjTzj
bEJJYnceXeNCK8WUh8PP6tH8H1Vc0nkRyOXHziUpQFH8YmNecWcAQ7EuU4qy1rZU
Nv16mVYdEjVZuisbxTpbF5mBmQDclpJmnI4hBgl8LSAyB3A+mYhSDNOEyjPU/P6f
yWGV0XuCQU+j3lx2rHDTJwjFmK71XzDuzUZcDDgX0DTRLUrRdiXZ1zwmWwHhA/ou
aLSbbYWfQiMJAWdw9GEjsQoUUNQWM/CZaT9M7tNbIpujA8lMKQm9HckVMPduAkfo
ooVpxP0PhailHqSEmvXxyVvIS1YWWpm8a4GJsVkn44PvRluUifDV5SOYlVcUjAXO
OxtdLCQazDLBNxnybLTyVxQRWpIZoh6oo29pYLfsd+cIC+4muFJ7XIKb+ytOMi/N
l3GH0fQ0MYSUQuDQh6m+a/a/Fz4RdecUc/suwcGB20TppEPbjsckoMY95a5jeSBY
9QAThH85/TazXlX9wsYZgARUYIFzRy5tIqUtmi6/DxTOZnOu9D7+fSboo0/XB9tt
2+SZkoR8jN92NsUaGg5w21ixfYIex29RQQiNoQdu2EskSQAHPBNN7j5N+kW0ttRR
xMOofVLHffPtbhCDFAaMXWwwvB3R3YrNfDeIdce+Sk5o+1ESLAwdLkhUC5J35QNb
N8qcS+AcgeL3fdIvYpfE5NJeIA46yYjGpPoxWIoMyIrqDx8gwf/fe2c9sgIByORN
UDpuO56pdgckgGOcEacS4iWgHWSMd78KRzmBXE48tUcLN2c5uOYxx2RFh75muw6A
IZo3stlKjS87rbLco5IXLhrKpMNWfbTct5NBCwmdfbeJwYjD9WtoXKwdc+A7YLaf
Hn34NtRKH+JnaOBhxvrQBHNQP88Yb/c8MwE6oLqT470hOt5dqmAZuZxYHBClijDQ
WGATn1N15n8/4B+L5lHnZ7G02KPlJVaxJ6LmFUHow7bTW0VzAFEqBqpfOEK09T01
q/5YNsmtOqq5B5JZiaelKnbtgZF5DJAmL03qIJxugWarT5BdrHlnpXnaiNPbH61F
GhsO9NFm7PEXcMSsibvjGoOl4MJOwEwRjJpwEc20GmML3CZXT2HllwEF91+n3DjN
tsY1M/k5KVL9V2y/QT9/vU8cTN3owHKvz4wU+GXN0gLzj4VYDpdl0/xmgX0A6gyK
/Ld4gKfJ5vR4GUfH+DGaDqA4xiwuOOBDajAUt9BGg6LiC52nvdvilq7eWx1cLlzA
6JmL/otv5ti4TSahkZuQFqy5iT0mcw3NIauvq5nd9E1WputflCq9lMCmfhNqUzTZ
DLUlp83JyrMMt/AUn9gHhp+5UjzkuLo+wO0eEFT3WzRsaUc5YPpRmrM4SbYl8wAh
Olk51Esh6JjhFdBj6subfplEFznNE2HCn+Gc8OZCsAvdVfSFznAolWTkaiW7VL0w
w6A/NbbhvGZJ6vqgftX+sinGtzWXbWqBs0tACuJOpRvDnF8HmUMy/s3w3j9oMxqS
czMnU1nhiippZpbuuikvGP/5GUg62JvTF/Ob+ev1NDZ3ICtfxtpo1SMbaB4JyKO/
jO3SytjlY/QFaUUqlKviRJ/VLcmEBfY0EdGeXu80Vr2B5PpVEtcoNZQwGfRhJSb5
HJX8DLqaCJ+tojBQ/2ucURHnMUwmqXx5g4PutUyNKA7Y423up8AGk9brGzRPGCnM
WZqPDbynV+ShMIuBxumDDsJOmsOw5tKKWT8b2FD6Zzk+5Drt2gnrcfKyGEsU0gc9
g1yXZWs1tOPnuGXVdmYQaBE9HRaREFoICrlDaZyHd3P9XCxqK43vfyc5cqSbwWXD
1Df+P+fqU9OLWMOGITmUY/mpo6x7yjGNuzXBM4BfEFvWfeATYNRariDkd8qViRSV
1/tfervuNSNVsrN0KvRCUCbIv6Nctm/EcO4OdjQjBR6ZJBTzujzm58ks+TdsEYu/
zfPi0baWvbokGu+kYCQIku+4NoaBJtAZJc9gLqwPa17l7BrR4KZe7he2FFEGFLLK
vL9rjSbt+DkfpWFGZzfTs8tlkVqow2tEn2/ngEBcuhhqryPgP7myZ22qZzD4fNce
k3i6Uei3ZQg1vT97qOwYaacCXB8OrOyNO6iFU0rM+XTbKpcajnkM57jgTIp3cxmR
JVTxsSLK0JW/o3KUzTIhBzMCnw5Z+i6q0QLIGxRm5ecRg3fznWnL+W2Qr595It33
ZAKFtXQzJBhWEH2Z0jqk5j+VKZMhel3VqE0+0ix2YBMgk/OJ6XywoN+WWZ7i4uEI
x++EIsWlR5HYEnBC24HLA3nLgK1F4Zctsyg89Tnz9glAeR0R3JCAECsti1juVpdd
NEtvwzk1+Ln7cljPkLSMQFWBuNL0U0Sy59S986N23LQNcBbcaz2ncNiUsTyMxjoO
lFCHJDVnTDVTT+n8ug52pd1+jfUQmq0taMcR3gCbsfMu5bcYu5MA+ktJnJPWdRA/
8eabhqT38R/De3SYHS47qpL2J6h+ze4MYIewIf9t8okEzMdEhQ5dPFiIFu0SWCr7
v/+GMMUieu2NNOtyXIjEvelTZAdxsWQkfSIWMi3MuueCV+aVV9cTsTJ1QLjS3mp5
YJBK3TzBufU3pgr4fp6m+b3QJhIOWkcTM6ZUu4VHj1Bn1DJo1dprHtFEb4S1Dnv8
Fn1qMFdJ4momsHZzq7tTUnMYSYrkuSseSliCiIy8u8Xu+L8zkjnLOwwpWpc/upd6
2aJ2KQ3RliJ1pM8mjI95LKSDJY/YjZaOWi3UW4dlB4fmqphak2AmCyNsJrW6SSQs
apeA6OHVdslPhlx/aDS1GsVoVh1d0NhgU3hzphtQFVWj+QBbXd/6e4TO4htJo/km
KvgeEx0nSk7Gyzo04Im+LIOz9KSZexKOfIyHV0p0HD1InQ3WYfAvEvmZ4boKkJ9M
HBa3PV8T+vDq6P+iUsF+GWGKy2oaHXnBdXMusLwDnJlPWL8RwjgHeVuSQjDoBXO/
8UArJIK5T/TRNxUTlKWPgmM5kXzfaRuubRF40tGA1jCyQu8Yl+jr/ibuQPEMY0YV
jdP3WcbMlU+9EhYskv43VJIYG25OdwCtezs+h+pve+tzAHaK8roytj5MMU+4tIUy
TFxOmXsPCkH9GtPrjtrLz1YbCykwbUf5Wdpa+BOZIa4VlI7Telrb2qbuac8yy0Fp
vuyhamQR6gF6WB4wXRtZUJ0DdIoxDlpN2jv8f0gwoQzNGkXUOS5eUwB6UBvnulfJ
2Evda25lzBbDxu4vqmzrkcIA9DTtk/VCTQdRKxCArGhQlOi4M7IYPB2p2gifxI/6
ex7I+JWJ4lQ+k8r4Fpc3KX3uwS9UUP+83nVMZuEx/XS6blQ3yc852h/EaUIv4/Ec
pG3mQ3RRVx76ZnJiejukeJKbGy1BP9649MhuWSeB3EaMfd/baKRE1DBYpUmLS7Lb
WFROcUdfEovzynWzfpNAocCcKUnJZejHJSYEqoxDsYpavs1DsV8/oRMXf/YgF8qi
Q4Fziqn9Mj37L0gQ3yfgq+JXx/766WIN/oGJ+JZ0LzbmbhnpABGX8LY8SHGEmhKr
mpiWMW655MYHanDL33Jxx5zOSOW0EmIcvEkAmRLd+LceFBo3h5aOeCWXcu50HDi2
sJ+otMcvrtr3/FTzkMxktJnLUotC5XQXW88w0ZwPRRC1si+OUU6IscZTT/Q0j8sr
roOlzvDKqWyCvJYdOs6veOx+AWgq5JP4D7DB8F/e7FZYu0l/eUnmaQ/XzoiOWAJU
QSX9YgStw0cNze4mvDUKW0luzqAgzhgvdNTUSEZ95BCX0Vt43u2AhKIwRy1FLDFt
J29sbQJ/HRTY1h4MRoRUNjGqicsezgLba6qMJtb2VJXc2XpiVdtYLcX6/asOg56p
qbZH+E9N8fhOR9aouoaEq11SldeS17HxGvfEAdT3p/5tNyAotKZh5Yo36Xv8u2pG
vT+i7AL6AMdAwxiPTJqWTLjBtTbkOjtdnWhZu6uHw9oUZIDfnHfITOtjassVcdaJ
JC1dq2jndb7hbTBvBqLe9AWk/PUz8+iBBSrsvNX5W0uwN8s33uPKFzXGb3LehRGE
wpKveqU3EPpNoKSpfKfHaMadNbvDynr4rI/F3xgxx5UyWgp3cuodsvctGiu13JHl
dD8EwMhoOlvZoxpsU0Mn5OJRAQP62Hg1cIxSqMrSFqAuzG6dinJfutq1v0Tf8b7j
V60Lh9CXl8mFi6R9KppN+WYB5OkslmoPgHXAaew5pVcQxpLGf//FWMNjtkgPbeb1
Ao79K+7lmUBDzENOGCbbDFSYXIQZgTRxI7UD971RtOgfy8oFoyADaLKOxjBHYIeK
GKb0lRl8EwtHIKXD0hW+658/uBZXdQdLpi+aBK8ghsJDdACCaaLyQNOEk5x+t+zM
GkOJlz+C9EOh9NJKw6q04g55CpzUhMvtM64vwggyfCWLN+pFpW4x1aXMHPWRsH6K
qf/dY7avCZwNdrV18eM42XARfeSzTgaKm/wJRFscUMP8z/7sfSIfwi8mGVjzDt2s
UMpC6Y9f/w9KVHoiiO+tYUgdAyo4f+Mr3ymE4p9y9E4695FcI9N+u7Gz9rg11N2b
94+oIv3WSRi/cPjY4GcwKUIJP+4JuwPnAVgU5UGPnUVwf9oyzVKdnYjWbNpdgn6g
STwsEyOm+YBcqWDWky3OloohXidpydWtqtzapiSciLoTJyWth1Zuwt740GFOFekV
0ioe62KBMELscm3yz8y5jI/kVho8XehH249RieRPh9HlnyV02pdtJLb7XAaCc+s8
WheCtgNwW+4jIsuHPonamv+gLZR9opTclCaREMQ75SZiejX7+APHN2X4i49Ivy57
2L2z9/4SyUj75hyyRzZhKFUZyFUz86dy2WAx4pHKPdDu0gpcTSAiITNOfQPxSDOq
4Jqz2qskkiC/YWOBPWs8VPzhT4KNd5aHP5FQG1p5cQRMkSDO95rB4rjTnYq7Wi5U
juC2Ki3oGTFsxhLIBwofq4AgVZC757oQMlsQ3JybXgcqL7kvHnjUh+gJc9fOi9rl
Tx7viVLxCh1OGrRPm33dxkMoMvTpB7NLWJT0V39Vd+yAyCPKwgS84nK3ULA3FU98
ZVijz7N1OyJbkAq5PtDqFstVQtukKkskmzSIxYvTJMR9i4HtPAjMqHntIlX+PSvC
7aubjTpDHsfQoD3v1MO+qrGK++t/4B1lG6cSeq7r2c4TRTnfvP86ivJ4hKRU+VXd
ovlp5znFllkJW9vCRlVV295HwQPWCs8TKPphZ75j+y033G2SfCEwb0sFoYafFRMO
c6q8Hv4Bah/hoUfixUKrd+hv2EKM10YHHBhKZLjzjXxTbGbabL9Nz/0rErcKiwFw
HKIINL9Owh5pj73+2iKThSMH865jZhauSHkrU/fMyqaHPnJewXJbuOD0u1xandjX
nbtnq76BZFZ8tA4gKaNL8d9X82fO4l3uaz77J8ACpu70iVaFvup9pBvqibdPmusg
FeBE1cbb/2vFsZvqJjYDdfou1XHFScnTiln0OyIQVbHhPtjJ+usstgUHnfe0HmVj
cZh6fG8QxQ3oo7aVpHesDBg2OJ6f7VMIAjQvt1HoOJbrljU+o4fUsYKk7KhjCJhp
mhVbteaM43ga4vwQCJ5KEQ0tkiqKIJXkw9OzJFGR0Tb6mHFjSk7Lqz2uEkd00Vy5
maBCOJWDu9QvuPKt990yABfh0sXGwR12M/0igFD3/qP4242pTO9HS+XY9JgwfmQ9
8Il9AOqYdt/nPgdrVNnaaG9mIb33TOdqCHXjvM/v3LZiWaCggIAobj17f9orYlC/
nQcOXcpILg5UUfOSuwBRCzC3xlHwfQ6yvbFUVwIC0hIWNaZSyD8wc0oy08zPRDue
qu+UKthiJdEW1XsQpsFYgur8R/ksI20XFR+ATX19DMAzKK3ZgPEn4dHW+B9A4FDu
C2WSQMUKWSvXGFzgAARAyaod0g3psqFFzfdLBKZALaTQpWFC3wNCJ2drLKWUSPD/
LTsToEjUo07FXL3Kn4ZoRb/W/5cIQANOVOFCocaMe6r7P3ype5OnMpwwSfM7HlXI
i8oVXLDwzdxlNfuCYvuxSwlROVgeUDnVb4u6UAKKBvKAuh3aeUpu+26SmuSHfGb9
qOUeoS4DFqzrPpEt3aAVRoY6Ftjbu50w7qnUNSBhqlDggHkxCW7NlTL0wLldDhVd
egZpc26O1tjafexBxNqLSAS0vgU5pM2m0dM4AeitNXpObJumF53GkfIBU4csoK0u
Oi9invaojdc/L4nD6yGSEoQmnB5gTD93+DamixiY4liaTNGAVmvzy1v9uC8xG2+B
NV2K+fslbuOhAfy6WoH4zvgLv020LC+DkIMAB5l585hotwtuRY9RD63ErozNkDf/
+YNw2fHIEGW0gS4CdL7ksWkCUqyrBhN4I9fwruILwK3uGor18DRqj9SECxasFvNP
UGty3WLw2Ro3FmkH0rVb9lZoQYYfQwG4gjuRwSwYEMCC1IlNETUj4MzKN4b211iY
c7jHIQB+3w8sXJa3CLPbvrYQJfeqVmSX7LH2W2/dXq2JgZLDQv3i0+XRlda0awcC
5vOqvtQyd14A6ir19SNIj9YERYTuT1LUtBKfTmdmYiDAuDRiZDrKjalxs4UHjRvs
c6Lhi9bF1hiGygn8FdV/0oRZEag/U5pvVKY232zHhm5Jg6XLQo+9mk3ewrpuIK6u
sn6+jU+Gxi7PBQFgaZnYinrQzq8FUxqwno/Z/DzP8uXpOzdNptx3KLVsN5BJkps7
ml/640yjd8f/d9/vQNbnxQmBkvVw+ToowmGd92i7MdmjgxjVqANC9s3YOrGFbusf
A3fXNKVWkd4CZbR0n6BXp9dMEWORO1E+A2KJ8283UncNXHuhESbhXp3RPlzix2bn
IYGFxw+PKhyw/hZDZ5N95Dc4zA6jAHmHcTKPLj/HKlSBWbyPndtNqjcBGlQTQsWs
lnnnnkIfoymPKHrEy4iW4jqcb/hioo0hc/mDRMZhIxmaw6+pnYKeSRG+csJAPiTe
BZVbpCb93s1STkIQTkU9k2e1O941epeH1Adzsqr/OZLyA8S2hpUX5wB+KvTNc0bk
Dc2C5E/gdw55t+HL9zG03rdr/urfMNDjmU8POO9ME/LQVGJGWv8/vOnqdcfED1bF
EC2Q97YaJeV56L9VmU37EYf7JWZwTTAvTSBgItlcxxVJNSB+mfB4oDp8m2UkHPkm
bftNHbHLRaqeccSNJSv1ImtjVcqMANywPlRaZs76ByGGvgKZ1kAdFSJgWc1sDe8L
MKMhw0ebsBSZt41fPX0+KX1TGTBuwFUv2Z9tw2t9pr4ImvMOYIS0Jmy6vTk3cagA
RdPv1yeSvVYyvIniU9S+3uX/Sib8QvmoLjH0wcC7GYpnVichjv1gFT4Kpj5WXUOv
I+mEBMfFl7FZKK1gM+ebjeUR0NuD/J099svcrOpxQQv9Geq7hV6sCxRKIDZ8OiIL
TZMR8BN1xBtzHC2C1JxHkNQmjOUOrQalWfhwyZphLhlJvyjyVGaENq3hROtn8s9K
p038OzczNcuMGO6SGRgWITe7R5hN9GeZSlCGsitTtPMmsHcgRtqbb9qP/HII0AYw
FrXnJsWqIDg/vUknmZWP2Inecsi0yH8Vn32L7GhADQz7tUVqQVUAT74ImziuMJeD
Pm0ufsdyzxR2sOossU8gi1K7iAwwwKF7OVyxUN3JG/y4/2Meg6jbC6GmRiwwInlB
xtrga5HVJ4x+GUAhuUnBsgVQLDGoKcEkgkriijyr3Tlooz5rrP7O+LMcXXdPrfN5
t+XulvOwnmct/q090caMmb9FVNxjOasOZV2l5ipzhZ1j/CPvCL7p1B2OrZljSva+
yVGtPF2m0Bn+0ctl2RUE+ZdD7/qLVlBmfHU3QJKkfLkTuaDl70a6Vkoh7Tq2hllm
IQl/1kQbGnKzud14wxuk6eELa3zd8TcBIsa1HrJpMTJdUhsKfGVDRnvb/IyfMonB
ndYSy0MQcaJ554Mu/sp90eiAMCjElpvzrAighXhR+IMKPK6CSs/MfywDaoWz947M
S9aUejeKcd+xic+DZkVvj950ocQOn2yx4PykXsVrXT6Mc+htw7aWNwddBCKdffwF
03trpPMLqEPz5bk11d0yQY4nZ3dMXCr/JQibzpUIgHA+wClU3EwEhFS3DWmLZ5Ag
fPGi0iSEAdiCtzUUzrmLHywY/ifhF4qQUyBuvFz1rLtR0Eagxjngi1b4itaZ1OPh
4Cj0/FtrN2F9kSliXV1VxH8sQySHOZJjzH+mTZscvfCrhLJCtnV+BuFjz66NU8Yi
cefe6Ghq1jic5C9iJduM9PK1mVca2nofMKmrJNMBKWAlzd8ZxKsufTVkg1C6vMDa
uWyuLFYn6snYzLIegpeLVDfo8ObE3N+0Ulhq9AazktTt29G5ejO9JITYwlM/z6zB
KWMkWHmtoIftCMxGHnMzK1TUTK3c8HlJSEnyVgvMNgyTnMhTFw6aaDgToqwxu9EJ
ZtQ3GQoYMPCEr8QrGJocORIhsFlNsFjZNzgnlEb3H5cdlnk/zPJjoeyToD8XjntI
yY1hjmpLAanxxvxuL4Uk6t4QFKmMPugRNND9QGBW5QLLJLmcBWUVX1g6J+t9kyde
chBn5LYuBtPY+zQz3QEhN3d/1MN2VRccdHzeLEKvpjLYA7nu0xEklDWUqFA5QoGW
pBj1P1rkCe8DTVw1QtaVzsMGmKII+soVI0yQzT+MDfHdKgz2q9+v9io79Q6vomVy
ATqfv/S2yCH1/ztTYeoS9g7AF9bVCmqdkYWn+z9f5geG3HSStc4ONTuDgLjQFLr1
BQT0/lPnQzrAtk9N0vypNEXIT7bMR1N0aUTWzkxJjjEobnAPH/9jl8CPtFNh0o7g
uLhZKWmq4TJLaUu0koE6/06c7mym+HCpRRCQAkyQ2PkN514mX7QfEUpkzhb4YzJ9
pS50gNObZfHQ53ydp7U1x3V8/I+C+PkR79qSPeXDDNOfTsRBS6HknLNziw/2sDam
t1yLdZrPM0eUXSa9SaiZSWb9YvmDVh2CTGvy4nWz1gyPmRxmnK2O9F6LUWuQ95Jq
ucFWvn2yRI/eiGgPnI9WPtKYXmiNI9gIRQvsgaDxo9G4iN3gket5+UtCcPXI5UUv
LjYj77+4P5ZAfQlaZ8Y4aczIHqh/USeHud2/BD5kd6MRGWLN7IynCWgTs7MO9fV5
Q6k8oLd6kVMdeflAN00IG6Kep5r1p7ExQ/ZsFOw24e1C6ZhH/CwnnTRJKJJvNk4D
RJw/flM+G9XFD+jLEd98t+Np3KBpWHu1T1C+tkNoWaWcU1x84Uqo1wUkCj/Mq+p7
DXSbEdf4mvTpcPbYhSM2qnTei1A49U+Pqh/Ft9eEuFmXJUpgUzq7tKdC8Ci+z5Pv
Lsn9+Fok1mMBo3kwVMveJNBZilMMYIRv1SQ/0KGc44Shn4TZIM5MhZctcU/b6/Vb
Si2lmA2o6Yr2L29fRpFsT4B/MBbqAh0E9U+Lw2GZFG7Kqoip3OIWEULeizcx+XGj
fp3e/zPATzIsjvBlnbSz2+FHF/lOwvgWDg/TjGakPu9VwcDE4MUGY1vj5JrYV27u
f9cXaC5aUlHW376e+RGXiYDTGrsIlivExCLl0hd3i8NbDEYgsEFakwSEM1VKdG1O
rqfkUSB/eJPG3R1teTUZDKkT09fKC10sQpXhQrRxT5VaY/3DcoXJsUWKdN6JjMr/
B6YaDPz/KtszbXVFfEafSxlEb61A+ZYAsltX289PYhagwVJLJQb0fWtOdO+K6wQn
nk+M0FFXWE2PLbL0yzjqA1TtVH6UWSZCasJbOoUNjkXgQxZ9e9GnFQgW02Jx6lIw
H/5tZNxsmNT6z+SytLXr07b/jNn8EzjVjuhwQJ3UZj6wByZ9v59c+RcQyOFvoizn
hhiXeodFTllfIC83S5EqBjWl6VlKrEY8RKLyUytp0Zvq3jJQ/3kCokG7Fd+P+u8U
hBVPXHKjiHxQ9L9wjTlG5gsMZzH+REpirY6c/1k88vToecJS8QK7U6dqcOL1V3JN
2kBbBol+hzrBKK1zVIZatsUlTcc1Q6CuR125udqjYi9GpD5BVDpcr9XR8LPvF4dH
N+Gig+z+FpSTle1odCPCW+GtM2yc2AqPOb037Mm7MoS/9DYfWf4bfQ7CL0BkiU4Y
kPbyO7mhvaREKgBZnMVuVNf8caL3/UqkV8n53eUszd/UpnSUPO3rIJ2yEsfIkOls
Bx4vStJ/THTewpyMEVf1FOsDdlIXwFrqhNDHPEGjtFFZckhPmujR/Ntf99rnsqwE
5C3nMarOk5y630ngEHtjdkfv/+iVmKwK9gdDreHE0EERDmD6UIfbY7Do/oghHBit
WCd/JLSKDmLbInmSQQcd3l9Pyngs98NZ+LvoRy/pgZyGaqnL5Wt+NUj9SMWHbSqe
OoayfAaXRdM1irayh5zfEeFO43JG5mCl63Q0hqYWrYVBhD/t9oEbUJIwdhy2aEHp
DsIoRuKiusrp9wvrVdHXvjp1hhxncmZl8W6GqQDdpC1noLc8RChXnMEiJKXAzAy0
clmr0vp58FwuxNntlwnDYzBZQJBwEVfKpaWyVUlCJD5ikGIOtg0wx4kcxE7dV9lm
XI2FYaAD/dKombXOoL1runWnH/RiE1qhr8UfGfm4I0yFgwLFkp38apZtOmeyCJFc
KC4WqMN3eYc5uZ5BJVBTwiX3eIZ+TRAeTwnwcGeMhFxqpfaHOeT/fxAwR2nctt/a
o1O+H55sUKPkTJMrf4dkVsaW5TSsnD/v1bwc/rH2PS3XKEpaG/8dS0sbmWAFNWvw
lqxN4NAEswsH5M4aXW7usrFU9SOx0GWHhZdKndFo39MAlVQBb8bQHnoPlz7Z3AUj
NscdKGufmpBU9M6bJ1eJLYJ+UHd0gwOO1WAavmgYQlemK/EGmZN8axRYC51SlrCr
VOSN13FBoGYu7Gz5arB2xLHaecHHP/Xm0ysUDndihHU/ReEJrqxx+OJ5kQd7Iku2
vhcZ2Vb66EWAFLc0LC9kEMv4El9eQSOGl7f5ZU5IJrZqJYAu9b0zrsxHhBKACpvF
JbsWP+rFEZ5gbvFlekrDHP1x5yezyed43LrbJUecGiylcPZIAvBK7SemrH12WUbV
OKyeEXjyQ0b55ur7T0H35F215cJR9Xz5Kuyg5faajRI4te2RG3SwkDexnnKUA9Pj
buXYJh6+2muf0SA+XslGUqbmtnr+yEO103kGnWI+qTyx4W3eSqgcPbTPWfv/4APV
Z5gC9/nT3A929f8FbAHwnn7gN1tPQfTaUkzt+0evS1XLPS6tWHBE1cXE5DtyJfx8
BG5XhfomgTd8nkrXimE+4nSuGHsIZKF7zYcbtOwrFn/0Tb2zv6J9R8gVw2doGSyp
J9rDFtCi5IQmXHegv0ngju6igldGS/NdVQTF4rbL8thkRYJEG8WjUVpi9fSX1BN9
mpM4A5sg6r4+HRu/WKxkvN+mKwrcT0wheA13e8Cqbzo6a7yXvtk19b798W6yKo+w
BFXcUkIgRt0tym6p8di7vvBDbf+VmeeujmwOAgsnaQ7kRqR5p+sqCWnzmHCybraB
ATZPIeaST9rxns6M14Ben12HyIqxs+j9IqVpys2KF9VVLR3xMVaz/5JrQ5aai0v0
t0T/f68x9n2WxfuVnSsnYO40N82i3MdZpNXQ48b5ZGVl5221FkVZCIQeiLYS7jLe
vrJa5/gfEpDZhMnF4QADNVpXPH/5qfeVKQgqHs4ZE42QztA68/hx1HfP4vax8zpi
a2NR3JBkRHd+7q6WOXFS+S9+ysl1SKCT/MEYKz3IxhX1oVyeYMF3vPkCODVC2zV3
l3gjWC7ZN/Gn0VeVwm+EjHhllkob3OOuskma4w+merk8vZ2ac5ECS4P5G5dr2bPW
B9l5y+ZYhlarRDLcywTgvMfgGyRFMSP2puO8zLdm5oTI03k+42v5VOwUW7/6GGjA
FAMqyXtMSQSf56BPMr31/GFcQg9NjEyNqMmKSPhCbAzfUb6qTYAPQSd0axMPFLXz
yhuQQB/RM+h2AgJyOvbzne1xETBpj+8I0PH2U/3wmipE6upyPSkh6VUbP2rwJ0Y7
aoheKyX/C+mVhxrgNFRJRrLePfNaygLRAfOfhDvHQ230Uw+N7T943A9/G3uUKhJk
5TNywVhM33Y5JKhY4YSsmvOPfImTemXVaI6INJubsFBzIXVMuK4qzp4kd6jUJFim
S6/Owb42RHdQoiReYM3LSzW7Ng4SIJgxpVyevVH4f+yek0yOatcqrGx+4P3nVh3R
RTvB8QOTfl5kUqFUcx9GYiG16lRLZG+VO8O2FrXGgQRu/g3zm6ZDXEgzy02DgmJ1
CsgbmMElSOJiX9aPubQbcapn/G+3F23daSo7jA4GitAQlWTqxqO5GYygH8bXuv5i
nGsO9Yrm3dfFgzKGkGAlEIYPi0TzOrZBjEtnCbou9MowJfSs2rC2n3FNji4W8tKt
FJcApK2asKp0/oq6WooODV2b0Z+3krzkQIONuBj3wdNGtTYK2xwd+Hwxro3jOFAg
4rFV8AYocRsF8GzYPDgUSr1lci9thN3sR8OrxaPhyZIVKRnPCTgHoUO4XpTj3Zp3
dgMEwt+dQ45TKopdZDqhzoJASI0t43wYIDt/yM6UfihHFC/m9yPbp9g6uAkrfdpf
WloRduaGjhq3O13rt+CgzKNdJbAEOhqpFysXUbzxDSu6kUTh6WTJaPoXje+ZGrAy
5ioFQUpdbYU9P6aW+CAlRDzh8hcxfZeIGQe3syLkXUPHppdbOubYxgml3KNBr4bC
rep3Jz6AQqbDr9YjyWVLNZMzyJKgSYQcBcMFPBIov4baDZUftDPzy3PortzeWYqh
meGjAiWjwj6HRSWtj/MptTLMZTiIpbADCj2CHHMSI8a68FO1yLXIMWfRAu+5MZIS
a70GpzF6HnOlZIFIiEjAva9fC0ZqTKEykYA3vGZJnWVkQG6VIbZjCAuAqbTkc1B4
dPPZJZPpWT5pkFXUtJgKnNheUCKEpLlUgj6tted3/ndadcDyDl/my5GcKKoXiUPp
4j9bow/aDo8C9/07oZ9HAKA30qAyHVSExaqG4ABB+5/5y6BkUrsUyp7q46fUl43Z
X5NujoozgTtXyzZ0W13pl+SUgKaIlbz0OU2sZfjHVQ8+eumM5mAuhevAYgqPxMH8
Wb9Vs584SZQbX1DM4qcm1iafngaPpYD5mZECZN9Ff+WC/dzorO+5oxbUsUT8ukDG
7zQBIBtjqWMyjRrktKddtEW/X2hj1Ln9S7Q1HZURkD/P1A8j9bgAuft5kGJq3j6X
357rR2lB2GWPs1Gno01MX9J4522/01YKNWVMm6BtNwKlACvnXX/cHCbdsutED/qf
nOt/nHiykFsURpidOu+M9hpOxvMItJsbuWD1iDjhtFqQGiud0/qQKX/STfmF0RWS
BxEQFA2d7CrSbEa7LcK++6vy3sKLBwcQQlqdBOoqBR4Ggu2vcCizJb+8p8jxmtXY
8iwXf4Ki8J4RM1Zr373s6efsSqgr8eCzBWIZ9KJ9UgWZZ7Kh1SAG8v86GQyEzdst
jtEtXBDLFt9JpQp6QBA0IAZkCYbM7Fcquk8RJweA+DQcD514y0hMHm/tH/iyYDBY
t0JFfTkgalXobVxtLwDaddgGhwoK7tTcrBf8ADMTMbbFryaukqxrb1i6jtlWQAdV
HB4wRlAAOH315ZS4P9uGwEiFqLpW1qaDN7L65YwIrHp09WqN1XIzwDT3E6ChCGTM
r1QDcyh1h6YeM8dYTSKTGtbkNnKXdwxsIVz+hap+ZOVZUQY28eyQVrm6dYBjhYvQ
8kEmkbgtqs3RSFnN62FsmgnKsm5b7GdnaV93q0uoxEexqIOQJi5p/yQnc5E0zKCx
pO0BJk/Y5mRhihNp4dOZl6WUMWHOKu7n0vQdWd4Kur8ccNxI0VJWRRCXZmm5h2qg
ZvAHDBakvlMhRgt0IDeSQSGMrXjkwcBdreX6GX8P2Dl9P9btj3RfJBlhKigt1B5E
6Z9tOZ7+j89xX+x+dU9GMKbksba9ocURT/nxSwOq2hciJjEF5lrfWHVJqawGlhFk
taA2G2+4EWANuxvHdCOvDtoaLvyxPgF/oZGCfWMCdXaq3yirUHMm2Y3QrTqLCEzq
+YBk+jxLvQuGuXh9AEg+FDQqXCL8A7/xGbzOfSZ68aMuEChCoYmX7pppRZKM+dD0
HOHItCt+ULPogX4fukYxw79rzjJjlG7nmL0vYTzXfB/9YhjXpUAPUUnhu1ueU63/
e6iecRJE/4b4JHqhdM3+Rl15sXlB3XTyLXJq5gJHckrkffSypbsA1vAWMQAlB4zE
Np8JlHi5/kmD9PFb89dLKAvBiwfNRWVlAWn5Sml9Blev/OoUv/OTa6OSZ4h9o1TA
eXzdaOKXIAPXRA17QUNXLm4YF2iHHMobiZfG+4wuv3zsAqh4wZr6uLIbdFWKFVjF
D+OrNZb7KIdgB6Qth4SEwoZKc/Uq8+7CMvUR5RI7WRmcdDg5fSslGJfDJAxhRedA
P2hw0sk5dMO8ixCXsVPdQlsxAjKB+RxLjnYQgOKyiYsNkPw5fi+a88UphliRm5U5
1pa7tQH/sG+U0WI+sgXyn8sRDrLROdpxCXbfCowu9SfuUlMuww8vvjrVDqm9w1XN
yr/nT4ZsZrSaLpQ95f8lcPAxnCg2g7Z/0FBW9/YLicfv5qSiS/IbzteBMWE/xRcP
DDkcSZ1GDrOZB4TtEiOQn54wRzfOjtfUWl/6g1a1cO1+kkGSMG2EP+QVU52RCslp
Vq9SszvAgK8rEiZncxLg1tTEuwifVa94TISacxCLEQybKfM0eyelGHllYG4p9Z1x
7G/8hIoxjSmqMXUPzVLKqXrQ93iGmSw34GyA9SpACOi1k9xagEBAZIbCiAFz6N7R
YWXWb39SerWOYMsNgaJALGuQHLNTYtsLkNt8eKAzVF6kZolNl6oO9M4SMhBfD9nm
JFa8/cI/Dhg5XqkQZ9gSKdd9ORWV1khOQy6XuzLt89gLNfpCiA7ArEkvl7pheo/f
T5a9NfIuNECLvxthbt6MlpwQfJAt6HAJ3B3a46UhoxgLKn6C2MabHUklzzaz15ME
cLD5SjJUMOgkHnE1+CR4jglSu5WaTURamyXpQooVSWNV38ApJBPZ1Irnbbi6bt8M
1TqWomw23K1lBbSXmve+rho5mygkrH6oJjQXjuwF3n+Ik8R6Jt7+TTfNAGfQlBqz
AHGHMdb5YvAEyAUxeGLjM1RvxPRBgQ3L4ChcI+FhJCSm7dSR0GB3FYwjsVNSL0f9
pXpzW/sYA8lusnuMyGDni4cx7ZrqK+m3MiJFxI0m5NfIgfZ3iWTayoWuGQpS9G5K
87exQuevMHoO8OCjMLxFET8oYjVb34mnRI+IrytuHkz+OphqntUjUlDNZL9YGAuP
C5506t2Xx2SY3To7zjpJ5MRU3MD9F90qpmbLsxf+bd/MTeVZCJubmvfiYv/nDE/n
zV1hbZRvfAhnyybTXleFBsPjpc8MdgCRtbBlzpLJRdgIBgF/AKF4+v9NZ7F374CU
TyGFEt37+NXadygh88QwyNsiWYoFNbmU2miVvh9LuJk9LzqdQ6tKlt6nhWvT50wm
4Ed+zwQNKmeFLcUx1HYo3UeAoGzadLQxeERA6kYOvd9nG6wY97elYy6ggmrJvwNv
a7b1/YNTp/JMXEOymgnu28EQHuVen9WpTUCdw3XVJawK2A2Jhret+M4R6iSmW/uA
Gozfb69Vgj3ucfywasEguHZ8LT/RLYEuQh6hZkuEk4MghmhmtSeXPFyOr/4SWAVV
xQt1ljRd1KoS4CeNE533dHdpXIeLFY25pw00JCJ0AK8yVEaeN+G+k4VkoMvpApoM
zd6iyKiSRZ9S6fNPQjaz5pa5/a+t6gcA2vxMNKDbnx1qfdcAdXYUbdf633dQyh8f
f4CfSAEgllGFyeBAiZvASsEanC5BpVgRBdr/3L0JSPUVw0uVX4/uF/5D30N2jAKX
QhHTy1rOPkrVl/iwYMUHIC0owce0WaksU8CWRIYr2QSgAo+PCIvg/L85v77Kh+Oq
4RAT7eGMoQdttxP/m3jVnzp4lYvgiqmlJkK5hIz3yI06gAOEFX7zKXIo+/l4SOoL
4tVnsQBWzKIAV4ul/xGlgL56CYt6eZOt8+WVp60YEiVUmtTdZeF+zbOWNo8UQ2pI
CjhZKfr7YtxtOKbNQySwt0YtqfMBqrIywFV2LpBhL0n2y81FHDVdr7Q6n5KUBpZ4
KVacn5scJnwTduEMmJmx0p5QcJlvjHDwfZGGKMGUF7AUHcjqafapfY30jAYHU+0/
nrnlgbCcUQ8y3uV5j+UpgpzMoh59Ui7KRTcZK10d+yMGnrxHsnm6LA688Uh21V6d
1XDLHR8s6z2jiWiE7VQGF/sj/LYIExriy6urrDN/oqk41W9EtXnyHm6aRUdv4o4n
MGCBCKAFh+TJYh1h2O2Zv0VpqSsjVjnDMvcalIOpehIce7YcIV8EjSWSFEKeuzMO
XghzyHXeGGtxKR3x+VX5hsRvwD9H1ZgX+HmnXlFH+wR8vS0E10m5wrf72IPgrDCr
ItT0/FOK9C2UtQYbUEYAy9TDJxz6R4qaj7MGUeDOjJkjMj7cjAo5w3dD6qhE8GgM
5owHhaiI5StZxmI7RuyKYjVUBawhUSzJKSmVI1V8O61IdrRrd1h3tCmSooM4bSwT
6G46oFU3PiUu07AMPODJhNVavqATfmTLK2hkQYzcSqF9VTlGbaQ9mEl2p/OilpTQ
IJupXUecIqZwVCYhgkoBeOkqKM7LC0R86DhCQ6v8+ZZF8Iqj136jKrLSobQcmBxR
Se3PDHJmbKNcCM8GEeeEVC/V7YXSomRALNvs8M+NmvfFVRVsaHxI98sLjb41c9cc
koY+75a9S8pDPkUGespWVsB/xB/F4Oq44gwpd7il9zMw6laZVxhhjY+jI3RxTRUo
JlJP2oSRvoBz6lSosHVC8FQv6W9fuAZF52/04+rDuJmdQ+o55DOxb5x2Lz2mcxS3
fxZ7WN9dXJh6l9yuQrO3m+5aIcXvPbShAv6W+8V5XNRlLHMIaQ2vizaftpmaRpl+
pr9GsCtqsgzpPXrGXHze9zZgvIHXkiU65P9kXYfIquXhJARjZJLIiiRcrDeu28Cm
WTw6MRj0kLQsPYcBET6aHa2uF2X/u0tdMddn/yIrct3udoHqGObdGZhvUwBbpJ3i
3cel0yRMtYxNy4plcjblP422Rr7GjVjF5nXxIRuxcAk6JZLehjX2hIBR/Y9yzd/O
KIjVqVU5NDC76P1U4fNkjzTjkMpODE3WGTEi8tPbkq3OP/gOfnJL41nKaTSGLanl
6EZu+/wCa2262R4E9NAcqbReFuM7iX/RvUfAiDBbSkm7xKs5VR8s+Ekp46dt9t0G
SxwfOCI/G61kIbN4bNmW1p2q5AaDGgxSjVd79NCHKW5bJHMmNXa6tP3I/EhzZdLx
7zELRtwkBebhhdNtvZY0/Q11uJn0Injg62pVPUGYgh3+NjoBHSJE1NH9LM5g5L1c
VtWRh3q/YvaqP3JJfaX7/fDDn0Qza1bYjcThDk8OjWvB/gYDM/Km/N2IinttX/K8
MrtI09ovgU+jEseumG1rwoeZ5YUr5uFRqxFne/p6qGasXQFio/2mOXgPr/KfbmKv
+wctfTWDsgoqhk5lZOr4lYj+KfQ6kt4qwB+wUpfqejaosP8vFZnsUPvmOXuStmca
687rNzsN8SBjzfCDlH5/P2QtecxCh4Tp8IH8ncNnF0VuM6yKt9LRFQ/Jpy0u1FgE
cfGVXzuZjErndoVKRN7vM+Xo0hztmpRNqSNx39VNmlGxO5QCOlt/HOh+BuJaHF6I
3a/JcDl1H6yT+whzEx43TOTFaMtZErqIwHQ2YtmgBLEBs6QtVG8WZ6CwFGaOKzGg
TOLcvvt4T5xfXnGQRD90iSvzf4SGJdcW2ORO1nIZehVgtTTpV1GdSxl7DeWYD7/+
Q5iDq3NVQISeqMpSw60HjFuSVa0nbov8syeOGKBDCUu1uQvEYxzExlqbahirmrlz
7oJjezTj+iNuK8K0CNzsXattAds6wDZlZpqo5CGKnRTs9KjlMJGP2lE1BxPyHiI8
VXlUgvDaES6P+SosjDtldBwzOB0XcJWCSsOxE9Hko0rnzJbOUHd9dQhbrxNs/SXE
bYzfCZ6HinfJZ0NbPeZcpLW9wKZM8yGveI2yCNxk7YZA69MvGlXyjiez9oN2WyBQ
vBOB0iLS26UyWKSc6KNZ0jODGYH+nomalXqMjNTtzmBCgmRzOgoUZxwQrtbcVWkd
fTJbnUBVglx1PbAVsmK7NR1jhfAc0uFfA5y4p0G571ODqdQEtqWYJaJhIpXoEhJk
Q4Gpb4Nt1KcjQWmLtunCdNmgmO2YKMEZAFu/oeVSMFmthr2U5TfruvJKE0Sc5vZ4
G9KGBoQMcbpstxKcCKY6t8Nd7jmhHEhrZDYj8W96/1DykDkj1kk1iv8n6IgBxyGj
eUklFCv4OAKBMfz/yVRGYRWy/CmQE7okxOdz3dfLrdnEfeUYLO36Xmq2Tmkau7qY
/l9SGpi/bMgMqC4hWBteyFe03bZdnf/oEnMSn2YpWnejtf8YOm0+xYT4/LFDOfb4
K54PwkLn197lQUsl12k1d4WpzFPACN2R/ufkwWz9ZbQh19h1R9AL1ehRRjksucrT
84w/Xp/r01j0+w9gEsP4lW7xCvKMMjzS5SCt8sTVybTa5aKOMYCSSKOsu0o3Vcj7
qBBryuBC2TQfD02rW83vu0uPl4Q6tHzqU69UfQwAwjrXGjnPEPRxnlNYAbsS+bhA
zWb3Y7eldlzCgzXHEYsCWXbqvegv7/DXsBmCi2PD5WEsNOIJADRJ0v8d3ng7bxCH
SMBNZsu5IIGaEN8mQG2sh8N6ovNtSA0dW78I1IQDHTn4cHwbsHSvD7hTb+2MnDjX
4RTC89Z3RPrnQMJNpmsg+AZDnmkT36GJnGuMBAgkjqXEX2eSds9HdliixfiKAD1G
b0rynv5OgvU+psTLC/5Ls7GJXUQwLrXTIQMULR+Pq8gLmtWbyPphHScHzVcXxs0b
itefJq7o/JPkOJs6hlhldwDNIjJMNOlMPlaSRQNky6rJu11n+uL5c1oAx+DeaAYr
d7ve59IcILB1mbtMDs+ZjjdCCs3x02U82QGQbc7Ft6LC8+4UqLivWeYOLVtwurys
D6DUnr42OKLF/L7W9z+kqQ6x2HbO30AnpXRIAe1tnMcVo3c/bmyULV+OBU5JNYlu
reL6LCMDNDwMlTBO4K490qBJW4Yf7iJ4lLeFzOAOwGC4x5B8DUIJ7WLeuQV0ezMq
OC5E0yOB8/H7w0vvNYXjzzT1KMJAq/bOZzLSTckzdndcE7SRJWZay2V0hL635OXw
f2QtX+j7mtH1uBv3WjU1ga3BAu3gimW9Z/e1g5z8OvINgFQMb081eAyubhmoZYBG
EUKDgFX3x71rqwMwtP/ImazWr180Rgp3PdlZBEv9J1lkCRbqMbWLJGP/HnmIBdzI
BwZtRqrlgqfRrt4WPzmxmwd7QIGn6cixbylcfJBm92sw+et5DcuR8RZgO4RfK82R
iQGoUpUIAef9u1z5k9hTapT5vwHynxhVhNl7oq5iTQMsVQwjW7RcmldH+4rnxiVh
yMAyzDWXZteBYjok+G3HQ4h3vULfJsSIq83FnfuIaAoQeFQrkBlFvim/jQdEea51
WO2918TlsGX2MIW6IJajM6wUIZSm6YHNZM24omrfDqaiYdczyE53u9hmYMPnjWa+
+Lv+fVmjs14gwZ2ysW1tJRpTYoogeaD/FxDIN3enhJy+QwTd9ipVeLhbGgLbqDUM
mFwp7wig+Redwhz2hH+CxBgNCVFaIOB1tHGITx7322d4csMbEI8r8gTE3PfGF9BL
ed5n8aGA9d4KnlcAmXyEGTzH5u1jPHyCfI9pQf7qPi2kzfGEPGIaIV5Ob2AMw6ak
CdbrmrVhCaJc9FfpjZeS2uMXXtL6J4CUgUklKPSH1r8CNWR8Jv1Sjf7zndHsC9if
CBFSf9rkrdKAMvs8FT581UDlyKhwuXs5aF0qR4inZ253pD22qcUwWPJiKxBR5By6
YTFpNvl4JJmefY3+5MyEav8JZh5CraPWyCjddS166BfZTOLfS3TH1gPbtHr7bnD+
e0RIjVu9tCB/FyMucJ5sIFWvLf/danhZ9Y2r8vo4YW7NphyZHrscG2u/v+pwmCh4
R6bJvS6l++1hDihbAKbEUBnFfF3HvzI3/4SgbS/EodqauusIi+NPB0Oi02axxyyk
CgeurNhSmE4qpZrclfWeNjuCZpTOIRQhMgWNq4BJVsTsi7c48oqaDxbzKCIzGFRR
5ovtd2ye7Y/suJKukZhmsVoLhmyngkg8rp08hke9vrGlxXoiUtmpXzYIO5x3hh+7
vy4VFGGcRBaD3i6tVAW8dj/AuzhOpvlx551pMFL8TVUt5qfzB1L1Qhe+NHC1RVPL
iPnVcMd3s3QrxtaJV6kFs0Z5+RuO83r9N+Vp1Sb7F8P4MRbiMHg0wQINNWLDlLoT
/EeU516nN8rR23aDLuxE4g3L1UJbhgSd53npFI48GDcqZbYyxbOlIdwwTcZEj13L
FbGbe1bVEWIQxUSlbmTWPLLP20+bGBo/jMt4kRSZGSyL+Yy5h9CO+ApTsHPdmzMG
ByJf87VEiKuvQKxKzDwxdcIa53+3HOvt+u9pVbKKn3aFDOW3Uub9ZHP4BbgUcx6e
VoJiux8jd2TFI0aHhGQ/kvahN2kZDCnhwYbaHeSms2idF3Q9vUOXUoLWcw8MGpmA
ZMchD4EDA62CFIgU8HyGhGn9N3M0bvaGlm5FuGa7zduYMKHu9E63/okHesC6jgNM
b6/H3hf+FIRXGLLgdthcUnqK79cta7RFFnLRoo0zxFQPYGrdAW2a6DPRSHV/1Ngo
wAfdBRFX8sVZ/s4AFk1EHTNgQB+nJTzMCLeGSZKbUrUrCdUm4agEMUN4aqDC2Nqg
FYToXEQxMcuLN+pTd83v7mUj9ujLZ1UT5dRmm7oxrKzJxn0zEqe4nqXlU9Ev2OAi
RGkGkvCxCTmU2l0GN2fypQz463jWrwHmZmhz4EtpjKwS6wAdJPDMIOk8/4k49zN/
FSlELoyQ1bZhKO24vBlKh3sDTIW51HqKFtH8wfMJVOC+BGyIcd1hNBds3RLNCnyB
bs9VJB4MKcrNIZS4MrLRqtw905F2UHiXYrL1vIsRzrqiQb6Iyi54SMjWlSd0DgVN
lSS7iuzdnLbRk5URbeUf0yNYCjAsHTi3yuj7Scj+aiHqSkCn2fQqu8cm88+E6G2L
40cYn3vhEJ8xaPC3+IxPuFMM5fk9+fpGWJdBYSdTSVnEy77V2LTPGNJPtXme0lT/
GXsdqJn5al2aDVmcpxDqn46GWDJ09aFcSJ/+ymWWrEzpkwplfX49tJD/+mJWeG85
/Z1jBh7ox4/klUCJ6h1jhAvUjjta81pSojU46XDKGzq/wrGh4QrC/OHGhCT0VjZO
eUx61NyGPuXf7lLf8et6rPwlHzI4o0fszsu8tWV+/afaHoYsl8VhUbsw0HZZvtsu
TS3yC3x8VQD+iD8eW25wPkPUHpK1evv7C7bATitHwvEpeR3PBag5dydfKn9X0u4y
AYarl8Pm45MwLSJDxVm0EfsUpJ6p2w9eev8gMPGM+wPtjvwPeFjjycwRN/t1KIqf
BHXDjQma5fF90or23UnBn+ACa6576oBE/XwHotWA0APs/Ik8SJ9NUxz3+CFil+9X
dCsmdYP8qgnzm0tbTP8VB3b8fmmaKLlRfkRgib9UAyMRt+GfIQzU68OQSELkLeGT
ajlZABoqdtxgn1OsrOeHxGMX+Lluy6nyJ/VczA5j2jwFnhXIhw1u+DCrBS8mzT89
uP6Zr160YV5MGyHmpIC5gEDrvNfjSTJNJlKQf6BQbzUAiiI8OgwvIgazLpB/Slie
j1XExQPR9cFtL0TPs37OXQjRfMJ8hH3VOOBOILEIf/8GGwiyvD+DLIwfxgixgkdK
LKOCttzbda2Q+x1wjcNtguhlGTi+zfCm3Bm7JHFtMGM1gXMgMCFTWX3WX0OklTMf
qyY+OFtNK++9umXqeF6OyISr3TJl2GTkXVkW3ZuLolibuG1vytwE4toCU8FOwBto
uW9xoT44vbfopp/FEx/J0mktLxbcNxk2abV3MhBotjmfFrGLTalK5IdUW6C4AhK3
WQzG90ZamhOYZJezz/b8vTVDwv+1JB1Bykc5NoQbQqo4+RkHoGjBj44UzXJiRmNH
LMdIszN6u5xn07NnVDn55uN/xj3P0l2eBbFVs4DSdKpRFBBNOQH7oyvwMKkPINNq
SShv/Zy5Ld4apxiYYfFuiIP/ZCWKrqCaVVEiX5mLt1AuCnDgfWiUmb9APnBsmbyF
21uUVRWqKgIC4/P0bzGmUa5YCmkkrppCX+gfoJIp3eq3S8izExvunfdvo/E3GaX0
k1d0gHj/HgzGRB6MXOM+GtiJXELyg923+WQBZOhKIolw6gvL36a4/Y/QNXa7oBFM
1XQfufONB/5MeRNRPKe58UBr3i6PRWs//Xyh/F2Xx4J+fklzbKfMfsZBj4+us9it
C849wYV7HFqPWV121NbSrDOxw948uPfpI2hxB+TNllfaPBLXUzYigGRv9PVNHCNu
2TgrfSVv+WDBRFV4J8rgIf5/HTrqVDWOlyKSmz+1mmKYb9oi3D8P+gdXa8kkwiiw
Sx8fqM7I8V3dYtQN3FcZ3BtJOaK2V/p2QikHAZQAcRRyEWH5pc4jrcBcGM7lPza3
3X0ZSL8lBA7f4SW0S3J/uTGvOHWS0W01J5bkjOX+UrJ8yl5xwWZmg5EHvwYm8NjP
PjRZHXKQhFM0vhw3wmJ4hIlJrDChEXYMdYIujL6dHmhU0TsFmN5QofrKOZS99a6p
QXyF8rcMITS8RR25EaRPB0kyMg1QFlP10crVy83jQk0GEnt1mQF7ZUo47LUXf8Co
rJrej+3+9nJP1RomPaRyHUKVVZ54OYE19nhH4TOgs3lZqhel7p63ju9Urc3VSGQm
Fdf004IcW0Gpci08sieaZExlESbTOt35kj1e/9zzTjnfgC0F4+NUlLkGVm4O0SGU
YPIxXVogKn5yp6QBqM/3Vfzr4gojams3X5pixMJDXHZZIUAk3l4ySuQraiwUTIhT
r8Jil/JeSZ2HzpMZhSWlroo3npnTfXhivUm07TGChgB3ZlBio6w2s7Vpj2taPksn
8x3v/LvqZWiCbkZeYJXGKg3m/6AkdX6jefnCj8dXEnQtfrg+gp+BIY6COMV5XcIG
jGdw4YddJXe+FK+vkgouCiXQr77JAKl36W6Ntm9oC1ETH05phorfqjQD6BbOIYLG
mCk5hR9xp7tNnTMxnfU+5AUExlAzw6GkD3gnsPO0fKkvXCJKpor3866gcFo2FDor
9Bk9sS9mlRvH9Nri/e+kG6tLzh/6/eFfcUNeA1NYKIRQYoD5V39wtC8ilQ2Lk4CD
75m/LT6Tq07dtLlvvZrhlU1sQlXOL2oSlGjWwrVGChFYkegzq02Kd0FGs5yrpre2
fXNYDDSsbL8bzwq/Wjp8fIKOOb46O9H7CCbdEvsba+LlWg0lZ+jC0DFjpYhHQ1Va
lBi2F5FRYL1FzO6evy46fWIgEVSv1vXX93jdPVFvLKpr57ZKIe+InUBoWgREFSgD
Lbz5NpgqLeoddtNl+YWl+nxLIzp3Af2vUdb5y460Qh5Q+A6i2SRB3eUUYPHiJxSP
c96Wd/3D4gsOltBEK41qs3/aEMqO4ecd07TXin5DKhiOimDIW+X//wBePAXLCDwJ
draawfCTCjsctQbC/wZmbEtbW/425m0amObnPUrgNl+WfI/1Tlk7sqtyhAO4iuxU
EJEg29f3SJS0vGjk7hsPhw8ZgvNIoq1O5DMIC0R6nKblQIFAfm8KRe3aXOBaJ44p
0Wi6su9WqA1f3qP0PuoCkfcF5Dv/8xPzLyP2VPwvSx2N8NcciRW8y6SFIfaY5soN
bZo/ufoTzpTckOhHQpf9XUDReO4COowo0aSXUGlYk1Ll7Q1p3SdKHaQ7mdLX4+m4
kFyzjwPGiv2cEAK+aVQ2y1XtfpEx4avOSVzQUq2X98tSTWfrcxN15tGfVnicFb2c
GlGmkm0YIucmoH4zUl+QN7akSToIbSPv6+kBBMRf+QGuso0Y/IUitFFseTUNB+7f
sG6/eOUDwvjTD7LA5xW3zR7RB0WFeE0WzgTmMpjNZI5KoM9erJn5pSc0R92UOfeI
f2DqtTCZlUCC1+P/GNIlLbWypGAs/6v5+o743zGKwwTDQaJtwPSFPlNBzRYKSqnJ
Jy1C8G8M4n2sx2q9evlLy6J9Ve8QD5Br2XDfjsU+R/Arz//K/uKawTM4NEzM0OZ2
JnQGbwtWPeHASSNd8Y+t8O4yVk03QxcApJJKulDRkjU7TdNL/jhSRz4BCkNee7Lo
c8Ghblzucqaa7T0giX3yceRnfSBiLHI3JaElC3NQLPCCu5r9zjqTfXCJ+XnTHHfU
zt4AlUN/vgMxCrMcuJS1i4MblzsnZMib6XZ2+rw8IITZIBqvGN2gqWaXhGEbmdCm
9R3PS2Pui2+i2ZYk+2LL0s0iLpEz3VzFYh+ax75W7NAJzK/heEYKVYbZ848BNsCR
j7uEq5LbCKklZ+LR6NZmlMQ4LH3rm+AiyAgyYqeHHiRd344KCP0cLQLRe/5Azxm2
yvEgpP41chxnX3mggo1FZLuZOLS1vBB8+3zU3YrLeviXTw59Z+EHvVpjUPrSYoyy
UqfBO3BeeL7OLUcvCWEUXDqFDVjoKvYp4ZLPvKxevhNxkC4tADhXiVqdOoxPB3J9
FdYmB8XZQnoDYvWDfomQlNXo2FLBXLc5iFQEpMOBZzkPj/PRfDfrJjRHlkPe5mLT
cWbCH4rqu4S0PZEVaig10k/aarDInPr97fI/SxkW23HxuD6ua5HQqoZP5Oa7/HvY
XxRfYSTqVYYfnpXt930cSOXepon9u6xUorVavC5r+hm0N48669/xuY+buHe+s/WM
Cu7a0oOEcqg75SGvSlmgUIHSrYSzu4/bs5gUTbX+UM1IVetbnF0hyY2AbKO6u0Z/
IDiMKAaeEpq/IJsvcFkyEhjycfWByq+rR549CxavWhUqVHqr7rDReuqxmRfvKVLv
pjQNWW8LEhL4gm4sA5/+jBek/1a0Kgmihivo9iWmmhJG97SfClga5VzcG5RozdLJ
OHWHbsXwK6M5/qc2OVujC7bLDrmoDVb1xFlEMxNHu7igLz+UnMnA9f91kbYmEemR
giAKoVt9LB13SuBRnW5iSZ4K4mw4uah2kOUyiWlGNzM3LbwTFruIOMF5Il+vhsVM
GWv/CqpKbyE+WM0efCmPQ0SvLvyIkLhX6kzuCkdQQs9KRsCyYLVqeyFjTj61eFVH
PzxOsYU4OhtglAIMKOORLhgH8tNrfHLw5JdUKh0WuxbbOlpFFba81kTFjxcnnSLN
0n6LIs9WmYAQmItb3Na8RNUDrvhOmDfNYXNeakxlNm30yBTtUVGhkmRj+wnKomJy
Ew8nw2n9kIITHvZC9gjqKVXGEOJWWBx8JcTu6fuYxez832tCxOuYevaAwhjUEVJ3
/39ZS4K+i9IEUrqliSWjDeN5zDlqaUale/zkDJe/v6EGmgr7wr88NPGIio1fIN3H
yCHeFdGxCK9gthe8sB9sBgpYKsgMWbO3NB2fLRNpM+ULaKjdlTXwvOQVpUJ+qMJh
0x6n3CXFmdq9CzFHPJXQR9+bTzAaYa8UHFHPzDkUaVtdjqGjO6JLZNrAJyVZClHf
cg027OrhoeqAsDZB2PiaNmHxjVUo4J4UqPwE+g3DiaVvopbFICQI+1HZ6tF+ZrIi
Q8fprtv+84kDpUyaW52CA/uLbFIEGI3f0f9Hg/Rv8/4tL/CjGk7okWBrXH7EFH9b
esuA7/AqlWGtw5W50p9kDI0yR+FtaGVmwNVsJmKHc1NAssbCgE9OX17sif8WGovO
k5un/MF3dFr1UTr+ecA8wm2X9JDzu8izadgCSGfqeSz24QuPqmHYW7QJFRp08yE2
wpGpEWPNXFb0kOXBefCnVMexT6kthyxoGmo55dKsa20ihVjN3hVNaIYwKLZ8XGvU
J8i5f/PgLkPOexWVHwkUN8vOr91COE4GsMaZUJXXbCSi+nbJDcFsv8G+Fw/uKM48
oYGt71mPtkus7rlmbTzFMU6iZJgMPwJYiDooAcNfiC8UazeHszmcEx1sxuCl5w7/
lUgKdhnvsxEN38SgUQr0uEPwgXU5yvxMfO3wXEYyKtRQBNbNu09ndfph/bAndwpA
hheUwEpnWBkvVRZjfIMzSMHarm1YDqxX61D+K396V0GsIE1y2fF7DmcSHl9ofKNq
5M2298IfKQi25z/laXYexMX7VLVJIetZ/9G6fZHZLUNYxpYi0hPF4Uc+CfPbrFWD
zoRyBDdHfKOezD9HPZBgOBDqysmwrMvjjjiIKbKJ/UxTPY92Mutig88eNb563bDj
ofUvAAWe0/At9jSwR18et9iz7d5njIWKV1Lo023lJ6BEwo2GqMrG9BI5MjmuqadQ
zpTyctW9+OOiO6vIFg/KGZbEJWjpPR+j/1iBpEMJy6Gjn3c6YrQ6tbwzSSpQdtez
tPgpzML5iFJaeDhTktlD3n5iaRWkKbY54Dj6dFqAMysCEOYM5tl13M5TiSrCkU6J
2ljH7VHDud8VTocXQzdKn+9bZj72gerAuGRrS8cGUVdEdG50yhm4sM+YOckBrUvf
DZvO8l+fLN4338IKj7laUPSnWUiCTsGfXQxCiEGP4fNCv/MRWiX5Ite3dCAdE5Xs
KjzJOQLFWyIby6c5C7SUzGA5c0FEEDiaj+20PSVwKaUgYn/904Fr/+rFZCdYDJWa
dthSodJrU52qiiA2Iu0egZWdUgzP6AyB1tb0gbMwigFgYIPGNw9c+TYcApG8VhMY
XQzI4oHIoNV2+tXbIS6ajCcbYzQ0CVKL/45r/+/ElnizretF9Ui1xj+3IqrB5jzu
S5K1VH+xgpmXTtsmdfzzISQajRGSkoqXzIaYEn6fkyrz7MeWWqCrNeaWAqVyEWTF
JjTpj6WP1WiHAT8BabU+GdFNOf9+Wx9MBl1qbo2phhELa4vNS37GQm/N5rzlN4uV
+LIPJr0k3NjPHJllgUZAy7GT6yVdfDlklB60vPyJ8BsBy7NjxWHIc0zjP00sobOn
DCIlUIuVN7oQh0jvHwrlPFajDKSM1S5kdSnMVoQa0CXA+yAn7jz1xtNIaafJAJzD
xPGSGyPpRVLqTU9dI3nWd6f8QsObmt+ObfAfbHrFGPPNOlzgUQOjjhVIhKluHQMp
1dexs7Aa4YLH74edPihXduPQf/wzzX8lrPePVRnscRJGMM3MlAntnmHJyXaJt8Kk
4Ttkp2SwjrAP0QV2uHLvzc2GX764NS1K3RKgb8+kQiY/yEhImhDBHueGCIE4rFjr
bS8SIe19pk9/6Ak9+jJKyQX19ViyRwFiy/vGDChKSQfogTsgMm8sswzG5U9cc35j
NHTgOGPtmvCTB0D/DyJQRJV/pJq+1Cfob4hcCDgro8QD/XhH1eT3E1z0dJz+uFgD
QegYqdOCysJd3YJIdJZCD0BGczZGdwI/e/usby2VovLp5VIMvTUuLT7lwnolc04D
5k9EujufNRnvBgzFi7CXS2oOT5Yaf1u4XScv/8ODVYCr5NhgBwPoYuZcuqIZ5UZ1
0pULVxJ47VuXnS1Ku7HlNpAUbkkzpBGAIdt9/Y7jcKNk1euQTI6/tLJ/XgdU3gdK
rC3lM9fLTvFxoKIzdr+chnWY9UpDWbrXMbSqBuxT+qZ1UvwHCpuFb2MCEIEEmoit
/vdOXNfOErPIn2TzjcF8Z/aEg0pT+izM1hdPmleHHU4mdyu320TpccyHFRzDFl8U
l30FDs/ydvGdvamaKX5BW9SIJr92cg0nxzObkKH+HZJvNCuZvNj7CuwqHnk0pcrn
g8lyu+AFQgxKi/tZkjvQ05b2AP8Hu6D2yd4UD/VA3BT4d27Rv17pta2N+eMZ6gVW
Lj/P9l6bHsc1gIhdB7WSj65yQ9wGULzl4asL8IH9Bi126A6VVEaJjg/2TLgwDpTP
PUtSsGOgDce+8HWCVEMWyMoS0JiZdpcuPd7BijGswKWisjQZzzrp4Vw51Iu0IxJy
IgBGcdEVT3RT+K4vsRoFjTM76/T6DaXVq7rCa2IDzbnxaujya5sHXYPmNaC8oViI
33pFJ0s09h9Ej/L2LiLUcx4vbfegXu+bJ6HPcbxCRvHVyILolRiRkiQR8Y9EKp5v
r7DU6NOHX+WD/rYJHCexYgTlqMn0UO2nRjj/t0goYHK87UlJj26h+mL1qqn2Z9D1
62FOn+19shestuaF59hw1sDlIJ/9nBh4vQunlcQNyKnCZY90alQqkUbPAsBJlLKZ
8K/hbx6v8vJuusiEDoEQsxO8S3j//1ziVlZjjmqqPYP5yz22haIXdB8nsM1d4jQB
kN22MVUF1vZiQ99OMpKwAP3Dj8KyBb9WCL0PPuftRyTRAbBi6Xp0lIGpoVNO9c7L
tFU0sbdQC3w7oEtcEOwKcRP81pbNoH2L/d1ZpfzJPy8RFBn73/3raqADOk5Hc/x3
pZD6IwQQapzSMod+b/kl5y1zPRK59X4dS74oLe0cdxHRrgWoeBnWOyWIUOkRswnC
8XsazrTNE4Av4Y+osIxalWjPUoiPmlFoYc/qKNQJYUy2mowoO/MBEZCNjzirHR+Z
ZGyoR83Awi2JGfZC3SAGyYUd27LWZaqMh7FWTyLFI6gdAOGB/V/iro+u3JAjTCvX
zDwupbXxuqccSpL4HnwZz9d58Lto4bA0caJuLKyLh3V/L5csi0wjyVcPdVs1wpgG
IkOd85NY8S1qvUThbnq/nUu/lhFk+SBZO3XrKgtMRs4j/wsXPv74+Koe6c3q3gUZ
rmYvaun1ycwLKKXJfFk23fld4Gdxyk12fZNBNXVvikea1d9CARUjo74cpUl0PW/Q
keW7Rvo8dEcmIXca8i2Tx9wwcLxUd2JYVUWB/+KWmvTJJUbVOW+Y+HECz5blP6DZ
vbW47Act4aOTA4YBl3PJdIXmMHMhqn4GlJKDsYW8cgtJQ5mxXq14y8EXe4n1BBig
tC30sbqSeQlaSUhtC4Vzt2C5a8J9phTpXu2eogPpHuor+ZD0qw7uNWzBls4HGgez
TMAbUep9KFEO2yNajV2UFx4FDRWZi3cqnwHaj2yoogsNo8kcPheRKTHSmenY7tlO
uitpNEafsGkTusB5AJA4pGys4FgLY38H0a29YOi70Dv8VS7vQ5tAapDW6BeLNJyZ
YL0zxjNBXvC838tED2ravfvSlwl9xA/6hzZtqUN/b5PryBXm1vjhDr7shz6xiLc1
SObc0x4FIQ5rLz7nh1FwNR+eX+uezofXM2ISZNakiLcUEvVNivqyioh+yxWCxDy6
NczFxlwR9CO7VIHB/g8+5fzfoM3yFWaQ32S3xK/PsOP9loWlS+lEMjrwfKZhxXSi
7/S/OzDddxkcspwouzs4389D6HA7XnPnk6raIg5b6aGjWCmC5JPv8cC72KnCj1d4
dtYM2it7ujOS9T5JO2f4LRpj7YmXEqiChideF+cAy9FG3mJF5CX1vX41xVjKcwEo
b6S1cX+hJAFfvpaWA6BpSIukGgliyI2xTAJ61nYsIiJzPL6evO/o6u++fXQkmAkV
G92rzMMuiVPuPrlfia5PXsWYcZLgBz/CSPLz1CcHL7V5IsQDGhGAmlQIUxCntOyJ
A93VTJ37GSRl16sixY+uid1A4CsLzk4qPTds2Q2c1k7sRUJfiJzClkllukPqAYKs
oMaxyg0DjFyrs9KcN/tMx3hidajsTgLiOt4j5VaqiEVGrpctkAeqwStwBNL3gII5
61uLFeOvGrDpHGTu3RaGCDwjIok+7t1LfjQ9Es4y+WqjeCxmC4mQfUeveUyFkxhP
1H/Xdm+gZfMljmBkwJ4tjjZatZeJqP1m6MAFdM6xFFIHTKosZnyM0/6P5mm47X3c
XiZA6pQoOGd4BiyghUxp7kaaUV3VAjutL1dzz8NbTC/jIGzqO2JEL+rvMIGv+m19
ahv7PkT41hKRL1BL3lyD9ov42DGtfM9fKdqHBkZtYGp7PRgIpoByNqYtLIjwR6gM
Evg/9xKD5S/YqNYV9qrIr+/9Ns9j9sk0Ze1XdN0kVin+PWyeBqFbNCB0g3JnTehc
KL3lsra9r9ZBbiM6AGA22vqHZs+nn/0NzPDC7O42mFYBIgMIRB5lHxd5m5LlyAXy
LFLuAtkFIEApLglfVCyWQDnEiQjFwkG5rXsIiVi230Sp0zStkr92dEuCIMD9x5Q9
RvdCOvG6vxyngcpwEQLjhf4HH7yFPrePMop9Py1/0LJnZGbHQ7mzeDjQveb3q7gf
T4Mo16swWz3Qdn4DOr39wBQFvqsn+hIElLqYcSBOKIyEJqGXfHu/XveCt/ENhnHX
lSjOxz7Fp3jY8apx4w7mOm11Rdp2ZgX3an3oe6IuCg1TVr8rhfPzYGcR1hZZa5PH
VgzmmVwWHMxoFCWOEw6bwSpXM2yrIcaLNjB4mc9e3ENgBFpnIQUB5zcJdifVSV9d
CRuOC+QoYsFtPCpw5nmLjpNBXZ+4iktuY5eP9fwSD/9ALm5TJMDri8gWfoeXo1xw
wKzaqGPO41QTO0YTTYJbSKuLoFakMOL4ZNQKOka6rZB3AjNVwTgKHztYHgEkYjAK
UPjF9VQNaMWU5TsSkvFV4jryt2T+g46NUXhw/KGDXDhQehoMwIP+4kqNwLFv0KU1
ES+cdAnA4A8qCALbE+rfK08dHSxe6hBKPqWzRfRo8N4HxNQTVsbeCI7C3Xp2/CAa
FRRRhCZ4RVJwd0YppNVJE+E3K0WmHHGyP29mJwfIVyn90f3uCpAdDzU/iusyto5U
xscqQ1qLa6IBE3z1/YF6NMaEylYaN3nRSvi2pP2YcoJUUb+oBCs1J395ql7nMc9e
QSI1kxdlejYH07wWC2U3N33g4I/vVVJqExKTZziWvHG3SOBXWqGhpWB0wu6DHDr8
o71GXIN2j9Mp3fb3j96689/Zfj/dUn79kM4HOOPBbGdzKC1b4UvG1LaY5iM1/rm+
dL6Ifje1fdtxEb9BCeEwfxdNuMM3X8JzKZ7P0m6F6nnJZ36WdRmOqoJLHxEIeKcI
rUib/LFa2iDD2blqaVfcU0h78igRI66S00/+TLsnd4ZA+N4OGmzYW2PvUIPvbGE/
ZFXu8hs90tFU61UVkpNEHEGcEQnRQ5pS2QimqN85dwxIvgWo4NsE4WajZF5OBbXj
OEAbjO2NLkQBayulQT6OhNzsyBV3ELueVtSpubbZt3ElO8/S4UhpAAJ+SatN+n1n
168PV7l0L52ozrt9++j2KBrSJKJ8GH88H/SYI3ildOZWHc9EOT53LuVllM7Vcq50
ij6qrLbgM+C5E9ELwC5XEWMw9Ui1F+fJfoneOPSVLv37VHE2EpdIHhqqRERJBSU5
QApRW5mD3dV/VsVexxslPQhlZZPX8oRQQ2DkO5p0CDath3dfevkJ7kiGDfKzrpsb
ut0Y5rZs4yn2r6UPAZZ7Z59wmRXnFJgCZIPInXpn9yQYS2kttGknkSnahWh+Rt+Y
+QNTmyyjA4N6xQwOM4asx7QW3LRewpppAs6cClW/wYuWIMosFP5HSu9Do58+5LsL
hCH94tKkBRDLdZfgsTGJJ18ckv+qyTEUkafvu8CKuZLQrfYRsg6/4Q9egScit7mf
3f+HeFsOpJyujXG6guMl2B6RABw7byFQuGPbDRZgnye1Z968DmDic0p0+JrQnfSm
7se99RTrIXShYUNv944OnHZTRC+Nd1IlEM6KTHZjYBKDm8VTJFxgrn9NftQAUbXt
AL724CnlZctQ3MnhZoPJfgeDEgNksMYjc5rSXmNl5GDZqSq+VoDWv/lfmBwDQicn
NGbyuyidgTArhzcmhlYtc7LdxKQ6E/xl7EsuBWFRWWleLER7iJ/kFlcCjxFRiD5Y
uEHtONubKDUV64GYAWM/nNbrRSc4xPof3cqdypQ+GwwtUd4Ulok4j5SkFgOM+k+u
bJ+LuHWbcEN0jK2CFaEBPT+jPcyj8XABujk05VozHdbi8k64n6QTaVU64I25wBE3
ohlkl95vDBeyWl11HCiH8MPQ4T288WNH1oZUQYIxNbt6wOQ6acK95QUflWApDENL
pDmibVF5bnEJZT6Tq3Th5p7Rrf4kWjydajVq863J9HfAfukTQ1xv306O9RpcAx1a
3+RKNQBocg7ocM7mZO3m8Q6lvh23NzfZgJYAWBvLsk/AC7rnVxeQ1YdpFa6F7CK9
3knq2ggbgVbl5d67yny5mlOAJCpZ9f9EnpWYWiC2L4r8jl8sVEA4OO/EJapkenw/
DzdWRK+tI2Yf9M2FTUomH37mtu0hpTGBYbgS7ObCwRkKJEO5dE6RFNzlaYOWqHvI
ZkEUMzeGoJhESuW1DaY7upqSsI/RWC/TkS6jl4m8uReBWH1Y1oviSRdF23CIIHvj
+U7Eje3rKohelR6cETuGofoCFjffpGuT14awtT99SwgGBOy0xEtvSloFAScYoxqd
I4MTOw39rYnhl5tHqLcu3o8IaPxANJvg28mCX4OgaYyS7TytxMEhwKfUIyA/K/Sh
6xP5Si11CIF3AgligElxGq8Qzz7dmwR/Ql5UkIo+xqwqB/9t8gvx7sCFMNYRlg90
TeqIK8DtR1X7hLQOJ9mLtF2Vlp3qQBI2XVOC8bflpruyEDjJMYpUJvWB/zqRwkaU
PM6aFVTO84ZuI9KtwMIbCq4B9RqRsod8+YEt2N0/IWsGuLGz0D8OVXqtOqMnNH8O
n+RYYrxMlATycczik1yyTpljgQXYfXK/55GXLg0f0Q8RDIJGRQPu9AhfKnB+TT48
il54u74dx4kExmXIp4/RKo4fQHPJZV7ajqJN6kp/8JF/n2eIHsWgf0orchR7X7sX
rcSxx5mD8Otq+COwcyiYIpGu+QOCJqMykqio/OcEktpnX3PGO4VHMmdLW+iJBTYo
UuP+jnRz7EX/tvlvSFDgCrbyjzktCRD7315TIxfWLLVL9P7vMSozdn+xa+KP86Ai
gmtY7UGgpKAxw4gQPf1aNA4KNJjiAWnte7JU6QOWoRk3inbDDLJYGc0bvcLbyn1p
RPyY4FUaHyisHQRTXdSj4FAfDXEcor+PUzafRF6dOCEpO03ryTev5KQHF/nEAR5p
QcPdLQ7l5vRlzg240OIUUH2Pyk72BkguUxBS3NgLYweyNOOy4CmrlaxKiUKzjVbG
YlQuSPd4BwSr5q5DGq8So/pHubz4gHi5TSsGl8dc6TRw9kFIpa3PikOT0J16YCkG
wGiHjgzCcREWT/pmGbnmGDEHZO/8MsET2L+iPyTG0ATUwvIcVuM0/CXzs2cWS1tf
EJtCdh1Xuc5yyhptxiemwimmPB3kpnPeE6HYU88H6xZhaGIjP8ImS2a+Gab9ybo0
fqptfSh/vDArSOeYM7PJ1yhSrPThzG7t4i9pcJZndxm1QnXl0jnc9Y/UCYt4m5gL
WjshqsbzftqQe0mm5b2kP/DPAKRzAy/iccMBJNFteFvi/OrEXLyKe1QouudpMq9x
BCXbhLaERBFS+IsaJG5GXKONjCrkUq4uTjuria15jQ2oFoUFHP3iFHAK1pEgb1+/
oli6vQxCSgIIhOu4MISUN8530xSeuXRBEGRS6ydPBM5sXu6IYinsEyrLC91d/2dG
9KzlBLGw6rikzOeDF24SKPFDhw3q+FXubShAYSgrJnaZ+aLslh75p4z02x+qiYVl
dALJWx7Oxr0U1ON2p1DrTaSgm4eGRGLysRKuP0wiO6g+MzWCaHdbZcqEiJvHb0YB
UCz6jjFNCRp9Bq5v6n09hIHcRt6fI3X6LdhIkXqzTiUyWFSMcarwdwgucJcY5NKD
j8AJ1VG8z2zlDC6N4XLsJU1i88uio9ctWaF5yMDkr4ICKdyqOGUXR2bKF78bDDbZ
YLBCl+6wbavy5ZxrqfRZ2MtWLp91l+2+IHkSC0peNBo0atd18VpBy6OAoJqzfo+v
O4LWyF7aZY9uC2iFsCSBu+mdVZ1LHFK2u0LNvXu5ZpLp2fxOdQU02i6oqWepbbmG
dZ0wJzPwndV21B47mty+5aPp0N2h5XB9BM72CK+6EXFot5fu8Fu52qoOGFgtKhj7
ST0XnCqz5RgR1faSJNRPaGQVVdUnUz1AzXh+Yrm07MHJx4ZbanKOgmAJMp5zgcvN
gDB26PvfBEJDmRUW0eBxdQNUWMYLU0ahnOhWJPmlpaaufTIYHjEJY/kbb04IKQWg
dZ7a7W5Su/NavxoSKSa0RCwHfxFLdPlo+41t0Tm9iiDsPzxlV+Q49qUfsXRgd2qq
z3MOcNsHZxw6wrSGbaXfg60ozvKfmjdaxCDWANiL4Vf46mM+X0HS++RxbrhX7CJd
LFYHEpbw/xiekTsWv7dsljX7HKzHNJEeuZ7jU5XjI/FjYxleYtr3zHtHpZCPx2xc
YRDWJz0+sOBnpIAv8NYSdLYhGnedNornQm2c89ovoHW2oVafw6KmKtQSRnt/y+G6
Xj2zmMfL/CCZK6mcLjIh0/pwRrrDlbOfge8Qwp/d6RvLydsF5wX1umBlUK2IFR4Y
S88dfcrFX+DqG43BYVFp+BSLr9uRLPIimYu+DM7CI9C8fDk0wrZ3egi72NVe8Ruq
eYBhrymW24D/ygbUMA5TzxeC59FUeVT0p+i6+S1jGYRPC5lMmPkMpzTg2BJ/fizm
8P6CYteQWhEoQRl0zQlJaipnRXf0bfzsr1frOsttJrhVFwDWC1yALVOWEa6CMWQT
/k++5IVvtY0Ea1lpKZWvlDxtFFf4Jwx0SbcnMjImfnt7kAgtHocKnzJRIuIfLzHe
0SyDFjQp4HaIK8ycp6/2Cx0/t8d7HivY2XmM2qgeHfj5/+S8D3x6VmT3bkJcvFa/
6xjNHByM4E4v1AoCVs+DYXc7YpUdsXsc5U90s2+T3ROAbvC49GF3Kqtnqevi5Li4
XfO2ScwVakQf6iICI843y06RpiQldMsnkwNn55t1mvv2lYpQN2mEp+6eu48YRy/T
6Ug9gs9FkdRMhqZKWQLI2C1Xo76ZWB1zMcVRm1p/YqR2CmFa8dhYTn2g/+MPwwKD
GPeYFaT53I4b632Z8kLYicM0vyov3GyIMhiIIm+S0dfPZySlmQxXjCTULgPJsn0R
IS2V5RrZ7nOeuEasfG8DKEAn1EK9gPdzwTKOVyd864E4EjFuJV14FMAkrlrgPDMC
YuMcLev9xA9tBDJ76FwbWG75s3/q+ilYDSEYOToCLM199OtvIPJRcUr6lTVHigcR
YA9KPI+8RjAQsi7JuWqSLFyjKEpu6XRlgNTINPmvKZH+aL7aMFWEBOoIixY+NbjT
mxSfVAB30xAKC8HbjxFHE3D4gZFeO3vWMIZRtCTHB77sUVWor89d6KmtLQ9VhcNw
OF5MPo5u3lCWvQJ972risx+hb50+xbfG5Ljz5/rsR08KI/UjoSW1KVFB1sAmtuPt
aqjEccyVZnr8afVcHG9bLtNyWCUHPsXtoB0nVcM+YRtO1KYLsbiC7r5XK0GpAvRL
yde58DlNW+42Y5eGz4S5N5JJYtbaJ62f0FP/9PpoM8dQp3aKuKFiberSLTkxwRi1
Dvr18Ty2jBUc5Dee47yKyOZc/Z6r+/uOWfkhLV+lR7nqQN1IQjFXlOpZZEgZdnwa
Zyjg+W7DCgN2fDKeuRyouIKHKoMkenG717Sc6vzQTOqTgnBp7pneeQMirIU6SPYG
Oi2K2XcBRANydU7lScv6PONAEH7MsZH8DZM/CesFPdcodVS/3xKGF049Sh40Zu8F
OuM4cd9oe+JU/E1S+QxmPZSDjy4VfgVLVCLTw1DP8roiZ8+aSBggnotPVnrO6skF
Lfh6Ewy/sLAUb6tgIGrUhwUSbH+YrX9mxA9mh4qetAri8oV0fxZSgoaqycaZA7Nx
d3D6RednMR8jhoeSSK/iT5s1RLdRL5ART51vOiVoRCSxGh6uwbgZ/no1iCqgk8zT
5CxfMea4EH0VNadjhtwlHXOYbX9gN/sO67n29tMqXHiYFe9KIii7zPVKfAnUY4v5
cxW/PySQ7afhxXGGgu0srP824f+5chgZccc1MXWSA4N1qHEfPFK0OB5N3iupRXgi
TQsKyXrLWNqhWDiKFIfIUekiL472iLKqtUnmMkDG+2EcB0sb0irADow4AdyrzS4T
86ziZAHqfAFcYTDJORqoj/EPI2YUlI6WzDriDsFbbDvNMrZ77xXSwaY/T3yfBww9
vIa/E7edm89lZhy7V2LRNrF9nTIyYV4Ma5w/gCMty+fCnUq8aBrvc1en3LHKijAT
/tJIT2Uw1IkhU7/LBZ0X1zwJ4Zutxk9wmBUz5M5IyMMRxS7Sp2A5iPB+88e/wuw7
htpqkqmsGnnL8QPS8EAK7a+RvJ6GJRrcOhVwWik/UFwZ5fVI6Ce76sdRTRQq7erT
zLvBRj8l81peTSz7Aw6Rr2b3GLl0+R5+HVip25flsztsTvt/S7ba/E1oeOhhHSce
Y5L/y7SradgkQNpOQqmXNlhmt+l9W00A1vjKogdCKCNL5vZu8oXJeM8Qgey0islJ
WclwZRKu+b9imM9TIgYgSfA2WkNnP99M5FuS6f6Znn8EqOKtUo42r78MU3tJzZMi
VRR9guFFmSshv0pb0Q9pMuI17CQba+JrIPxSyzrvaXs0mynb9DRQOK4+xVZB3SiE
vLRRWUit7zKxmQ/kF7OTbrzduvlW9R3/QjEfYkJeE+ZhIEAuBruaXkA4mM8l2Gp+
SIPi6UfhEhRsFXcBt/el4bt3ei+ZOqgYMOxtopq4+xlueR/XDqRfKI4hx6PWDq81
+J2gFLbo2ivo3yVqoPPZzGIWDR8EXS4idINwcVmlDA4ktrdnD938xxzY1CZmKzS7
el7OpR9IM8igsVSugUWSXYB7wY03T0+nUVxfOh8Z5UkAs78+nPC61d0jLpi9/DqT
+Hu+cLs047nh4flSmBBadnwQYBKbGRwKaQFBo6pK5lkBATRgLJ65y78V2gQdSixI
reyR9azfNzCfDcKTp/1EqM2t3OIT/FB9ZdIhgi1lgEa4CcnB13O0eiTo3MKIJtZm
IeGzlCG98Fw3Db37xuOM2PsA9utpPttgRcSDRXEvgI594P2WHZi0suYLC2X2aIrP
toPjDYi0u5ewum3Oy1YBMEYTDjbNFMKre92inRzNa0wBZdV5gy9j8YWT6e3KU5pk
g0F9afRGu8z5c0y4V1EjbAqDfxSTxdkEhvtPQSL9l1NbeDJumKrmfoSnne6sQaIX
3sol4KKRpbHAUfEdL65nPqj3B/8w4b3h60z0SSIIWed/PDVCxS5ry9LGaHNdzDb8
DXhvBP3P1HxzoY9yfeoS7DV3hU1x5DSNN4b6wZYaBxnrXT2pwdFk2UqYMLic64su
ZPKSHXwtejs/BDPuCBqE/RJHBg94DZ80b/X0I3HBvkhyynAdukUeRpY89tOzvs5w
vdv6y1pwXoLGMrWTbZIdjjniQcrPSBdRrKoPRIOwbYgXl8BM+p0Kolayifto7veR
CxlEDgf/4MVg5E1Lg5UVg3hFGcsycwSPvofCvjozuisLSzEFlLZJe08JXb27hYEF
Nwk8gkKy1G30JUG69Zb2udpqtQkRWbRlx3HUPRjoCpnipHa96jTiDL1vlaGGU/kd
fK97urbgwgZF6frSmq9wDuHUKlxsGQ7kz54NeHUdNJDV5qQf5oFGmGvsxrh1uQsi
4UfxoP9GvWDlt4+TsWBMgryLdd3qm0OLbkb2DUYFCkHlDRDZNpLRSTL3EEKMJUyf
/Zqh2sgj8sVLsxsBGCAzZWKEGJNpFJUoD34ud5dd5UdGAOZnEf7bpb9AG65+GzNw
DU8/+g+MZ/alMy9GvdOO8DMeFxccLCYVFStu1NBdZd2JD5Iclk36ZYXC2ZKKqic/
F7WOeKEn38GtJDIqtudEKH3cS4MiQqmNxUHGY9Lykyf6oE0xWGr0fDHiveW1plx1
XTVOhUnfZw3u1JCzAE5EsCduFW/rGoieYhTF+8iV34YBQw5PsI1v8fxs1eNt6AfI
x2X1NDEJEzhdcz7Qw6TCThJc+XzCkg22UEF//GwB+z/mvNBoZHbTLaBbug4bKyHH
JQp52COORdAVblTeREtG5tzT2Q4wiVABH6tYFZ8oecEGdggU/mrI9h2sCpTWiCUo
96eS22dPkOp6RHKCw98n3o1ccF6052Y02gYEw8KBuigspJ8orfzk3XcYod6TAUPq
qEougQumfbtYtSdFcHDyLXA8ydgWJMC0w2UgJAxajbgj3ZZCKDWMwt7FSbLYe2lT
Ky0U29P6dhYCef3GPmMwSov5mWH8masjxxEEuODaD9xnWISTTkbYAJdUBg1dQzVi
uc42U4fIA0hw5SCpcGb3edtaPtqmEFrIodKJmtgth7pA4kGVKwkAfiUK2rouoLw2
G56HKnnQlTgmkHGUJrvpyq2hhaCJihDVS186wmVzSbZU+Lefv3iN/lQHfGJKm7ok
Hr7BxEQsqv2cR1Jvt+3B0GXdT2jF8l/9A9jIuIGQIx6h9NYfQSXh471PWGO91aEd
Ko+r9e7Iws55avRv23X6fJRhzI1iutLPkx7PXOCHHZaWsOpwwEIEVkEaumh4aQnM
ySCAbbsJm9Ix0RK8HfZzWUtwhvwWqLpQYrsyrayl7GXJwO+TiiO4t+6SzsnmzBfj
rmui6hoM6kXAGLyJuALdQ7BaA2bf+ca2Ar8gwsFWBb79kVaTs+mwKf1oKFvUn45e
wMgjxT3Ns+DFxUKlrohmuFTo3t4G8tdVtqJ3QFGAdwnVKHQk6mA2y/9dy1mCsChe
05/fG53X7ylpHe3saQI8L4qokWvrClRPAoie1NdcyqCEHASbVgBMgNKLS2o9aZYO
/Mny9q2bgfE+60M6/QKGuVbN9/R4pxPgxFXylbrdzNsvrcxChKzeG4NmiADM23eq
jTth19p85K6d3RehfKyIsd57bV+ABT/GmwDjGhIbFXWgKIFT19t4LPdsB0ApjeZ5
46bUJl70iOnR2Xj3aBuiblGj7ViCFJ+vcGbOAsp6tslJDdwz6s4rXE/2qbDlDP3F
X6829APxsqwd439eUhyQWHuhK8dK4Q701b2d1Zt9hjVaG4UOdytcSUrIWJy1cw5Z
9wf/6c0hVgipDWS4R3+D7OUEZX7L3IojFvf9IWMkLJadgJ/pt16LONfQps7/U9PY
L8GRVduKolrbXbQrmBSb869rrk50hUvq+JUglZ5et3Xt5ZLi+NMbJ2P836gTiUKn
+hsx8YgQFIY063WUGujEKSX2RR6lbQKAry5P5urvqw9LFfvXa9wPyNsphgoCQ1xv
NuEraGdlu2c/PA4173V6C/6PsX7zLfgmGjOq3vE0uqFnfcYzrNaODbrV5Sedq/Sb
u1lGGszflbl2/4XYga4XF5eKXMi8FPuBSzHQ7I8BTK1VfIAoU0gx1pV5xvXU6Xmk
/5S8AWD7nHBPxWL2LpmHwWg5ttOPg19jAHJz9JGYbBDcdZwJKpcA5d+IEguGooU2
jRwZs7eV3ax60D5ufSiVsaTbFTAb4yIoWv5KdThxfbA21lZJ/bPMeXvENbO1tPet
yCdr3TsiwvpIoQ5xW12/0MSR3e9dAXpUUfZLQBnRrlHz7FUolkouWWcvypIu8PXO
uV5uy3qPJOOkS+ffx4xMmnFs5O5kMpwys6WgoCs8ZDsNqL1WLsxRgsx0ZtAYLQD9
clutQYd1HEGJfsyPI+iJl5EEAA3W8xde8CLejLr6OuqRVnoGlr1UJmHmi6QDjS/T
Res6JJOim1C15+x/TxdverghuOyu2dJZ1ESBAgoep7q+PEor5WqnDRHnTPcM/L9k
19tX746XYTCTWdOh4Ap0JntGNAS//rLtfEFi79/8JrlXWkS6CaYOkiAAWHsw1osE
9XAZhORswWTbZl4/J5lRDhrHlMWC/9IwjjSr7D06aWOdYcP6jTDDpA0cI3TmDXa6
QpReAe4Oui+0s7HVL2c2i1PFsgUkBbw/JbVGBudrlGU8H4QPH0ko1dgz/OwMw2Mo
lwy1c9qk+vXDRjR1gxMx/O/4+sZOB0HtVzE+T+gacHxknICQqQuuy/avkUPm8aI7
PhHC0r/1ioFed2NgObHXJIfqVykQc/7/M5sDzEzyD7PsUhzI5mABp/A/kV3QRw9a
MRmPlCg8sd4MfaqAJc+xj8TNwM0/YktgAc35C9w/p5K1Bl5Bhk3KLC4DN7UlDYL7
zb0u1re9tWGlHAdnWvDFf0S+JEqPpcxwWz/HGnmRvvjuzsfrx7PbOORsxNr72Zsr
xGbgpc2Mfx1457948zCrMhaNLWCJS26Sjb3DTsoKaaX+nuIIOLVxRGDY18JXCqvI
MSUkSaDc7O6ZEIsg+OFXHvdicK39paQW6CczGGV5LS0PYt06y/ejgaY3+zUytptT
E4GHfwn5BKH+w6L75WUj1Xi6f8QRHIxS9aGN1m4qeI0BMjHvjvovwKxmVVbQ5Rpo
BAHJEwqtim+1MNLjGzVkRJNOgOfFQizELtUFcIcy1SXMmCzj9U9JlOed/x/qNBKg
M+8sOXuT0I+btMk/qlUVkwg7WK2K5Ch01Fa/8qLp2XdC9lzAVN3FKHfzwXVmBPxI
8dG7qHui7ZyShhaLtbKy5/J4um+nZz3Dvspppc2p2DBsibMkYQAQBpQVTaVC8jBl
6fmB3fxwzhjOJGEXOHPyFJAFgGEy6aMGo8yo4+JUhYaGUkBqTIOvd4UPq0DXKYP4
a8165fWmYE+0PoqOAyhnn5KSjEOqgqNPFONmfNJ5/tzJa2F/bSo7q7SK1sPzSOry
rOi0fzPQyYVcRYWlZFh7Ta7mqE+/47CqWZ+LO+J5y0YfTSMB901ya/26Fb6wy06u
KkLejgjD2snwQHUNp7gn52sq5m3kLUOu4gWvURbcnpxu5GusVSZAaFYAh8FGhbAI
DjNsbYHXhpsbPmFBcanZhW8BmRiJHUW+5ywjLMh9OK4tOWamqQ9KMOlTyNIDZGW/
4TzPxfdkWLu5Nya9mHJKFqGgh0Vv/WKT+0ydS/k7kUML0Jw5t4whnHDY6mD0t5xz
tPxwKswuCA16fFcnefazt8MeJ+17xHyfeh80AN/UyIicuAJW2zmtQ5e+lHpP5gDb
fhY9pAnC/7PVK23wFWzMIc3fazLjImxyQcU2Wx/qC62k0m9FYPFwg4HWDQicL6mo
2DADqnrNe2ezp5fsq7+DutpaYSNO+X21D9fRsVSkj8BG+PLx449UMFx1+Yk5pxa7
TtEbuA0p7l22xQrmGxuEs8KaVMwYi3SciKydkr/I0ZD9qwWx5C+74E/DeanV1DR9
QY+szeYZ6sMSSy3ZEwz0Oujbk+FOMwbpUKu9tPgUJGRAXDYWfAdYsyw8FScEvqr0
a3GgB6XQzDeNANU8GHNvibS6zL6SJzLupl09GSm9WPc2MF5iQxFr8pNT6/E94i/4
7+6aFienWj+JArGLbZTSlD1W2sc8pDUoJVn4T4L9b+uISRDIY2URDejnpdgNsbQT
myfMXZyfHSTeKMT6uAjsaa/No1NKaDDQ6Ug2Mw1WbrOPwsIVudY6K5MwXfIEWmgV
t5FsQynWTFLXu1tsAiwIGv8xfbk5Lz+j8OSZ5Px0rD0JqeTSbC1zfgTqw/41KPAB
aH/wy2pv6f3JBVBQJqdqrPv37lBJh3XkQGIf5AEbvl7DsWSXQUbVp7poXFXO1rSe
QiAU0N+ASdQkrKv16wU7FR5asr0HrQ5iVAB4P+UVI99JvGOGxtgaSrIBhc6M/W0W
nKGCJ/AQ2SnfbwgcVi0Gn6IbFIc2TgJ4udMr9BBbguk7oJdsZn7fOwN55uAz7qig
piKUFdcE/ig2Uu52R6+TUgjx6oLVouzpq7gyGfBgFXnGO6j5BrO22vZ95OTBNAp2
CMFOPJGk+6zOr6wLMMsE5a1Qg29b+E1FJ2fu7X3z1X+G49gjKmaxy8n/3vfUAosZ
wdTsyg1PJsUMOYFNFfkTsPwL2C+uOrqFCMOtjImpUflSeVUIBQ9236FfS5jTjdMd
Xt1zHFv6b6PpVNOfjYnL4IGsjNZ6+S6OAn04yot+Ke8xZ7BX6KiyDRaXaWeIH8n9
I3ITYe9QeNCztQaf2big4A8KnUDXd9T6jXUceZc8Sw6CxaDoztYRxcYxyg375JDS
N+C35PaeHc4YERCMQomEcEilUbQqIKpRsBoiA1g1ffW2TmCIwR5W1YxoVxjcsXGh
2VoODklChy2sOXmt1kyjUGM9hCk8hUUGqblSITlVg5aDlJyxkV39zHmQylvO4oK3
nCxNIijl0RPUwM8EI/dgPUwA6x1iR1lSlXTYvht0yxWRLv3wR2+Xse3RIDyKaxK2
LL13Kdbk7ug1lstZznIpqzeONfxXGpNP3BAI6/QAmCYkoClEhuNPgWmQ1iRnmmdJ
rL2GBbd8HqUrsOHiS8xOwQ/G619clIatCgzV3YT0J976ZfYDeO0+93JhWlJm9Pvi
XnFfBo//2wEWIMQXm78lVEDRgFnHXKsqQYtk1zifbXbXWy7lJl37cfiPmNR0AIAS
WsmnkHytGhrOMkUiUFopKcpHd//I5y1bNE+5c5ruiZZfGYRNofs97zp0atJkx23u
ge1XNg1s3UTv17Y6GqCBGpXTRW2sdyye+ald5bZRS1Ep3WpfaCDR5oehIPxUk/oj
t87d/Z3NgB0yEH8DnCb4riQrTRmsb913kdLQrD9Ne3RvdtuKtBSqQRdaev/h9V8Z
xlYqgeqr5kfMx33GrkZk2nPiFCfk+OkzCp6t3rt8ETWgN5UUMhqHMhYZ8vyaoW0k
yd+sFvDTIw+LmoNxFLfNBShFQEhyZ4JDjOjNUVuDL+ojNSfQ4MEI8+Anij5jjRRL
zJ72MsJHXM42pWjG0XV+vrytsqEUDl95CiWK1zJKSCcApeR9c32e+cGFB/xI98tB
aoxr6GG1mHsgafXk5Ao4CnUll95gzUvyVljHk0Q5uNgqlYExctGDFnmrbXdXJUDk
vqchazMscEJr3J5MT66T6iIY67yQCG7ym237Y7nfVqxGViZIoetTqZt3bpJ21WQd
Py2nN6E8GBRmiEYhN2lHS7Ju5a3fNjnLvOGgt6ZLwCmhvelFXoXU+pIW1SEmHHqu
RMs8jkK3JjuJb6Fjtqg+lX2fzMxWfxlaYQyfU2cRnKQ5EDQ9TtxKgbQqhdQ/1ThY
SZjnziWYeep29U7mK0J22ZsQmo+5veAVIRK3SsMVsaO0DLLaOGc81+e6SD64x6oe
tH1/3i54Rn+pkpHXcUdxcH1RgS/vQjJLp/7WLItBGbOxZJmppWBDQb062AkeWAlt
3RP7PZdpt6UBhmeFnGUCtyGgDX6kwKO7zMXWvfFgc8e9nySwboZAuFdn/3S31h3i
eLpxbts+7zRoZvjOgZhYfBpgn/Qfrx3rxw6jDi2JZ98rhvYDExemAXcD9esRQNFu
SVcfX54ekl3lRbG/vuSqEXNwXAijvdg5CHacQ4X+5/hp2SgBFNExSq1d+xeEW5JK
tTwHoNIgn2EYR+bX+IN9+xHw5CBRm4K7ZQkp95OxS6cXpUroqq+2qFgogKFXDXc0
SJUNp89rxo3Z1JOKiBF5jAUfCAoYJm18v12QLjzttmd6KdMzSq6XbSQ770CqzfO4
R8LbsOPoAdxIWtblgv1miOedp64mDsDAMEMaw50n9V/w6qrG6djVywQ7NseepNsI
OfHfsiAbTM8B/kesrTWfno9fHt1Bc04zMDIxIPhvBY/Azteh4fw1heHbWKyLc5W9
FLQSKMKwqslokrJP6q8K/N8PozqiNwPm+t2EVk4d6+Y/t3c63N/bxfQFJRmzabV/
ulJR2yxdk3cWkZPk7Ps2Yjk4DJ2TnsIhhnMbmwInF9xj9zXPi/iKhUuqaEg1bbk3
dHey4CNIwtXSISInNJ122pCeAZ96NB1bNzf6fOzuELbTOJbc5DzKZBmg96Bkxz9E
VAg6eA8y/ot94hDX3ivhLQRiskg09dMbEoX0ANUhGzYbgUWiP1PxWu04Q/wT3Iik
BRO3P9EAeLKw9dGlAnUrlv0uiPzWsJ5ESma+S8B9ackC9Hwz8khtJxG+YgYnoLCe
cEfZal+48e4KBofefWojHb8ZPZWZ0N7MPa+pVXdt4/fFSUCrN4Ff8v7zgw9G0dbV
D6xKkqLwiW8MqlJjgVl2tZOEfpAeY7G7qYiQRzPRmNKQSFp2Ir8vi9b6uXoRa/7d
gt5QohwL3nob2I42MR0AD1LLHcMhI4b/VPoipWZNrSNkBM9Osfp05tNJ7odH6UyD
K5x8DpOTPAKOwUHvLe2Ak10J48tZEi9BN5VjKN9mUDqIhwLjs0EO678Habbcm6hg
Q2+TNhgN0mYntSwfiZTaHdBUtMkLbGUOcdZNvSgiOREC7j0dHjr5lLPMxHtWzJMo
BCMzX6eLGy9PR6lWrecQQsIjqQpOI1EKZ3exzoMqKXBhNUscOBvZeqRLLYDpZpgt
OzHvyBX3A60K16RAXTHPcvQi+fiod1LD/1MGm0WQc1PnkxdzPVmbpZXXW8KaVe3f
GQ9oLYPARDfSDUD+qxhkk+UaHGpPOZxBz2rLdsIuZcY8WBcfuKB18R8GM6YXILyy
hhnfNSuq7F22E4v6oJa4ieRcmJLy73GFDT7QsIABKVoMECUESipWemMdq7edRNLF
aPSpRAm3CzsuSQRHfkm2tTmESjhX7mhrv4HeGCESdt0KczXJDs3OtDY2qqmwRGB+
Bl9Zj0aSbIiothJYDV15tqM0mgIBS7j0sH/IyABHzLN1EuD/vJOkw68okK6g0Vm1
DPjBMocLBNBXsDbRqEtPUykq1q2MArRNdagIu9mSweQQMSECxknynr7j111k0AGg
V0bpMWhr2gUB4Vh8mRO3Q2f1vfryJTLIcIEjQS3yQ01mmFNT03dBfH+dhZPpKKAN
qjtmRFKZ7/Z4avadcVDR0O4DWBoK3M8BqmoBYcsn/Aj3cC7Zzh+cCxLfiqhIvozZ
kmhEJF09f4ikGyaiXd4767q0O+NCkYONJKX0m5guJ18sFk/MFTPBP5hDwf1oENeZ
reXsuWtbqTurw2qg8pRlm+xPSV/czi7vhN8t0XAt6/Pn+be8qymNeeIwIlM0PhHo
sO8Zrl6GLhsI4eLh0WZ5qKnlU9KiaNxREIrIiVmWoqD1F8m7ntU/ux25KJdgo7HY
K5srgigh4/XuSHzeZ+mb483tJL7A7Dms90BxbhM1gWlLHg/645gb/ewe1ZxDFLvF
NfT4jcnqm3sBvzf4Kt3QM79r/EJmIXGYjMJraKyfhY3t+SbNZGlux5QCSE3bGuCm
Ji8J/HDOluOS4l7elJine/zNdY9DLno1aROxSjJ4jvKC64N6HyVy6GRlMWZazj5X
LMfzWh+PAXZ4koBsYOxZxTjzK23TZOyRL9ydGDLAu2u5yVLL8Q3fkuRqCrOJ6Dlm
eQmhQPgWeZn3ChElCVdDu3t7ITwxHCJ6Iy1or+2Vy2h5CqQH++In02eqU8clIF7t
h6pQLQngM40V2g583r4FUA9D1Bzep+W2RniiPljuO7irBoqOCPT4nphwG5aCydOU
1TsTa7KS7f5S+QYly3arYuB+gmDiIG5jPrRvczoocAnp8PMbDHAu8gBWv5mMutMU
Wq+iT2bs/9dh1o2UeBCSRpL0X+bMLyDpiZ+dcknaAj9oCtRQQ80OGQjFb4SHtbvf
z+D0fcUmQilh3KfQUDEjKK+STWK1aEY7QD9VM+9Ew+OwLilXFDQ4A9ADsEG5WPmZ
AczfeMiOVZxWSZikVu2uRbPjvz2lzn7KZ/1apZd3HgFO8LSthtWfMlq3LT8qS6BS
mbG5DsJLm+fMOKhGRfERsGTUCTlbod3RdviuWi7Di9iDmgi1mvH85siK2dYbBtb2
wmWXey95C/27KAVqlcm6IDMkTsom2u1Jvas9oECI6bjN1JgVhaf13AfV88Pk4hcL
wNc2es9PRZhywsjqUq4JnmMtnF+CyAuD7QeljE4Kjr1amxh4AleAubRKcHvEua5r
oR1IPasUiFhpkZlY2o6K2hAQ/1dtFiMbRz/xpZbV83SBkuCtv8XMakiG6KsGqimi
jiApQ0xJ456i5K6xcp2g5xCMR1jqJDzwUOMrBvKI4Ka+dp94zlKBo7XXS7VROQvT
WH8pA9lbPGScDUXxLX64mlQ2iQpYMIqzevkfXCjNEnI5x3cvhB7WmCihrAweWoGt
lTsEDo+vpAs+573ihPAUavTzKQhndjSHbTf4Zk9ee37mvR9QlRgZlkVdGF7uVBno
WpCqa+Q2fUb2wzCjjnLot/c5Lvp8XpBkPTNiObq7dlzbg4IHS43X3FmEkrPrAzOb
r/eC7AviPJhZAYbEZ0pA5IL09JZB2kpDSOci73npDM6Lvu63Cjyr6v9by9pPq9hR
IgpTMEujz6uCzJaxuYgnrMTp3SqFGsO3/2HA9PAOGOUny7xJ3HI0GQchkutA2Y7w
ZAxIZJzLp0iW3A0abmP6jLiJUti4AtUhZxhyqoZlfzsla6YfU3WJML+KAvRfkEYm
H7JMeFSMQhoMsB0D+6wtIXo9TllQVRwLmBD5qgvJBPZ01Us455/+gZa1BgXyuKgK
MYPC+HrgKYwlgejsf9O4tlVqOwR6qcHx22EPURQxbTgoOB0NRn5gDRnnjpVmLz4D
8UbCQxhrPQ9i1yLnbE8YVaCDnIbDog8jQY1/fW6aB7k3BCiJO2d/x8SrzplMQR/N
b2QGW0fjSNbhTHScWDG/EA4IZC1ev10W6z/LQVzMgtmARhxi10ZfQnY7VHFbrsRS
hRvP+Bo0rUSr+HBPwDzKZbkRv/38IdEpOMl0ZbUh5d8wFCWW71jj0uM6mwjXPGAt
L4fefb7yiEUwInlnEtawzWMw6uNjTwwZcvLmO19juD77pUdwh4gGTg8ekVezySFm
JmoVf5svxfnGI5JwnvsRlsbi6UZFHqr15Su4xK71Sqc7HOIXqNWgisg165a69ljA
6qLPrbhJ9G16VC22i6Xn7S9H/x1+Flg08WtPpFo9F7M5GlqACWlWQYnPMNB2pVxm
ArNQcXmIL6nQI4xLdeIdaBjV3E/7zkHvC/hAdwkwQ1KqOz6fhPuRDKaUiAiF+3NR
0Yqe/XTy5Sj/+1sw6mutvnx4Z6oiRe1W8lPX5orHofiR7DCnFlP21snpmTmLwJth
OBm1Rp+ixczFQXD+lYckeaoTPqGdOF0dJRc8DGDK5ZxMi8F0FonjWINn9qEn6vDo
gtW51aKdDhylYfqRZtVXoQgvY6WQ6v4rDdMPdho5/OUEMEvnGMd+uWnEBsztZY98
U57VT+AeCKPoTZJ+8Jsg68M/F0BZu5YPeWphybubJN5EP4UbmA30BCnqeYsF9ChB
G5CTfCHwRLvIt+SUS8Hk9tAsiBFxv193cAEljIRlKdlAhPtBHjelLXT2q9dcpuU5
SGrgvOnrDq2CfglmXVf/jdRsxZfYjHHPddqYk6IKXC/jRnYvhJ5+Nsuozw+1M3gI
D5GjaSaK/DrIfGLeowlas3iCUmmhFHkMSO27lkWU+98ZeaweBN52EWdzgvQKPTYb
qK9LAeh3cCjxVZTaW6Fmqsy1HF8A2ATdZ01nSvQwXH3pfHdJXuiRwAZQLz2hviVd
pGiK8DyCCJTBACmjE/H/GveZDHI6QCV30+sKrRz3WI3fdMBSFQkKDygRHk2Ema+H
XY7Jjbl3/0eLJVRMMdrK4QSWtWmBdhBUa8OmMWCUah6JHZENTt1Szuypa1UqGsgk
Eer5MzsrxGwVcawrQEAyO/XD3fxBa4a10RrnegDHhZcoeiPhoDS1OuGuF3P0h+f7
oXQ6IojQbVg9sWwBzNEc+EuC7SiwWFz0PnoejLaGXmdJ+K8NCJE7P6KLX02MYwXr
Ocjm/k+7VQkmWaRSwNJI/luFSjSUJdrtRQ/vulSc1gif53XNO83j6zjc1mZhsYja
gAb4rVd6nukVDYhxWGpteGYLz7U5K7RXgKRhuvUcI+h103XGr2Px2femNM+vxeWB
TXfKXNB0YwHhQUQCqCa39IZ41ZrBDb4i6iQXL/By0ieyFIs4bdqee7zaUGK0zmww
kcJW3f4P3eWSbfEXe2LubK9WPqra4zArqSO1M/0NIc8Qgf4NaiNT06ElCpZTzKce
PQWuHI4UHyDoMlQEaBjbnW+yfqXwJA2s+x6jt9TYRY+3GB4KZ/g20EicWbI3qSVh
2pPofuMOfj3qlIXQyFewNcYeeEYRtOnXVS6DzRulvucQky8heF2W9TL6ZmWCfTs7
z+OaaGWILUEmQpIWnHF8VDzluTCGVkzh9ffRJUtSUJntqoexUFBIC8T4vwSMl7N9
jmGTik2MX3EO0AQ+6qf0PLwZmfEoA+hwFveRfgAkSf5QOBEiEzOB1izPMKZMNvNz
8Nauf3uHjKyMzPCA9zKoFX9FwYEr/W90lAZVVghUzryo9dq0rC6HLZ2oDfPgBNtz
AeVM5FuBnnsWNnXR4PbHNVgBubgf2K6ZHQBdqPUihX+KAN2yxERh/ihQ4C3lNtgI
sqf+7HB8KhYmBm/qBzHk22096C2axQY65UStXOUJwj7GYmwrZKsAkjPgye6pTx4Z
bA8GfcP4mbgYjSkB5svft26UmbmBIGtCGze4pDWj4fcrOW6krHKJRzgMLaZ7BbKe
v1l39iUVo3+CZ/ejzY1q3pbix5fvky06j2DXWFgupfB1lN5htdD5U+8r22GsWasi
8MTGaDdU2VgjPPwjBwYMRtVnDD2VdzQwcrLkkmdcBdtpvix3uo4I2k8RUHI1rPKA
TObLXhFPrLkoAKaILEtt5rk2cuRhydIdokCCo5ogl2090Vkn+9+9n7fv0F17SnTk
VaDGcj/1xJmrULr+8MYkvJEe+15eJzuaJ+rwHa/6ghhWWVI9EMKYtkLSYPrfTLXx
XqlptUSiu9s2iPoJS2RMitCmiqmR+z98jZRNhwY5Uk0mszVawjUyQ2gB5VDlg3cd
Dz+ykWyo86WCxf9Vva5MaiR7wAXy3t5YhWgRlUYTEFtYLL3PcvcH5r9q2oNAK+g/
286M/qnSf0JKL4LxugzlQxSjlyVQaJdrRqW1/a/qtIgc0ebMAYjqk96lzJ3zQ+LQ
YbLQMyudI26vFfGEt2f4kKNK99wJjJ4oSOdeOUJWcHa84AAo+HHkIxqSBMoPNp/P
29M5VgHcFPCbb0xhYC7hmLry0CeCiJYoO1iYj/5s9vvJ2pLTyO34fUnTEFrA2rMd
jy7Xof6q7YjCmmyaTcwbFBWs6bIqdilHfmYRHaoIaIXvdgT/xDTtM8Fpn1TawpKW
FKqLxN7szHO9WT/JoeSl6FZCbOXi0T55kjVGnMy6lcZozTNNNFfnfsCv5kXPKWaH
67SVMRoEZKFOVFDsib4IZqxnoVIz3yuhsg9K4LJVa3L6D+YXS+GFGP6G6fREDuRN
sU1QxOM9UAVz1JCj1n+X0/hauzP9pf5uOv92isXzdlh43zhO96fSUY2GtADbRG1b
7+i2z6l0TKT8Z/064iNYH4n7d/e0Ibtv0dczP7cJ8hNxfSYUCqnuG5gBxhQmKbwT
6p53X1AGo5+6v0v0QRfnBjpvNbH49Lo91YgR38WaeltAw5pnxLORfJ4oQjxR37gc
zrXzNg8JrkWGmOpeiW9BSIGAxYX+vUqn0nVPQ9SJ0b7sR341ORWS03RPzxWoe4el
qtmYlRCuZwwTlOSo/04zjjPq/lZuXHZxlCLEGlcknLHOImu3fX3m0n4P+N5Uro4T
ZKjXURYTkLD4+KXhP1udB5WIWsGOAEnbcNRQkvkJkr5lxB0O+qSYheQpyloeP1vk
bd5IVr2bsWywUMWqLtMlbl6YDV9Wwj5EuN7czVZtNqIdMQPCfnLuMxbqXxoaBJJ2
0umAG3A/3r9dLnD0spKr/U/b7TPlt1OpgVm+AImijKg/MQbJ/CBQoXz66hNPUq6E
ZG8LjV3SUaOgoMertERnE34IBDkvGnDf/BSdT7pqlPO/prgNtYz9yI0kFXf43aiS
L1w1lxw/QDkwoMrWpRE8pugdPp91alcaVbrTUn8b9zQfwcgCq+ahB9/nP+SG++oF
cfXW9KdadHPCnh6nwjaB1BlAhUGV0wTh0QoWFwdFXAo+f2MnYKCns7uD8Rj2yc0N
Mhg7p157IywEh/LOh4vdm3QzwM+HLgeK7GOBcQ8d7C3IO2p/B/nl0bdMhtv0SQhP
k63bdCh2zghlPWDMJePHAPXIXorUiE5OOJaTr4yatDZeL2KjueC+Swux47cJQnTk
9meQBbYNWXS1Y25Un5704+JeoDYAfmn8zQRQLMithyexTKB1DzdHK90s5sF8cvwj
aYkoeUbAM/hYPXykdwZDo32fHiR4tFnrdgiimBUCInZNlaCuBLG30bLDGn9j+jZN
8c6Na9sNOpddNoM9UZ0O9zTc6jJQxlDorLud83CowlUxI7FVL9pwT38JTBluZ2gj
/zow3EMBSPhh093I2ruqLPXIadtDGVMz2t4/YVvG6Ove1yVm2hhL2iV/iiqhQ1g2
oHCD/cZRlME91+Z/kZAZmR2UmcyHxMrWYQ3tNyGlwQGOzg+dWwP0s+Z1+MznnKfI
7A3xoyL0A7V5aWGJ+RV88/SFNDGnLh+oynV6HFytty/9kIUn4avyg0KsauM7v1K6
YsEVrrHXfEeJ4adrhwM0LWiXmgcFATUrE6cjtunf3WJd/M//YwSmLOtqd86cMwhr
15+GoC/Vn+4nQDY9Sxukcl0Xzt4aIoc0OI0Nag2e4j3OwEZmG8GC6jhY9ely/l32
CohOU41tbgEBKrn05fy1UNHQyLEEc7Go+/cCtnOqwHojjXnqpR/Cbdqmvl52WmXB
M5XqkT4KMq9LNMM4cIm6ZexOpLT/2p8xBzJczAh9i0U1JzGr0bzJlQm+KRUwa5hW
KF74estEoQwLCSvMj75sdbRcf1tRtk9Ls9Z0ZAZoHrg5r0zOI5JHUSvyOM/OvyWG
58e3Uk0axRoUZz5jS0tyFDNrNoZFqg0oSN8JwXd9FpuHoaEexBlHfZKeEUVYaGVm
J+cXUKzqXZ6nnZpIdZ8Vr0Zi11yjlmnJOpr6L5JhI+R0aDz4YPyh48/6YVlxxYFl
5CWrZqklJfI14h91wF3vdRYy2VBMKjN5Ydq5tDN0a51Y1NVf4Ls8qjF1P8qvqXAs
aW3mznB1nJOCAikVsKfhe6bNK/rBqb3YndGpIQD45TNXPIW+91lB4dHs1qffkOct
wpJBm1xF7Wh5kZEHVJKQz2PO813yLhzYjrXSqUhe8SUqP/Psdfyq3dlD+faVASgM
oQmFt16Y2n9DcubvNQ/HZEnXwx+NYby8WZsZK39v75h7y6KdeYX+8qt+Saf8icPu
4DLy3C9gB8Lo7SYIraeHEyuIKiEUdtmqNDe5C4fr+gbpKEjxCt2+PdR+F+MaUtgt
ucevganbfFvoh5ETYxI6x1ID0NbPx03W2J7TrcUXwW3KUN2UzMvmSCaEt0OiE17l
AQhtwLlcisw8AHcL9p7D0bXF83CAAss1iRURw+ien/cNTeSrp2nZLdYYdVkMjpVB
jTLnUjeIW/PHze8YikMzY/lvqezsWZUjMChOT9AWmPcTOd8IxYhWKOXtpU+7irxl
EnBRyHcF9PhMYQgQNN5QXCG6IEwCHDpfQNejmdtfaIBiZ4jGodV31ykDj/7WwFFw
ilyLIjBEoTJeuRsBBRh8PoUJLTnNBJ8mR91fIvaTCo2ExgrVch9MV9J9UjbKMchS
S06jgCb0FOvvo42Z8nJwAybDfHUNkEyNayyKJJy010DGpoI6rNSgNbTea88zfnAF
/qSVEJbO3M2LlKWLITdXGxdLpxNwqh4hcRdSgpwVy0ymFSx1pglo5CTvSlmnkVM2
7PoYhm7pH01YZ62rAndK3vbYM3sdzkNwSEdedPt6n+XABT7DAjdmYYFhdgnwYkrN
S8wGTbxsHUa4cwYs9ZDQ/+TrhmAjL037Gw51er6IAoLV1m2iA9W9JvIrWvVnBUIx
bxrxntXr7dhsQZm28aozOdb2jjlo9hMu/5CGyZVcNbjtpVK/+ZZy9viD6el7Unqz
/qruB3271qrcbP2iqUZnv5IUsRZWKHoLn59OvKuarGMQCdJlY9sfdJ9QSZVOiQxz
HQuAlRvxP9qc6Oc+UbkYUPyGIIqeBBotv3FwxktE0E/aMuFwrV/IqI8mFkYKn4FA
EpRX/l3vy5ClXVvFUXAG7bqxZqN/x54idN+q0ucF1AWTcCIKGDHmvzIYXt4Lq/Rv
YeC6nw27FJoXwpB1owBgnabCxAiXYk4FNSkVkdH3vGaRn8UAjKT+WUu4dLyOFUnI
64SXIjPr+JlJN1wb1qynV/MrUMuH/pkNLbdwKmcR5hixcLx4qMeIoMcsMO1HHpZb
YV4o4YzK27nhpVMp/h/AhhYwqQUB3cPJEkxuAI9teXl6fmxcqaeY7esAcV6Tzff9
kyqjRBY8CXNyKZpeMctUwqsDlQCY8JI5dhQqPFvyJKlFYU1Gi3XVRwaU3xeXqDXE
0OJ+//PpxcB9y1uXSSDjYsAEjEbQSxsCNjnw/7GTp/lhGaffS6ghlfp1Q82AWfth
xboAnGif1Kajw+3dJtpyt6g/oIMaKMfYVvRqHtRDHXts1qmoS0gpxv4PBgrIwvZQ
gU65dR4ztHDsJCl1U/nK7isKqMtVYX4RzAywAUMKHgaZ/wAyCRypA/dS/f2x++uj
3f962gmK2IFMxxdDoWABRdcwfkjDnMV0H44Qt2gZAWaob1D93n8LqlWiMDmaHCur
NyBXnMcoab1DRUkO9YRssnaBI1E2CVA4L94QHoPmvZsOaj88FjKyYNwV/O+0zl71
QTlSjmbzk/hk4xHvX+GY5zeBgkZe8m5L5JQYFCB5GE7CfX/CQmHhgDgvvZjMSauW
lQQLF+9MH3c+hMrQLtkShHwBsTZ94m//4NLMOdLTHA6RK/2+SHzI0sl7ddLu0sqa
66iFfGRj+lmH97Y43c/YwUFw+ewNpnS/602fS4i/gC9C7fX5BJEk95ZJ/LFQ5PlE
jTM1waX170iKl2GoaagB6zEr4z/DrByq366ZcunAWdpHzRwwYLGgeiAy+FD7PBgE
uM63OmoVD13rciII78MtaE+0lf6Zqdi/LNDsZufjwP+2aiyqL8/y0lfAcXiZKnXT
4lgOGl28VftwSRFQqtibtClCnowdtYOilE0TC9CmTYVQaulwfgTIBRg3uvQn1k0X
wQJttYYYzh0cMIcDQIJpxsexmP31XJIZfBTn2apxPMMN6Xb9tiHnqbFp9LshT1mb
OhaADvCPucbx1VEjtMhi3vq2wpNPZiJODjaUI9Qb1V8WnIdgVTAjV8JUGayK2Lzu
DoLRKuMhvCV5FJNDiCpYZtdRTEL6OewrrycFDcKoOzyhMsJEodKTdVIlLcM2RqJA
QwYL0L8S6VqmEqTYBffAhXL1+VN6yV8BMfMJizBRjNHvkmEABkeVFJOT8Q9VBILd
D45S9ByRdLtCscSNND3ipF8xXthcmMzKK2R5hkmwHAkCIEnH5nCaJT7LgiA5VFE/
o66694fDfaRQQ7xL5mzhRYNzC0ORWCKkvchZt5nBaogPvDmbiYWkMUuDiL4qWPr5
O6yrjcpLhpRD1zPo/exEn5G2vsyrLN71PvU30WcMizxxSt1eCPbHGrGv7p9T/9MB
4XREF52kfCdntz1KNd5wa9WgdofddpKJxWDu/BCJULkGO2DwKgMmEH59K7aOGBWv
FDbFCe7uCt0nc9Uy5y3/pomk4kjWZuVp5CtOe2T+Q3X/YbP7JEHcKyeOuxRUboE5
DAgT9cJ296n/ladia3yMUu0xXr+Rag2HBhJGkAUY6b80iVgrt47gHg/6BtGXzmdd
KH/OJIVdOSoo5DgekSQN/gHNBp906qzxBnXaQPHuHDW6KiRSKCSl8LTD+Um1uqJN
o+ewEur+DpZ58Wc2ixZf18Y4t2DjaieXW51iiugdR4hQIjOaFtnkumuOtSZQvn2J
Hm2VJf2+7cAfdqBKd2v94zEnUVXUsJ8BUbI71BbUWxcv7Prq23JtGfGEKQtIrkwk
C/Rwskni7InhUWlNoqSxIOlcbOXQqatsL8dVMH5yMCEJvHs3OuAO5nC6oX7dwlC0
joHYudSXBd5w2gBcy8MCgGThxSwfdXji2V4cCB8g4gU5QRxoPX//HSkqtTpe1f5U
OEI1v9lGfMYSy22v21+ANP2/EaycVh+PnbK7pZVoSQ9JnBgxg/4fSyhv8qqwS1t1
xCKQJHiK1IqJ81dppIqV05aO1p6tLTzAmSWQDmpYN43H7j3jsp7W3+S5lHAGNZh4
gzQ4E94qzoh/cKFcfogL4n3Re1DdOQH+/TqJm/eg+CM9onb6RcJwnSd3/HCPK+Yg
27RXEbeZZPdjlBMBZHKspP0LTalr5dKS9IKqffewOL1J49tenfk1mOgTVEvcLKcQ
jo0Vs8YxajwxKT+cfou1tNAhU5nUmBJ4VkU/fBE5D42vQCwYZmEu367KinUdEctU
wU/V9+foLNZUlEhNDXa/9iMAJ11FuG/0c7heutW2g4MyZPkoFg3HxYISrj9tgch+
5GbM4MHizpigoyCyA3iCcprOgyYYJXMM9Q3uetQWB6QINv1a5unIbe4g/Dy6tRVl
x9j2YvnOaSGO9mBWuXDOCMlHA9D7HNk9jN1KFIKkNBdeD5Z8kfdxxtaay+SzY1iJ
XxFa1O1pZMlDvXLwQwGHmuqY2w+Pur8etT8FRs7y9dIvhiJqIRavpAYa2aH+gHcp
u/oQJrgDO1DYrZeFIS+LyVNdv7QFyTcmt+x/xmm/xYLsddtY2V2Y/DgbYVs6DYXf
TWzLuxGWmg5HmGzg8fq9yRroiZJRr+Sg+i7SlkFayEpMDOuUfnQFf7nkYBga3yUw
huutJDAT/JGNLH/d1uAY/EWfJWwZ68k4yOH8mGbClIwY7TJFafNgWH+mmteCKTad
6j2baxsXfyxg7s3SMg5VN2phBm3I2/A/Qx6EcH82dXYlI6WpXDp/PlHsOpSpYyN7
hdNJ8zdQl61UVhnvq98uV0Rsh3ukytH5Okhw+QU6GFi2AOJ80MHFHLn2s7u9v0vH
CtEBMF7PQBIOFCKM24cpL+x081VBajYP/2Bin0GR887gEtJpMWqvpGsq4F4AKpEr
NrKJjypQGY1XYSQjoM2Kdk+tpiZsZzkdBFXyFBErE+0x/pXDPO2vo6u+56qunBvc
o/uDWlITlkWWgi6XSOX+fY0YYGO9LtGy8PtKxQimNAlqmFfPQeKiGA5hov67c//w
RyofjsvMpWcC58ere7dcEkSKB4+/US8gNlN/hWKSQ5He5eqXiT68kyD8LyctaD1d
AHL7qPwU9cRabL4rHd98m+7s5cHKixlDbxVZmGda/bmjTGrtDn9Fyk18rCP5h9g8
FtHb33bcHy/R/MenLj2BbIACS3aL7ZjKRSrM89DFLonrZ/mu8Bo4RJ9ZlfRTUjos
gAK9nVURHIKn8z591u10LoNmZU7yF3cvm/xu5hX7PGkzqvc5ONUQl5iM4FSHkcrV
BO+R/RQcEvo37L8KRH3k6wRS7QtjsPQgld2KS8s2KBSzglCYmrgustlUQgMpdsOc
6WoXcJBQVdBT6124KXVIZr62fPGGx2GqWYEiI92wm8PaoXM1Rz1dYgAE6b8ky0Bx
8AAfgiZBnxJjffioz4bKc6HUGSpp+/O3tBbo+0ptOJ0gYjxqOnuDVEK3D0uEmVJG
qQNwwgEb6lJrdK+zGn+HN0vlbIpGSJ8PSeYE7oEJJnOuRFvNEju3FHS2aMglfrrp
fugfDWoNc9qJ9Gyl3pFGcoHjDauy7Bq3CngE9Txn/kj7LEkcvP1PWwnk0OHqZ2Zo
7SfMCe1ng37EWNRwOO5wHuFGPiWEaVqrbPMluuibl8KZ3utAs5661Vi3HY8NE2WX
evs/NBgPHD6z+5H6ZgiHKspdjxSoewRN/T4LbdW347M5mAA39gusLz9uamf7rS+T
6ZR+yxLKt99b9EybQsi6AgrfENaHgNH6Hq8rdq9TdQXXwFHew4C2WkieN9f9gPL2
At+RFQZQ7x5q/bxdtpy0xnFhbV1+cqofUdrM+6efMh4lLrtTZMjqWnQjVDrRuoCa
ve4JDsqwRau63ptMfJGbFynSfpfJcpWcRsMVMf7p/UOXDqiity6FC9Y9QfB5jeGK
OQlX/pCu7zyn548pmaaHe44nbKbrCND7BlOG9NG1mySM/mNmkfQvipAO9RHmaPJY
oVhxJcdA4IHPP8khG1O18Dpbw+TLZBWfmMFascrVyUB5PTDjBSw7hDm7hoaadNca
uNk4T8jU9U9uE27qhTBc4ZyAR4vUIBs0KocZJEmKLgzS2PezKXvc+UHe1TXey/DD
dsrWrOpasK2dRyHMcLnsfEH8fmaKmOpAGDcwS7b8P/0aW4Ne60bJPM3AVFj4zzrw
aNBugH4eQioYwyuI8U0jYvVh4YrgZBH/C/f67GE+vN6jfCDvzaEIYUZdxlL8e2+A
IJWD18x+fh7IkSIcI+AedAWOkOa6tyBl4/C6eEM712b8K6SoEAs2CcX/Azt7I7BS
ji+x0e5azBfKwop7eR8oKyuSiSBgDzXbvoFiSx3KhUKhKDNNzBbSFMdPuGxhDcWK
LIKZpxBu37SRDkKjC9OB/sCXJu8Em68j0kKcNXUEjYW35oBc42pZncPenPRu1pls
O5Om8Vngivt/XGY+i/9zLPjqvpsk1JdCeRf9BMHrl1vwwM0IK2E0iO7kBkxrRBTb
rYHq2njyaWqWj5khdL0pqgYEbyyhLOVdOJfbdMBTBhhbI0WCkQZzuyZD6HW8nJfM
Yw6G9GqC9+5Qbs2CIsqyTwn5Yodrf3zW9Qce2FxK6F0Ke+XJLPBSw7k74RS2CebM
MHQOkY93Y5emLLxgzC0M0rmU+bhefolGqy2ZwvNHQwvIfBUWBtKn2HXOAFMrpMsH
Af6jEWBcStAahgKMQMiH7TR6n8qiTZST6w2N6pSzDtHl2vBlEPEswDv7Yct3bT1j
oFyZuSVRYwRtOt52YKEFLN7bSBHRt7ulpd281ruvk1QP9jVmHsU8Q055GyktrRVi
Bu41u6U76i1JblFaOU4B5m79wDmthgE0d9u0pKJbOfdtcRsDNcNH1kCGdSMyH9ns
NkB4XbyqgLj/n+8YzQwjFhDtn1QX6UtmgtpZ41n4DnA1xut4gt155dctFw2c1lsB
VqOKYKt++jTIE32Ur8bCpKPvplTnMfbSg4N2AkQ9+sO+Kk9TM+zrcnt97xjXlf8X
ae+1zSArtgvDM0gDauI58YuLdvVmm/POEygrvVsmVgks7ccFDr7fD63fpI+fksNN
pC7kxI74eB4ueIqpk+RKhsb0IulvpDjY9RVWLvz4/Zhelg2JJEBXytFghkkeh4uw
J2l7yaPUuOJ06apT2SeRYdZtoBFN6jfvbBF7Db3MpaZ6ABsEx2EdG8V4VYWLdEsk
m6Fg1Y1S3H7oAqXdWJxMhRDttfLxVtT/hlArpaMIv/6HtG/jka142vC3DWcO0g9+
YHes/vLXr5R0JKjhYzQ6LZh+OKv3Ab2uOw0XbIEIG66BcjY8/rMCZ1QEOVA930P7
5+Cw5DI50biBxTYn8YGRGoPtLi6kOyhrE0rqvD86cdOzkZhwKI2XkbMxR3swwDhT
kYzbxeukX98TiA8H1u9E5BB6xTZoIFV4lmql7RrVa82iM1f+EfYXnp+mCF7YXHOg
98yAP4IrIuTACI2a/H3DiU0dY+Tjesxdy9DpX/B0r2EJpYiqKgz8zFfc0shIYgRb
IBy3Mn7u33YVs5/ovnzhtHwUxwNLVoxnyrakvn02D/xep1ZttzCimm+jsFK12JBz
O32QV1D74O6OQh//igzeiwjrU7ywSf/i/Ua6HO0gmXn9l5b+k51lysk8drNlXRP3
r0sgW6EHMQEpgl+cvWQ0RwgvRCWe8qXtTuXlhOifcfqftzNVrDo1EZzXDq/IclKt
78x/QcKOFRKlw7lz47etisR4T4f3/dKUPI3awicYRZx5f6lSuO0p0049572wYEyP
PX7f/3Wu0xFmlNvCXT3hooT7AxD7ok1XNzcaBbW20KUSLfMX3D6kbEsVhWNbTuwZ
7oUtYScH3iL0IxTHaNO2/cSNuAVFKc+0vdMyKfW1Z4raAJ4bfGSy0jxbnoWHL1Bs
CqFHj0VE6bmR4uMLYD8m4RDEkc3/ENlc3c/KTmX6YyZdJdNEqiJN5/1UeN+dD1hd
oOLEoLbBOfHRMUUEBR997qPBW8lzf9AeXFsjh8g/IT5O8uAZr8ZuajgXIz39tgax
9v+/fQZKD8krmuGFEJWBGvLjxDChdjrEf5MLfM4qOs+LShdBvy0Q3q029Nxig7e1
BMO+0befYNzy/Cg8RKdwVccLxO2zP2XI6UYpqK4HnqRfx+wMnMF54zuWDQsaCBPw
N/P8tAiG7pixsjcUK9zLbcoYh1p2AHOkoM41NvadnxB1dh8WisgFhHzqbPRc2+95
VZnQwvoW+WWeuZIlYH/fQDVStKgkCDkpUjKyrojK35RshTQtalpUXJIts1Q6qIRA
dg/sC8DPpIASNS16u/2kq/aBxt9YXt5xaC7QILBN4BJY8edIe7T3FP3HydF1ttBl
VYoFtjmAWJEH/wM9tqKDT4jucw3y38o5ukcCdWwyqH1hOlJogBO5agaFuR9RIEms
UGBu+cBjuYR2gQRsoikYdpqwM4VFBTtwyyjSGxYYPv+jf09Yg4RsZZ9hLX7RShPj
k3qjOGalefQ+xsiYxHZwg/FSAh6dfJuUXiK1PZDNlcxgY9MSiRO4RIje4j63EmAJ
L5/uopo8gKdFeovwCgr60P442r80KSqw8hGdPmLZ8A4Uw92Ci648Dbm30mY3oQ+0
lbcPcuvKHU5qter4bixqjBUb0UWB76PPFWPnzd5bR2fOxjHJHDNKr2b4yUrVslLl
6Xm87M9/mQ9eE/vwvfLBsORY58L4lpnunVjrmSzYua2rhJIaHUmQKWEZ2WkQfeZc
CJNbPo5EDbkOwBbIGPoeSiKBr8mxfRkLlWiD85+vA1/qlxf/Wlh0KBkq39Yv0IiQ
Xotq8KGHHNECJqRbogLdp6hrWn5x8ZKc9mxMOpJCOXqrFZaNfRpVbknb0dqayDiq
CucgVNpQbR2at7l+Yh+6nuuisy8zQ+0bJFMkGE9vggoFLGWPwpywBPSgsgLZTxqS
M3EmiU1RnM6fSjkNTdrI3HJw57OjwPgLmcVpnp0ZEwG00yA9zlawHW+ltudRReV5
2V7V+WxiKuPqbM+RcoI+qcnEW6sn07YPA5N1j8esZ9WpTEXx4LKqyl7adtPf6/60
oy3icpaF27lyLKLp9pqXyWH6G6SksFDlmGHesdALV8drrBh6Soj/6htRrtH3t18P
8GnakuF+6SL0vjZRd5GYL56PCfGiPSYMH0OFUTNOIYp20jqDaYc5quNcSK5Oq8ji
4Smdy1v6gyKS8i6M/598Tqp/cnuRm5ABj+OBLwKnI74qMq+hjj1/OhlPCJlOpIJP
B8KZQyW2AT1UfHwvVhItbGTgXlOUlIekLhw8c8NLbnJrxPjt5DJhYv93r8KQLJFq
1r65sNo8YpIC8DYlaDsIW+pywRXGz7tTzo6dFwVoU01rIN1UT6cRK7heSftIVRe5
D041qh/iclAZUz4vRyn67/fMSHcPDQ/WM3Y91zSn+m8EDQnw2I5Jnzm33n0INxtM
AYLi+Vz9j47zT3pX6KOW7ZrleIi49LYSPpgGNmVfGDVUMaaDDHR6DrVvnvsKdro8
ZtEZEvOz0RZuoxDVAT/fIlS+DjcunEuOCPqqCxSVb/ocrPUPTDb/e0jyeEeEX5M6
2AT9Ryf5TyjatZqNVUTQQMSUgHYOFwdg6Sf74tZLCT9XzxIAAmMOEsxGQvBX65hR
uK8+XePw0KJnokLYw3KxCLTKIphOz8u+xt9zotO3jXx5dUwo/Mlys7dQB0psiizn
1bGgsp0QbM4dkVDu5awWYsHgCgWSduY0o/IMS+g13xRC1EeAvB+2kGdEV9pw/E1b
mDGY8hZlRvZQpdm8cublsfJxC9MaOJcikzqgrqoX/addWv4+Ft9BFyf+TdfSwQ75
qrUjGTQmmLmfSkHS+5Wd3oTNoeWnGWjIHmL8E0JujZ0O/3uolq/YJ18dXbPdAjG2
fAY8P/T+vv+jj6Q0ofR2cNATmyiDSrV+ol4u9v7DTCFLCfdmzo5JaDmB4gBZjMjW
tJ7/uk8kblDozi+24IgHBA1IRUAFrYIoZBaC6c/ZZnPe5GBfrrPDDPDOd/VBy6xw
yQVDn86SvI1j7AqcV0+uSjxUbr3M+FKPwh5iKPAxY+1IRbf2QHjvyv09s0f7sWX9
Yz2LJ18UMlztK+Dp9aI+KIjdB+kUJInA2ZHWCExodgUaDOLFKS+LnUiwwyFMG98I
A8DrWi7HNhXhATwo8QZCgLuCUYR/qxzC1OZ/Gtf8Xuy8+yEEJ53WZ2nHJUKD/juU
66NiG8R7B/4fjr7N8s5zq48qRFbc+KG6U7mPTLpOBqhya8NfDMNWsZ3OkJhvkfJY
wKX8TEsJH/TrDtO7g4wETw/W0DWpReAF0+BWsefjMYZEH1EXv/EHbinktTcuqmbQ
1ScrZqx2/YfH1NIk3J36fAHuXiYSBSmfxFMdF8C1doMAvLdYzwbnnljsaCq2N9Jc
dRmVjLyKjoOSc/Qnu6Cs84h8YpdXqLfJ7geTbqonkHnFg9IZ05VYJoud6bZ0S3er
pd1PH5O9dIbglYUy3l3JG9TIUe81lKuPeYf+ZeFwGRHXVEozl225irU67SsVa95N
E/BRxxWggXrd/pz57JFX6VcGZoyDuG3/uYLzH9E5oRVvAJnnWTqYY1O+YCywqsFd
FtXEjzCQa6Y6WLxaG4nrCSSMvfH2lKAMOwcLGNh+2osl4uiDcoZhJ+g70zEU6bBQ
G8XdkSIg+zGuGTkqjeLb5v4BHU5JcXrKVP5eeMg1cxl7p44cub/6pLXL9R5dSd0F
7bNw9sRE/9taxKxnXB5X1WOmRuCY1RacwRQXyubZfQ2afWBCERutdE0xIlXcbG7q
57p8AMC742MAhLQp7upjX/TE8H3WhRlFy0T6XMkZ9NtRgwUROefAQS+CG5P0zzGP
L1F7cv6p7rFYJn+2mCJQ/CX2UShnYC3CdPKX7SMPBZM3qMa1UPDLpMOOvvtFIa04
EfTGqeptiOhUnZjhElQQfjizlPOJytOBiJiUToKj3ZYKb48bim3HVdrcHf2+Jejf
ChiUBfVC7gS6pTIPLHNG5RK8GhVi21Pcps8KLay8M+gtfg0EB/EnHQsmdIksL3iq
QK6IrxxStqjqxtkC+12h52HluuKrFtNgDbD74288g4uiOuo8S2jffidouAEid4nR
fbdyzB96Zp6okAPtPJrJou931qFryMjZOmkUepmNoP0y5Wd+E4nqRqCZRpCKsW25
ocMGLZ8T7QAsQcdYxWyVkWk5XbHs2Tr2/Zwi4FgIJX/ncBtxM1Kdc4yBv+Rn23ec
pR2H4dxlckg0lxXblW6E4wvOYaMHz21XxCwjbL7pPstN2/6a0Ng7frJ1g9pK9rEg
JiFE51w4gn509y0plz7myix3AVyPFnuKBTFmSKZhx6X85CeMd47KfoPYIxdv3M/U
7Z4auesfYt8v3lAe5gYZMDcRokk8pKincCyXsCSqkHw+QH6gZ3BTro/ev3QguSIZ
uuZoFfrdLvYpdZYDPBZohu50D65skI6hsOVMvr9TPhRMMLjWxJ0Qv7bdisM9ZdR+
SWJOcZKgcIeySgUWbYqTjMP9TLvVYD84EoKXrAtxPSTjdOiQJSDx03YjK3dNQk54
6l46gygs0ZQCsQQZQrKd/RrGAy9/lyVwfxzet5Q8bCmqAIlTxWwLZC5dVQj4yz0c
jB3H42V+nn28co51RPOFhVCrjUBfVQu7NjlUps9XEuuuZ16KjuFLvCDcSCZ4NV6y
SXazZpd7jifr4GySKU5A+uUCBYmXClr6lv4nFJsZcggsymRZtwvmdewFl1S0sixF
Nz0mBnVzUkF+svZv9qRN4B0QFGGUqrB0UcY/8VdM1pxF64fZPJiLCqPSJnYzO9sv
OO9nvNLWyjaAJBOmFQNa3aoJGm4oQiYGKaR6N9CtnfStqd8NiIiM7sTjYOD6IpdS
lXvSyMpSB4uarOckyR0v3I8z7MN/+uFx17ZzeNCfe3n3x3fsHyERKA60VfwYgml6
mrKsEj7bB9ntAs108hbOj0ohBn9QzTmfKjaJvwvj78yOB4piMj2mfKF1K0CBj0ph
cypzZ8gNxj6vwpG3/wdFebUdw0CeBLCsGvUvuFrzk3/H+l/UH7rsEqx/r51tp5DT
2HsfvK/0ZjkCc/EI+BXuht2GgmtuGQKUB8HERU7vkRjy+DVd80XjKJlgqlWA2dm8
lkHvRYGkg6OZj7QftLQKUazrLHjaw1Y5Qev/hgrEX+MPlp+QmuUnVN5T77o6lcyD
unoUIAVSOaV03HC7pBNWRO7HRiSrs5xFAUiilBI1afDyGr3vp47gGgWUFCEBP7bF
R3gqY0kZFCJB49EbdHnQ8obI5CtXt3ZJe3WBP84LuD4Z5meaSpQkGHcpkfmL5jV4
F5K1G6ErUOG/icOA10j8d7I1WaImPMoZYLdrv1Jk2Qy9HFJEeOm3oHUs6oKIIlZr
ZZJK/cph4TM5VfVifv5ewC3mH8zZRM6iTODikur8PJFC8ZgvGx8pb8M2cE8EVLVm
QeC753tgO+prF/FMlJPtTp1Z+qq1LqERsjNI0DennUmb0ONzFtasxSE8LQil6Xnq
7CsJd8Lz2pSCeEbxKfln6+zhd7BLmp2tIlOQQmfMNok80nNT2lT/h3zhAJTg1iw5
50iRRfuXGjzkc3++JFH2WKi67K4W1ybvlNwMlz//Fv4E6x9i+7q8GkA36LVt4uqu
bJtVk5GzXQua9NxFK2lqZv/i4xLfNuFS50zTatDh7rdlRm8e67rUHinDuFudxB2A
xwnIFr7fHzoFu4KSgNfT7mnc84+WoETqjC+gOVcfluqrPvO/ycmc+vmKYtZFEzB9
8cThFWvRfK+yQ6nPmoMn5QIJn4nESAKDnjOxi2SGWEcHzS2aCuHOYH9ZdX9I5jwH
ZwEWFAKIDE1yejn3QBfGbzsTclfx4lngUNFxWyS1BPQLoJX6P/VJpY4+vA09mTfp
Ud/b4uVHEJ/fBYSsdlDLv3Ky3i6GDB8RnPCIaZgZZ6lo1LImnh7xSmmvgkyccPLe
jE9i8D4ayCw6qC/6AkPVM2SzVFBH1mkWB7erw3nZqt/wn6SUpWCr9N6mrtCGYnVW
brWkm/zLd36TPc3YLygk9Da/1Zt7OdEBcE/9XHplGe/slkMDdkTRYNsWGPIKaRKA
FKCOmqu49TGxjVHuDN+XVULM/GwJ9vP2auvLKMsEYz8zp60/DCKrx7RNWeHba4SK
J/AB6CPSQEy+8tK6bNvjTc8xERspGHMUKH+k1AY5S/6izl5fhi0b1cozDitUkzDG
8okNstw1ncz5vNlah3/7j4R48StihmG9OIwtRPwby3VzuiDaBuhHyRW51Jtpzhik
bL3KuJi8blFFKyoPxxPGjQSISuEv6ChXNh/YiV1gybbpO3P61EjReAHtRWCErlSX
DS/fBB7xyLnKCXoOdAsOkFxvJZ9uUtNDab/Rcd5HtPUDu984dKhQo12+15ELUjHI
02j+7c4qAm7gHO46v5IENyta2zXPYV9CNvic7D1uG1xyH8zsRoW3CMet+GnpSsjq
n1a/deZpACo8PIr4qF/jcpR2ez+W0eQxq7ftVb6fwJBB+HV4tLnc6rOl28HZIkv0
tflELLEzjHJG8mbsek7EhtWu4LuZAtO7esh9OQEq9f2cPAbei4utpGmuX9Zv873s
CkMG733ZHRCdYO4BFDdw48/6922L339BUP751bD5e+ttt+cHSCLPSB3MNDtHDiS+
Ahif1cNV1A57tZ4lykAJ89aZYMPS7kVjk37muHkyPlARpraWj7xmYY4aMAQkWEyh
e/+ysIZcOiD526MhVd3jdGyIdZLX1A+CDzrItbU3T4BV9u4KmqPnEJ4LPbtwGtI3
0v03UQiUK13mGAJQn9H9cmGr3et+n3TyfFFyoT8qx83/NlNLwZGqLGwtnxYVEDKh
s78RxXFkh2uHzJi3r91oUCqE2UqhQZBcpsovi8fTwJwoLHl2TB8iO+G4iwm0h9ai
N8+edDumXtYkOWy6tTve6tJYU8fRzvZ9f7oHbdfeL2ZqJaiDUqlvj/8/mH7xmUhO
Viho4YS8aNT33mSUkoyEv4Rnqz4JURhI35HnHHPdm6QPrgBKC5tgxL3ejCsKKZvF
P0UuUYVW5V3dRugZ/hVWSfVIxpLvhRL9dw9xHzAg252o528ISB6sZEz/TEsmoOZZ
MmD7Snmqox5Zb5bY3xTVJizNLmrN6u8Qcbh36bX7PHn45Oci7n2tKAy4zHieCfDW
Jmn5BDHssYN+1ipulPZ9x68OSbp+TW3QEONhkJwZ8gdAVUATT0r/6Wbczy9Fl8KL
SQII8PclQwQNyqBOtxbfHq3d0+M3SZxb4KXQH0WA4RnvcJpa6F0+zggYmH2izemf
iSmCDzXqcdCj5F6aJfRaZcDW2Pp/HkmcdU8rDH9mamk6By0F/+rdKcP4g7YNU32R
nef5BmA2yWj3qc6ND9ZxiTJ49QOB1nKfFfFJ3fgaVvjoCsHn4Fd1a5bSOn9+NMhK
HuxQZkVi35e3KDMWTeES1Xc2eSgoE7vgVElIhLiKV36rQzYNEgClzRuyk2Ibl9mP
crOTpHUVsW1r2NZhUMMbMSgjNpro94DKPWokKHt8YdNcmZ/mtCexDPnILUpCm2+y
SwCDCVlHkyYcWJA1OTs5AeinLz33LPWloSP0hhcSAw4VXRy2BuxdHZjGH7wududV
ws2s5HwpVex42YeK5wbE+1j6bVVRvcMYgHqR8KIQWMs/U28//+/KW90MZCF2srjo
CwatIsVTw8NmH6cD1a0OSi6d66DJ8LTu2nb/nrOraQri0kYX+loQjfNK+oLM04Fp
KfxTCV/H5jG9rtNH/+DVYSvLpoSb6gTX6YJbUVPn354QLvzmmW5I99qSXXjWEO8Z
QEQIKeMnh1JSYPCVxdKiCzUMPdRNcHGx+lue6J2SKzLyNanUVU/+0PuKS20toLyk
5/oMKDh572iO1zdsYfzQzHdm8nvCC9sEsJBthod2Z0XI9+A0K6xPaXAFgwTG30WZ
BhT6ZViOsZGYf0CDpQwEJu00Qyz7PSel+JupnctKaZRGv45wmywQRN7hIfYnzmIJ
p3IUVJducJbvwY/8wfQO/oHzwtK88XQ4u7zHGSVQCuQ+U+nsT3UWY+gD4Ekr1YUS
EQerBrICnzjFPIyo9IQeNO1EKznAYgHx5/K4QLZnO6kUmJ605Q9mzfNP+mhMSmZL
l63GpShN6yIF73Ryf7rujWRScsm98hLptUyikvYyPUHTChtPJGFsFDkwJUdF1eFg
6gSujBSRMgxCiHd6dMkD6aUNuRxK7Qz8SmrKfUKKpoVSkblvwAXsCPL5lT5S/goM
OJP1eqCPe5SwR+18m8nEekPjfbHiu2yp4nYXYAA+pubHUnJEVPyWHCwmnL+K0Ulp
LU0etLAF0dwfqS7wI7CyTZfhUZ/yuxuhjEOPdF7DCiskh2kPXlvmgso2rfuCsG+M
hvrrGpvotK0sou3E0fjohsZQtLwZ2qQjnuNwzBSd7nGpeGjYjXE37iW11dLYgwTk
kQkuJu6nLCyXK+RWeWIpPs7bkjagQ5qAYZ+2UHEwRRGCXF8/2lis7mkNg5c6kySb
jekS9mtqSQhZ8tmAzXTtbVeTNA5xfyxCWwvb1cBh00sK7jtWb8P71+9HIOMgs0HR
jRDLsDAHYoy1HM2RRmqJWfncsE7DWagTY3NbkVkO8uknKT4Hcjf6FZEtbdWVh+EL
w19ftrnWzexmKI6TQGk42y6VcmXBrVVXvPM5I1NVUMF++qgI+wCA7QrnEMCabyVq
2QR5ABl8tUZYgE+4yzKe4w0YVd21TxnUeF6AMmJiMjj45/J419L9ZlWcENbmcfX0
Y+BkWRQ0aCBjgCut2x0ZvdjXSJNs86z6O81LSfBCD/vN+Nb0TLWh6pThuI+RKlwO
`protect END_PROTECTED
