`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRCCUCZFkBCU6sGNxuK9sZS+dOTG8GRMs/p0jdylmhF04rNJ1/y4pDtpx66J/J4G
4fXHlNK2rnf0yD79KSE/VFGSM5/7YmRoiEWWAuj7B8GKUM5nsmgW2HusVdxjm5Yv
o30hjORZhmA4AGcfgxFR4NZm+qwq3Qkm2aZqOGnGSXRBsAL5/eGDcDAqLK4YT40M
1dY38gtnySA59lnJl2IlvSTQUomHz/3U+wIlEXd1PFEk7tNS6IZ/a3PraHWjLRsd
At5CXaXjKhv7TJzdcVp3HHUvibi4pv+E+djO/UW4KnjK5TkT8t7duZPw9f8bs8Tg
3B/+7qJaS6ERUHKhQ1eZJ4HULmyqV8PHHk1iln2Mm4pR+/ZmUVuDoLgjnjZPndnz
nIaCi+cHCVtGHVlm/eF6AYw54f/zryUAQRBvYKoPXMUjPFLWcrUk2JBOM02JdHGW
NtWVhpoKRQA8DRdPniihlJ0+d/gehuGlJkm/DNvbF1VzqI5LFqhQRfjE4aVnjQd1
ceo1BwQYnGdE7eQpj+AmZVO2usXrOo4/qSeiyGFi8FzELTg4VKruOHOSMDHvgHW/
JREBRJNVr1k2sS8PVYoin/c6FK0YI+eHCtYlTAgTKJVk7qQfqgZ+flzcLPN/3wO8
5uX1smX9CA9veC5pT3TZSd/oDO/M4xCioXssvlOkuoY62KHCf4EMiuJOeyScwQfw
px6h5cTn5TxKAZVUhMcpyDG27m8z9Kph0ejaEhGQmmn0Af/5XmbL83O/Tgizj2F3
Kqqn6a9JDwZ2VfkXX2KwKYpvyV1VQdFFmPPV9jQxavwNLT1WoJUPjpmDzkwRhDRM
Q/Px1ly+M75Y1k7ueXyEMg1HvnlCJB+o3V7Rq4W/lenBvbFmlvouKanV1/fB++yM
qbwq7ETPj1JngLZm3K7BQ5wz1OBtbwcxJch7ovaoit+fOADk0PA7/pt0pNaqR73i
v72VLKQRHBzIF013kN6MDONqBbvOqx3zdF4UjcuSyVHaQHai13qY9KT3b79KriFF
+vE2c4m7KZloK7FI8ZZytNHSN0VHs1ciRkO1Jd9yeBcGnBNMxTeZBNcubJ9bSP+3
4saaNVQe1tlHcrr4LRQfZqcb7gf/ILqD5lWduF3aOxw8b+I1non6O9vXbH5pIOje
6gU6YDU5fFMhjnlUflfh42jih99yr4TGFcEKqSmJ1e7zTLeYuHZTLWOU5+SV99xp
jEZiuvFchz6DNHNcRfl5skYoB+N1zGibM1UUh6w/AYEYn9IvO8sYYtvKlynNHxel
uNQoQCrhAUqwkvOQwNTkNHWtYGY0CsNFbYzTxgNLOHB1ZxUim9IdOZmYZAbpBRod
Ixbbrm2NlccugjvhOg/qJcLxzf37yyJVVmGKmNaP+Sxnl8zx+7q/H1O1jR0X2Dla
2pEGGiyL3TIIU6cg0B4XwwYkMJ6PMKZEw2t466PukObB6PNKVg6VfaxO7UP0D3CW
3+mr8a40TM0oIq847ch921B5u+BeCLX/8KWSHWgL0IRkw2Pyfcp7tSIVMCEt5kje
1YwM80DAQyUR0nxuiePMeBhhseGE00Gzk7gqkN07piOknd+enuqZHmk3pJmxvfUs
a/x81CSEhA6DXNAb7ZXrGIa9kA/ex6vntSU7bj05PaVPoTV6FC6GhTijfClJ4YGt
ak2fEiCMqYgPhFPF0hpMU6MrxSUu9h0u01VMzfmsZHBSdC1qL9ukabWTgx/4ZaGs
HtVFGbZdiOPVPu92TD7FdZmv2XCp6wwYK3ERy1HHGyF7pm9U9VNroiLuMVynAGSS
`protect END_PROTECTED
