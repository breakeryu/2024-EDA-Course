`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RPzbRrIs/4mPjaPmbPnavlZ6Cm0CffW/E9bIUeUpSuRi5/9U6kX5DYI98iAaEFgv
pZxLtFjYzlWCuf4phI6TkDEZhSf7h/96IguFw65zGuUWrhORHr0QPdoSPxgl56CV
C9HiuMKRdvZ/YGHGJGDdw0SyiImYa6gsJEm1S7sIhH8Ixj2jBvVxsPjph9D4jGwi
PF+QNgDlGzbIiio7XIqbkNVl1qP58xN5bW55/foKK18tXkE42tdWx8+/qXHMsAzF
LIX7smTzqt5FZO8+iYqZNqIzC3oR2FOcnQt8qanhkwpRrjjmm0VbaGak0XSoykrg
vT4AteeGuZ+2BXvNhkieWOhLveHV313r0P1zrqltvfbJN5HYcFTinrJ4y1P/3t/h
imxiDK6W9we897s01aYh9sRmSAqfmCvrv1AXfMkMuXxFGHqIW7wlpZvLuSJux7T9
aAOrFily5+SrdithkI2IdML4ZdNtlkTgaliVtJUDWb33+Ipm0q9w1hxyvgdYEJzf
CUzL89KCzvZR0oeZoa4BokAJ+pEglMuM76ZMeBTnAgTTHpa6BiC3w3DCsLMqp5bf
qSpkHlaWOUe9N2w4sVO7/kiHZ9s6NXEv9Fu8s9RXpd+HpBQ7q2Hs9PKODPaMeZsD
UIjc9Gnik97CR3CKn5p+20WYQYHu8JcXi5DXlSaBXIWiwhc9ZUGLyTLUXGepFbNp
Fmh2O4QBE/RlbWwAO88yP2VAhFvgzRaGpGOQHUhdMuiF+u0uAQ3tO5D7W8CPINiT
fr1bNaYjRcauUTsUr3wzDJIqDohCkNR8bEa3ji0Qy5UpjDYQjGnJeJDjfHM0FH5v
fGG9k7M4opDBKAaXh5O1apoLWw9wMTd7MVeWCvPiXhFfgL2FahX6lRQEFdYa6LRx
U3VYOafbwYj6H8oQUtJ53wNGtvOZDVoUZQAIHu9yYsKUkFXOysCVhWlz8pam6IPI
c4D/wd5bWnJXiSW5gjfvRDsPlJ0lccL2vfDmrMJS/ro4GM+iz/C1kRKMkkImYUwY
TTZQsNUbGaJokFG6pbwAcIP2HfOGSOIJ2P6O3KtIIvWTB5G0eBDvT5qjElYv3ZSl
fQ06dv7aMNEAHnM8UaF7Iv/AoRiBno7DviFTpu2S3/o1BCJcT6R1UMv6swvDco3X
hey5jlFLcwiurR+an0t5se2B46KoQYwcqnBbjbp3MnNcXjT+k1c4eFz2kK97sUm8
fFnY+76YWidQ9gLbsxhguO/R2dyD3ajQgWdT0AClKVA0LqEzvOpdKIziqftVroJU
`protect END_PROTECTED
