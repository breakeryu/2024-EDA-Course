`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JFnnK2zLtJpbLDXIzAj6q7auEiSa8KL8pltdNYr5tWbFTJ+VwqbpJTS6678SL/4G
aseio53Kn4s/OJyhwZNjckv7PCEH1LOi2vT589BgIBBYgZ5A9vGniC8POPWfmtam
djGVY3xuOK/FoeFyjUFBk/QWlcav0L23GNeKX/GL2MhZBek64LCSYwbTNoUM1TpB
hA/CRkHdgGK613ZtVzKydF2MHyadmzufbu1SJIG7Ll0r8efw5Kej0aDCiwvK+kCX
gffevV7E6DyRqiit9m9d5nsa5DR/SmauFw7Wjcrx1piQTu0hYCJ/1H65jUQ7EbPL
xV9lDjhjedXy8LSLjnBu7qRa6AcfmuDckVB/Bk/L0z8VKP1ivuBbBDuAKarZwIzx
w0W5Al/XcgADqs0IqwwHp55t9y2PoutPtbSA8U+fNM3LOVMcx/ZcO02SBTzKv3C0
7P6NPGKhxKPbVPJsUMa+V5g9wZReryio0nXd1ZT6wJdHmwSImNsDGc6JYWq5Uxhg
fEOUj9OiDhAZgoK3uEPV56kjsPIGVrND/oMqmHrC42/soXEM2r9joHhzWw72qpW4
GD/ZL8WGWKRMrB+KbjmYcG0gQ71KH4kmynMoJfpvgm16b+nYxCMkPnAHvYGyguj9
oU1ZH7uGbqpT5qMf6IGV1o0Us4Xh7Hr2Jh3At8Kr9VekHp5z4l3wt/JWwgfPCwIC
6MJM8VusQy5VoSzBdalrW4Il+MZXYlrdDKveTMCShyDJkgfd+IRTrF5/UwzNY8nf
mi+xvnbb/3qQQl06XVHEzwRcnHZHKbNuD69DBuhPvqRiUWFLdfW04H4M9JFOlA46
v3lgx+P3uVb4JOeHrMWO8Ko+/PxN7OsHqCuKbv53LFt2UACO2i5qG8zgmSiwWnBr
2C7nQ8sBMIuiBEZ0pWIHfelRPPVjzLOEJWYOgXokWECKAuHNdQRnPiIqTxkRG5Av
TjfsdyhxBT8UDOv+2DSpNkzoKEbvMFS+KEFSdc2HfILd+2rmgH/zX7sGUteL+iL3
oFKakwR/V7vfJnon4Bgmwv8KtmsG0JvkCtg4vPtV8IiEoXePP1NFQXnid/OFgkcJ
TMyH9KpQEH0CRvo1f1mAPU92OIW4CAA9W8TwY+qeLuA1iPYmaL+VIoI6oToYVB9a
c8y0BmfKaR0D1RyHKItC0GWnLFsN+Tx2U9La70iFubNmSb7cMZaWvuXmx/suyyhd
Nkq1sfWJtTyfF8a04APQlouajZJDexJq7hLlL7/mX3IsCk7o+VCfwY38T6ZkxCeS
Ru8IiGL85SSB/5WfWS1VBn4DUqpRwCzM2YQa+LO9haf1NU//+PDsjw5ZWwED2d0q
CcIwCckh7vyUZDQfforkJJ5Ji8zPEohmmoF7CBPOKkHlvz6lGDv33PJYq2KI9V5B
EfPbt2FoFk5/QqZOXjpt/J0kn5icRWwKfMdyPNjHyUjJT2x96k3SO1BmDKqd48ti
vBBcd8Qj+qaRbH5qnTrej5qLD3XP94UehR1ubtHtzRc=
`protect END_PROTECTED
