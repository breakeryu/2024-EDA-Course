`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wntUyW4zSlGSK4/xyYohYjH3Omccze9fVqIa12OrLswEI62jskaTLVpulzp5sODR
iv5coUCGqoaDy7sDZl8tNsFdhcw3UIQJCQaRDsenCQtjTs8dzFJe03UaokMwfcW5
bbLi0xMoR/6OkexmAr2XHOFKEnDav0i9YmqrzmimN/+zHySVhPozowt98duCzMur
awGWC2luNvlTJ4LVRXEzRBn2My4Bpr+yJrotsEcwg3hD4evJFi+Pwtvwp/+O2dy8
ek2mM7yjfxuqSMgVMXxDRTHTKMuMYD+rsmhxgN4Jj7pNicxhoX49TcTRN/esGBie
9LEqIWGUIDSrt+bzvdU18UAG8BOwedy1kbBPCH+Y5y79jMrP5J4cs/t8FRRyWAIF
lNarv22mT/bTipT2yIdFNexPC5O99Fb1yOPCURcS0RuxPZHA1hQlxFACmuGKup4s
IGqux/Vi3x63MZ2bZICRs9DLpyKpBOHu5/JyOe+4xuwYU51rJqe5faW47ZdOWGJd
mqSNypjh1ys2Ul/a6kUgQkSp05sXSvXcpb3ChpUeBe8ISsiThCpY6y0O4TEJECtg
Z03dnJhHeU4xvESZPKKySkEjlWwQ4MYTwYvnWpn5SCxgzEqBrmhHfJwgCsYxs7zp
CR6DX9v+MhBCwWsoKf5fNjHcL6aMLXKFI4WK3NbrRcyUWakPUbKYPjnxY+ZfhtQE
gnaXuwvmks5Mb1Tj7pqfZRgk9h93v2vbxDOMMUAn8n9xMVB/YKmSES04Tifn6mVL
D5ERIKoXYDvnXVHsvfCu8KqvbRMzC6CwdszoR4JwT7v2ZL9M09UPoLkFEzWwzdeQ
pvj8u7Pi++9NkTmX8vwLQa7xsKXAxsnDVcSDX81oyZjZmNRodwem4vqYDf9k4JPN
4rO4MYuu3vGRiyVLmlj7f0RQopZHZaY8Z8+otgpdc6IuhtQtioz12qQugr+a+dK2
lnynv22j2cH5lKdMbIM+qpFHFHBLYTpidPn+WZba0S3Z5+nX+lhblMtLzxn0l09q
Me1xYMcdmfsaYf5eTOkiNFN0NuGqLYIGGjTVRJkJTwrJJPpVE3JW5NnN/pWz8N5L
UtxBFvj9DLZf0eh78VbOieko6hdjv2uFWKGf1KuhLxtJjaT8gPcR1wxpWtKoGfwC
6mPaHmAVdYVRpmXVpg34twY0Y0AzaggEMbO8c7Jv/Tmi1q5i3YSmEmLkwcrkNzuf
GXPwqK65vC0700perwKIn2ZCE5vKVco/Uuwk+8MBg7i1P1PODw+qlXv3RmPrlyHi
r1yiyd4aH6T8ed3paXGTxB/P5XSyYrX4WmgMyPDeo7azt4DBC3diGULJhCCiHB1G
d/u6eqArxbhtHTgZ8lSdt0yBlMO92K2OsGOYVG0uRLS8aOyfqD9846jRh0urySO7
Fz8JQHYDoWw74uI/Ay7Td79NSPg6UkfbgIdR27nn+NZmrrzKfL9HEt4UV+q83KyG
ODdhn5LXMs92fuz4fTyzPt1ug43S7Sr/aGahX9A2AMWQfWMNFDMo7Qmg7FMOgw0x
SF5OQYihsagQv42pdTqCa5ZgkF9yOOz8rh6SQTTkqowlLEjOUQEgVwjCwUOTKr7n
1ReuYC3wYbYGyW9NMHRoN8nzLzGP2MkXYYKhJS6JrRfiwYfxSeKV2zDden1rZ8oN
PS1cZk4oeQLGqBdrBndyzwOdIlKUinrATZY/hDOdvcjShwoaElNVwJCoVeY73r0y
zcrt6gxkxrIuw2ukywbrEznQ2jq1Bu4y9tRLyZNO/pAb6i9UWDMaSeSBRawDah8T
V2mL7GShiBEqxVnfiGfiEDokAP4Ubde1TAslro5x/K+zYJfUDeRN6A3IUuVvUpXZ
Ph9nee+kL/udwQmupHjFXOpP+ZQTpiuwhUN4IRBxjgrW4PjWS9ROqiJA3O5732vM
xRqeoOpYjvPRHtGPPZfIIg==
`protect END_PROTECTED
