`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XPTJcvi7IzImeROPK0DT9jXc0irC+YKmAZBS5uNmfbYAkxTk/OorpTumL7pOp71g
sxnY0FXH3DzSt/tsCm1CIuszwvJAGg1GU7XGXYhN5GPhgWtcdjCXWjh9V9nXcIzy
Xj3jjvvFGysC1qoxN1CNult2wvgmR1EYugps4M64SpJvXrxUcXgb2DHw6+CwEr6q
8cqSahMFmSALpcjYRGtkBigIdQPBG1B3OH9AwSNWCMPhCSKFsNnHNkE7F3ZI9l5N
3MQ1ip+P8K/zsiEr1QYF+dvHFwQ1n6Gi1xpHcChBxwsDrzYU6Q6IBwzdvM1WwKSr
+pQjgR7cw1JPLgymjCYRwmg2SCyYauHRZ8K9pbEd21XlcZowKtMschJK0qWgSWNY
JRlksOLEsDBmtB4XOW+RxsMVIR6dkypljlS1Ey+MQzkr5SIKYcXmfLqWo0jxsb2M
`protect END_PROTECTED
