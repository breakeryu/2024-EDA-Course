`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v7zAbP3dZUsBGMxaRZ9ILNue/SpQKpCxbw84PITITqPZyp4WvHx9ne8t+ekRkpFF
gF2W0Wf7NwPRMQZnHjZYJ8K+DmbmbCoD1rzdlMTaxb+kYAZHbGPtNpUBLFcQFsxd
6kd4oyQKJD/BGg8O+Tgaf0eLp0/kzTEHvm2jc/4yuAHm4Q3suPOc89fxiNq/pdvT
6CEEvF4yCx1NFfnHN5VtpzSV75s45BZ4JXP76YHRO9j/sjczshJJX1G6LfUO6fh0
2aJB16hCxRhruH+oN27pfiKlOTmQgRReWSO/ktHA0ty6EEN/Ng9UqNmt9/5d3aQf
+oglX7u7LmNdPrcc0FmhhOn7sUTD0jWPHedkpFdNhvVH8Egk6Ad7VgLau2TLgi4Q
s2vbs9SH4Q4cKbOWXzcvjrrXPGhLy+Yck5SgBOAC8sSYlEw+iZAdsNq+NVEDcWpf
mZ7I2K5syva68bzgDuMJWWHgC4ET6kE0J1RE4cacOQw2peUn4WCipbME4gzr/jZ2
pK9xxPnadVJ9U7FCzdTCqu3wh1xvmzdICycCfFZ2pjdo3Y4Ld4sBgTKVuoPRRNAb
qEwRPBnli/FidEwuoV0xdQ4QauptNgugZdDbLXFN7io=
`protect END_PROTECTED
