`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcLyLozgOohM2Tfiry5bXlPdsO48Tm4IL2a29y5dtGUYyfhc12AVs4MM3uyJdHvp
bSTam911dfWWjLIi/+IujxmM2TLggR3yA4bnrTz6YmtNtCMMMEesVKtEPXOVo44n
htZNmjDlu0J3M3y/3NLbqFz9jvnpNr6HkFFy79HnWP6BwQrHera+s9TityPtWwvx
aNoMDgWl2PExF0yeiBkomxzjbm+inqzAxBiDqkLfttOhVLRiipHLRPgX8WtXnTnT
qrZJJGEvhf2lPKJsi0u40wsgw9qFl4xvXBvnBWsfb9+s+jPRD6t9IjSRjxBm0vtD
eD131TFzDtlV3N54jVtVHK/F2AlyyHTlRCiJsYrMfWfEg0f1b/uNv75AD+IjqeV8
eHY1j7BmorVrDzUNUCd+RossA2sagmZZn0ZAlJQCFFLi10zEid4DqvV0uid7ED6w
cDNu79jL4mCZ2c5LWGSBVk4kUn6+cVq5nZIOMs/F9mprAEfEmPjqpYgftwvdSgKf
bdZcX6r/ZayARQdac5No0GF+7QdvVrQfbs7EgIgXN7HALL9z0Jybq3nYVre/Hu8V
MNNV1r4FMFLIS0EaffZcFTaWlenJ+/sDP2g+pC0J6ZykjQ3c/uZhWfutRt3lnQYX
o8BMNzTIEeWybWCmU69/p3VAddcKVbFDFM+kxWncMlVzzGmhPGOKBpErEWkSaFYe
7lDNt4+FdjMSZQ0UdScbVD+gTYu6wIbRAlYK5QHd7Fe50qQGMuA2lUpdnckUdzh+
pFdU4YTqniCqVzGwgK8EPWimKt1tdqBRfFfpTSWv4Rc1D5QQ6Gfvrac+tAYw7IfJ
O2MYyN6ek9h9nMquTpapPi05xv5bvZjnVbwZfTJZPhLEVnJPUukr2nTr9MDdRFuT
ynM9awhgRQE2ugqWkOCLQKCl/Q4a5q1fFvzDEsPVbxIlGT5BV1g62v7ZCrfIoFBG
SxVpWmGqBMQv4Grqe7ww7jO7WdFAN187gUcW9gZZNEse0PbIFnU7g9+tc1yVWi/l
ydFSsxlL4MiGEN78zcNnY+qUSWw8g2J65CwEZsbagg0+sR5CcSEh9RmQ+m1g0wWy
iEEf0/xGm8Isoeg16N6koYoUBx+s1hqWCC8uVuYp3diS5gto2tL7/TvCfgna8LJH
Ye2hYDTlufKGKIrLrfzhbHEfgRIdAtczN0kDWmGuTABmJVOT3CvH3FG3CcCfhi8R
C+/Yd3W8Btwk5tMzyE5La84Vp/mXHKHd1KaYSDV1EFHRuCe8uIHLf+C8Dd1BWngJ
d4/nfcqz3nRV993hZwVy/wCpYYwOo7gOvhCRykqRsHvZ6OM7250ByvEH0XTv4Uq+
mKLXG/aUAKON1kUwY06QRRQG/BZWtJ8N/CUilomcoVaR2bwheqlzoW6SO/uSY4VX
ovNTe0kdcNaggd499aYHXdGjL8Hi1qpWgJMmC6MAabq9SlCX8demrghjSXFbrRcH
zRQfNunRLQdNjOkuN0nmlvICIrRDZTRDrKdepHIzK9BOexUCCvY8aTfKL1CTGyXA
jQnECeHfWGzRwoGvyufW6Enj6XMUDIU+JOBe0rRyYCGWJZhApKmYiAqrI1Cvd70k
/XuTLw92SZCEUsIRG3F/tkevqX907ErzdnD5tpoCiyic17BXOu6GsGqKnURv67ZM
bhGrvDX5msQ8r3RTQlPpv4NqDOL2bbB5AtjJQu6zdYlFCumjwocb/2ENDfQIUtyW
1sLZ/e9SLGc8xPKFpNM0YfWr/SwcyKTr39Af/GBmOJnpZToCLFYdqKFH1FFWUfEa
BQjOnxC+i5ZAeijDsIYe4WKKjoLAFHRbww3/9zKgbDfUWoH61KSIUxMKrrdV3TZn
OW8s/GipDNwzJS6iMfXy4yq5O9ZY9tpYDniRUfw/EnpoW0woDm/37o24zb53mX10
7l3qS+S9QyIMLKK2GCyNa2qACDChwIeP5vd69QR61ujYkeFunI8I2lA5o9rPOWeZ
2YazSSSK91ekpe7m+RaEHG3eJwbocKm9UaHLc3YzdacprRcs3ZYqw39jbgZWnxv9
spVYgZiV5gAOSsNjt14c8ZXe+EmBLPPWZQn4wOuE3UiouRnwXyTeke9nkIWO7PeA
ca84OuwrnfToHc8aWHLqB77JjPKPpOstYFR3OZnT6S7gn2D4giy0bRVUDfMCj3t+
5ZfWPCGShGHVMfhbC/RakhjazSuh8mM4mhe0eEokuJ5vIEGFpUuSM9j1Joo8z752
AsVx+p4NRUUJ4fEHVxgVDS3wV0ocwcEW9TMJRY/m6N8BeFKD0Ijl+IB3Ml12baL1
oDTb1TmJ6bSp8+GrpchC3w7GmidfxoN42zJFkmMBUeLnwg1toqpY+z4+BrjdwTQD
`protect END_PROTECTED
