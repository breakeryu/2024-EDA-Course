`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vGYCs6hxYU0RfKUvxkyhuEcJqhLYP+GlNJERIKyAybFIYvxTMn2ta5AFKZQZb/ME
fbdCft/TUzAZ6QmpwTsnJzV93VOAf7SSaDl9WgeSudQCFZihIR4FUmtohN5T6Mck
44ukkWI95WD0rVT2Epifi+8l46LhGsnf2WPneFxnJ4YjjoZOBX4u2BFBFGJvodJ0
/0ewS9iEpBm2zVSulvxutgjeh+0zqNa2MwwIiZSxuflvZnBLJPGx2i2mM62r5RrU
Kex38BZz9B8jU4V/6otwb80nShg1TyCCaJi2u2pRhg6xnv7RKQVM1sfhWnvayMeU
jVPbVk64OfniseubP6Y0MrRJY0Cazxzs1Recvi5TYHBoJCjSxuhMUvvb9lNiuzWJ
sWCsLosubQcYLQSrUybWV9Fq+VGXwu5YMepxd2sjO+DASaCiJZIT8Q/vUwNDQ31z
qyaH7xokfdn9DWvqIL6DeBYSbAm8ADvejpPMMdu4qpUAZFuF4IpwE2R1tklMlVJt
tu6pgeF1v+XrHvGaF6Utm/w0/rveBai9Qh+iAknPXmw09LP2m1e2KHADpf7snlYY
jFOpWndnOpHMTPUCgm8698qwhF/5xmGBfbsBVYUsEHR635DshCyCeJNeTcyxR9G4
B2Qdvu7NhjS+KvWlmTNjakj5zYjEJs8aOd9miiwQte+g91yeCUxBxsURBHJLbFVz
YLnp/sUKwPWYCXOhjwDL0Hao6K44In91BHKpGMzLkxVsAqLtTVSi/YKTA08PXBty
ra3E41sm68vnU3OxiH0TbjLobkKwopPvTvHd99Md8qtqD5PpTVmq3PahTP/oxvwO
tQEuPwba9NZ+SwopearjzgIVdgtw4zvP6jq6/V9h8j+rOKmFiIOTc3Ywmrr7u6xO
g1Q2ELFU3vgm+m969eKQ4hhLAOf1ZcGUNxKh/SnllHbvvhwku4HSR0N4IjTl1ctM
ZVz4iE6N/MMhOVMFnj/jSa69Uan743Q0hq14xYmklljrHL5rv6NrTVPRh6wwZQiH
h/8gTyhEkOqR0QqhFXmrAkrkzrkhyRgtntQWu16Qz5ORNpFRVlAQjhsWKmPoAFY1
qNnq6Er7vRrkTFQGqw4e9DS9aNjid835PZdl5uP7b7V3F+yuIZR4AA0KQ5vs9+F5
MDJF/1bxzDossFiAsGjN7pW+qyLtp4aNiUxW+M2M5G6cZOSFvHa3IPzmnz4piu2i
JYMK+cWQk9Ss4muRF/3ffRfo65pTafsl3GWzWiSv6AJOrctyMj04Ekkeyyw89Hsn
rtyuof7wB52TOJ/p9VUVnpbC4zy8Z7bxymbJsNp7zFO1Qru49F/L7bHmYLCkqBWp
I8f4/IVmiCK0opxlzHmLBFmJ8cpcs1YPAvXoylctQEbZLA6OQpQYwbjAqGYMwLkl
d4Ysy9H4xRiVytOOScesFG0svFit8qGTSP1rlxFEixQeXI+/PcgsPElDwBynKrFA
ktuw5WKwb/P7bUJrslT+t+BCt6Qinim8luMW/Y9OFI1OGuyjrZhSWFQ72p/evf8E
r7bnDWesYAMA+OnCsOenAIqZcqhWk6EE57RaMl2Tx+WHaELqCL04s8vFD2etnM/L
Bi/A8ZgU8dReQxrtknKz9YLTFib+SWN3fFlOxawIAX8dZEMPe+xSeM8NDnh0yrev
nc+x4Qj64I7SSdifa36ctzoxe59lq4JFzyQG2Dw4GNpVFmgGVKTnE0LyfB1znrWf
ihXCz2IpE8X4IhX9HP7x6T/8sYFjqrSR8fpmG2TZnLeqc1MSl2Q7SpEJHw1Fwi2m
62HDXH+wzzQGiuhzEddQayg6AbyufARHovpb1op9SPHaxCnM/jH5ThnFbGE8honC
GAVMFRL16RnIIdfInxtjiJ71j1IRj4rYxHx53L4Oxw3l2kCP5b+vy0xXnzUFI6Ix
oX0cQuiyZoQi0UN8LDB07P4AIpmp8UWPM3nSpaXyapW4MeV+CA139K4zDAjbRFgO
fqhMbNZkGPED4BVxaRce3PHeaVeN8sUUo4WoykhD2j7ekkS7Y1Cswif62y42l0HV
3elCESvSH6ZCFccpMGkbjZtqsbLe6GYdi/xMpX0ZxFNSq4fVCdFs2al4DrwPohJu
aH+7SIS0AhBvIzn2AkdJTI5AqOS29Lipg5gKxaXh/DktBgL6MKJOWi9Qn7rcsFq4
+BpC53dKSxZpGcstED9yVwP4jsUwLemGAIDZR9hrRb3qo5TL8mM5Dt9CbNBMsSZL
dHYinAbWP3qsumN1aTIbg8kvH57KOQp5Ec/FZloVgwcDWtmzSPwfVGO46Iymvl8y
vRFha4ghHrLx6pnBtD3W4vxzD2DjCgeogBPFl/ubGiZZriNhfUcLJJZciaRnIPlP
tb/jP5rfeu/ZcArHOrQ2K1DvE87f85YfnAG8WCaYnRAV9idHsNhGTd900Bv/1AkC
PdQaCd5bxj9h4ZowUPm1D8u1EZX5Pt+5AR9O67AUKZoEpWAti7lk9VeAOJBpc72Z
6p4D8kSLTzNXbQsjaP0y1kd/nIgVCm89Ke1w0VoUcqptg1F/IwchO6TMIlWoGtsq
IbkNzpaeA4FZZBwwqi0fqXdnl6LSjDerdi7XppZSaPHpQ54U15dp1AfiWjRMLTYe
bAkJuCU+M64eekL22a3yf2oqr0j/NJwYVVQZ5MtWc5L+Z659tzwoE/WABSovImU4
t0lapKq1gR1/MvaGGi+ei5kbBXSmz8fQCp4o6O5h1h31B18HlbyTzGyhGVz5OKzI
cn9TVQg3y47EiiEI/9lnEprOkhY8kRLXoH1n9JQCFOzGsBKsz8Q7kpxqCcD7Uqc1
y895iRNT0uU/CXvmAAXE5zcp4lGOD2eTFSWuOu6LZY0pPEKn5ll2xfTcf+H/4CMV
SnAwsZahy71mEZxdtVOV26+VybRXJVKEWiKvObLxNg5heNXk1nIX2m0FpCjIluql
pG4n239stmRxuxfjCtZrj8O3v5Mg2a/56Y+rBAeDW67CRb++wZltIxcIu4AtxxlV
s0NBNS+4UWayK4aoz2bhJKWoeeXVtTsAeKp4m4yAzx+V5IdfznZ6WlTarSvbAZwB
TglTpUOMpMf9a+0wZheb2Bdx5fiYTkRoTZcpS0wJuokiAfmUpFVnEaP/pCafE+WG
aj+MOEn1KH+b68eRD2lYtTULtU1F/j6cZ9Q3TfyRd6Ex/YVn1NDOpsbgqXVLCvAs
/QfWLGldQCweyZCK/yk2o44koXJ1mmZQPgMty/L8jbL7DvZeHYMYEmRIq27uCDk/
x5s0n14oUW9Qy1I/5cVBPnuLuoEmNVeVyqn4NxfwaUCZCtLe9/dVqnSXASWLWa65
9fxcCcz46Mxg/x/JO/DftWjWS0WoAuT1BS74YSjWgw5FbY4ZXrREx76Yo9bCJsQG
kn/Ltm/5FqdKXmExIfblLQ6WmHhMpUOhtipktL/CZij5emZnon3OVZyvnT3cu/15
1ijk03PZsPqA5258YZT+HY8A0C2JWNZSWBVaBIJvOiieyXeAm74pLB1BJNjREzqe
MkBx1hOTOG/SN9uvQqZz/TOgi31L+j631rKRy/BVdIzlkZ+g6PmQ8/fP7QGwN1yN
JTkizEBmxBgMDsN1B/xKfo29MSfVJOquCRIdkKea9MVH+9L+IK7k7iIoRDzwJTdl
0awfYyho5m8Txzw450Y2AxhUYhZoZjj4nUgn9VZwyW2C9HHZtGtBUdbEdzRap6jQ
IV/ol9W7qa+2BBSxYJQeAfIDuiOZ2ypIsaPdMIyx/ZzJ7WFwHX1SrNg4nZM0sOiJ
33ek+vqmklRWqE68VEgT2XW8xdT8Xsf+S/plEXZpxwbj2GrhWi6rTbe767QQVAdc
mpchz5XojW32xx5Q6VLyrX1nIAFKwgWMAWiyZpETHdGmHdZHeM+SMmtWfYsw/UwF
6EMr3XD8O2dR26Uep+LbuZVqHaFI1SOzBMwF0BcCL54qxfLa3aPgM/brUam9JMGk
dDZ2U1Ke82oM8HiEBMW9KyMv3pytDQkab41HDYhqix2/FoC25QQy9TuCcQ1zkQFR
E1btfT6jwV8T2GO7JwLzUv0e6KiRcWst9AOnI+qbNLFsOQ6wqc2lOzk4QRa0FodJ
LtqGQb0B+QWXZMxg63aneVNilZkCD/3tIDzBnS8Mg6XUdv7NOJf28uCB9wExQ4df
U1JhNXwR4MvTW7kS9bHO1+Em5IIHG0D/as0EEUR8lPi5RGlaf0V9MpjthUyL7rNt
ZPwuIxxENNv3ZC4f7MIaCGkEKdTbnWvXUBleoebIRLDwxGEDF5fCQmy6419IFYST
HBg/QfMhj+c/RnMhKWmS7wAxLjDViOjcDp2RYUiOegzxcuoGoOELbd94O31KoaKT
c7g7cweJ0dtMy1CQfsNnxBYYnYk9SVRjLYs0SvqhnmcojngdjTu87kQe03rW2YSy
X1t32dO42Q470XDXjbZ8MhhX3E955bNfpbWQ7rKtgJDAEh6WU8kAGeMqeBtD13FY
50V//6FVoOgxIg8mlFKB8DYu/1FUNDOzZ0L1CYrJ2MMBGmUzW6zTKmkrMIoC0ZU9
wCCimdZlM+yEuQvyMD0MKHS610ww4BbwdGNyfosgjZ5pljw+2qwejBQq+VpS7ID1
wQZ5s+M+pklmxD/olIX6TALPprZ1bbGRm0CDJqslBzsgIEDf5w9rA/+YfUL8IVWH
2ZPjWlW8yTC0UnosNnEqCOQNaxYvGxkFcxV3/ffFYPXHgrtYppUHaqrnuESjSvOG
NRKEfDjIkF5kGx/XCoHgEOnBEz8Mga/DjK8sO0Di8c14X3M8saUKDLrp2nYFRWUq
ouqrfFEoCF8l7bNDc0SkocEX7WckDj9eZsK3Hb7qf0lxA4pb8NriXz0F6rw+okPV
UD3WV+8IMfHCBfvSL3vOCVZJYIf0B8W6srCwL8dXqwRoiRPJ2CvUzjcW3K04za5A
HEG1UXoLRz7F1FjXb+N6VJB7RiXPf3vA60jOfp97AQkzclH9BEkishk3FiRDx7sx
vB4Rh6mUbTIhltItfxmrVT636yw3ttB4IPu7TJLBDmuD27qQeyrnhGBkjAEJAMpa
C8RgQpraQ9b18JZln1tEDCzBbsiXUEpuM+OCrMN2CoEAMATQ9FfyxND45UFN7fvv
izOBqjJxW5EcCLDLnPEnOt6/QNZpxt7D8O4doj193rODxaxvjQ6cHfJ3NsB6Buqv
g3j8iWkf8k+gT7EsoFB/1xNJbTFzg3Zs25vMgJkFcWbEJUFa8+8nlpVW1E5qwUtw
cJq7c3o6RZktJ0Q3o4vW6A3RBJtiO0fT+k5euXw20lp3XAg27P7l6eh5RZ+RalhD
FxAyMjS8KStON+V4ekfB6jZjB/kLSwwO2ZxU0waEztPmLo+CX3Abkc8ih3z1LLNL
W1UzirD6ym1/FBiy8uoQAuu1eCTjzIsBqFMJ8vhhsir/g0FTl/H/UdSvYDCampPo
D7HkX4lFuHr7LrhCzyFar+sXcMkkS4nZloF5EJQ5uFgR1E/4fIS2fob/QPR8c4SE
pdJozVGmxzQSx0i2Hc/LUdwjRzIdLzm5U0IspqRiHrej0Douhi7GYNOkYt2CA6KW
neNESjImykRkaD3DheWRQoQZJ/v/H53J/sbW53pkyEEmv3/DDGg7hp73oySivOTG
myWxxvnxYqy/4rwWwiI9ZCSLMMoXDMtB+MHeJVBm8EHfsxisxvBlM4bR+rp8LT2C
eGwgBUGFSkDpxfDI+VCkThkF64+NHGCB2DCWuBuyjW1XhBBDnPDz3Q6dAqBTqtTe
27oBmEMWp1hbBcoJuZcn3R6DM2AZvqe/aPnzj6HbTLQP/2j4NO8ZMUwvsN8YMP6M
lmpgxq2KLhK4l+O5zu6HNX59Qy+Zpi+4D2zGs/6Ql8A11N2TTci9tD+vy1q6mYgH
T/CztsGw1HZkx7+yonqQlf9InlTwSYl4TkIpW5oRCJfph/D10bfn5PTQ01Gp7n7q
ec9puROWVA0GL1raZQBEm4AajR1hrkQmv4AcqjpXNrW0V92fr1BgcTbAsGGTb9JG
bdFcRLCdk3zHHMyP3mujuC5/M0oHAkBzcoYi0wYYC7nQrqI5EfqkLLtirC6WTUTf
0RA6J8yZ/u1n0Pd7EOqRk3d2YJwISiol1rCqjKUX5dXp8QAbxeWCHxiiz9aiXP+r
ir0stkJiDEvXqKXN7RhiyJLqz8rLsGi32lBQfkZZhZndKvUbOLL7vwYFyBBvk4Fc
JuqA/IvwGKUxsgPNLwoJSWeDIAzLJc8huwnjZKwAlG2zXtUROWLPbNPDRMQrqVbd
ifUpxhIORwJ7xlDS2H+NeeqJxqnGfFFfCXccISIMpJRZbj4W0WRaYaBGzJr7ULOi
h/hUzIKpMa8vhlMc+6dxYbPwTnSxlSE6jxxPpigpnrJ+zQDISdHmX1tCpmYuPYEH
KWm6QomoupiL3iOg9oP2VECWPEkfC8uOSa6KGXspTcxtI9tbt2yg5pdIZYLJNK87
+bnh19rYyjerFD2dSBWdhCwPVMNZQTsHIWP/4urqmVK72P6RgxFffJLXraPgl2NV
NDMh26UYMIn6+FhHJf3/pYeVqQ4Gb5YPUq76TfMKr+tMX8eA8CNosvXmDgoRNqUU
mFEV4DQkKx7+GraN57z2UXIdyDLOdgTCNfbirguuia9jbt3A3EMKDTQbdADo7ne+
00xI2Nz6+hep0erTfexH7MngmsqsqxPJMXVkqmEuwMq9NWiYBn4eI7lUG/xqPDJ/
qeMGVxAT5TbOMqFRHIBCYbjgl6++N+KwCMA7E3NFGX/w49q3jEFzXp4JJYkW2zDe
7K/e7t5xfcF9gvsZbYKdDmf1AzQSXXbpk4rMSdMfsiYFgEmyYrVQ07j1TUC3Huzx
kxZ9B29+0pW0G9UrOIIyPA5DG+J7ENlk+Hq8/TMzUyecv0TaCdPqE7D0lNLUb3LP
7wDigRzHoeErzlt0wcFopH5pw/c4TO0r8nqfvhvVR1vPE6wZckmVre+NGiLeRrXq
TGcN5tbAymCnlX8wvqD6eCNeZPgYF50kHsBj9i9ioNGr93RgSQ41i5uvAoPdb0T0
9WgJ7vsgJPAkoglk5fXyg/FmWpKe3Fg5m7xgQY5HwuuN4NEi0YgFnc+44ptZCeZS
gpPaftzILJTdpiMW7QBQ3Uvy6Zqv0cOoyROSqfGK3fpcIt9oJTZSxHykShuT5yCI
TZBgpfta6KELaHErc41hzj/GcoPCyRmX53MUXA6Jcv9OF/BpI4B5qbA/S8qqhn88
e6KoO5xwYpmZuE2jfb1n+Elxol2G/4qgEojq+NpGa0I8EnTli/jBs1gehak8uHYf
ZbbRBoh8YYvT7fg7QVLrsTjzh3obyHh1nMi8eAT4tfQm8ZHkfXO7RuKGKqlg2Env
bKULf+0mJeZwn5KfO0e7ci8SNvhW6nsw7mwnSRcBTAiPktXJYHGQ04HMTHjUw9Ka
jhkjRLTXQ7/tWyR8pXlv6K0l1QNOwM7XdGZhETtP4KuJRu40ObLFrY5HGLnkvEQx
UCs9Q63hhmO6RCKbw9MX4dbqOAZskUlupvFcSd+U8E7xQqWIlNoe9z0Vh4rVnGd7
X+Yr+4Zme47vXqTKOj249UQpK67WO8I79ALxqYQ9RsOrj92DL23HrLFzAg6dUBVz
Rv5gNYrxAZ6PjGbSUGnRiwnyZz9kJIF/AKJLdkAeamvi+sjIvo4i4O3QNbvbe1qw
kOV0CkekMISon41xaezqgOwV92jgbPRZWKYoDMcekN/nmWGysCFrp17zgSj2dzkB
TN3faIC3ORD0uCx6jZ/6W1RkwCAA6p5iMWWg17crsiCn339WILTaZRI7XkFHMPTf
UiV3N7Zenvr3uIe916gWvvQh/26sX3/dL2XuXepfXafoiLkXRUxCsKzxratUxiat
uwaDsGexOO+fwy7G5ItSxioyoWcy2n0uprqrjAVteZzAaUau+8rgVzJw6kNmvlZK
/cKWU/g4eTzoffBuJFo3k61v5l85tqXdXtB07mP/OJvqTw7PFrEhCDysjGm+P5RV
RzX2TzM6h5X2+kCAs1/iEZRXocCe57nrl6jJ0GjJkrkoOaGSAb0AkTVkGgZ3uQPz
fDVKJi4DdRYfywotcxUKOUNvs2n8Mt7Xe6K/KqvEfanEM9P2IVGGQFW7UNgT8ECo
Y9Kfdh6gqhv6XJV8EreBfSGQgU/IEucQW3Oyceoki5Tw0BEZZnJ1c1rEODcFO/VM
w0UdsTbVu36U1lTuY4ylnkFUu7rCtE/2C8JcrNvCsI+yIp6qSs8G7NLa8+dzCJ13
uRnDlF0iKty2coK8p0niMEUsfTn7GXE7CA54VqgfN+D2Z1dnMCc+5wWPDo8a2brT
ovSyM8dqi78wEqWShFIZOAevqoArrWb7SCYb0jvJxacAFyb1zrdV5RtKJqyuWpR/
6ebhDS4YuVIpQa9u8QK/lDMuJXTT2gvsQGcG5J/+7SW7qYF6DhlMN2obP/C2bC+r
C55GCVyPX20OYXJRR4CJNZa1gZQjmTOUeshht6iO39AuGNtpceCwP/A3EwQ6Kdbx
02S0JJa1k5lESFYEQA6Kdg6YUIGzzE/P6JmzlkY8WQiUpzrCFFxBJsgQnGkB1XMa
xKEsQG/TtXUCCJ8P8tCbw+eJ6cBgbiKZkmPLpscJrbEPc8br3FQPSvcgp48SzUEh
LY3RZ9Sp08f2I4Wh+4dUtRK9uYbIycCv8nlsW63kUGMKUkCFk+9qKMrwwwN/zTKf
YHJSHqeUKN7nB/cPoPMzqEak4O1k0/ScNVksVZEkNL7iG7yFALTEGAknbQ0scW9b
pvGExqLNozYBfOyqOkAJy38ddrKIcNoKMRZm7NzdfURQ6AxRZaRoZGPK0GcT3610
sc/2ALGP6YZLseoP8em3O6DS25sACaZwuUTCph+OsaZN99nXAMPvKNXQTcbfSi5l
bsnFjZCrLkD+HMuWpQtVpsD1aTQ2SLTa2vB5Dcy3AGruPqQHbuXt29GfGuteehSN
PTPPqV/KR4BfJJJeS2Ilw8ZCj085EfeW7N/n26sKqySfWELg7N+PhoZoUyqFNTB8
nfgYR7kSX4GeCeyCIspC6q1UCAqCRHzdgHNn/PucDE4xHpi0JoRv5UjmIBeshR+I
GqmJeWQ7JBvT0cd8C3VC+yV4NepiawGQejypQXw8z5gJiGPfF1sJNIyeGH3z6N8b
rP9epjKjc7BSe+cAp8YxmmEYUMxmkmYfjqiyahgu9VAJQYVQrw+25WG/yEot5K0M
IZHW9+Fjfw8jc3f5XwG3RkIUYUnGShdsPkCafC/kESY0Jp2IynlrA4ijiExfvaB1
kXzeD/38C0r/DD9hYFGLSuUG6h2ICBxzuncUzPlGQ9o4rll+wKtOKlww0IkoGJUx
Bav6JrErjtK6hIkWSmTXX2xG5Agg4YdYOdmnVJEc19dBexTaOsinccWAE6/zzBit
LOxkQAGn+xh5Hag3xnftID5hbE/lV3r6mkDTg624riiBeP8Cq6bc6EhIWZOOn7qG
p84ttCPoJpy+Ni1HiQ5UhvxpEftngb4GaLo0yyaCQPGl5NoGuKetZmTQYY4dL6JV
GJQqW0akP8uIxRi4k4rCemAvaoYsQB5Qa4t5QC2KTQ9K6a9e+m0G6h7NKBAQW4ty
SLQG3XVaVmL6FDL3Y7ASLEoks/deVayhZfKMX7ajklFA2KFIotGPGWIYyHvBg8WA
bzO2YryOKaxq8dLfNZs9dbW8/mRQ6D8Of5LuFNUjCzV6SpGbFNk/RwqvQF/FzKOY
+S4xcfcVV8vJDU2uc79Wiu7xNVaXcGawFDr4+3YRav7e5GkDzibTy265+C06S/3G
ql55TBXpMS+uwMoav7H/t2CSLB8HEeYAK7P2gycJsqqSaTiHmrAns4O1oEDR5e02
ao26jIjvQD1I+FZOgMe+Vk3HAaR+slWGD5mBNcUz5vgRYtyw4EkT4oxyFCjSpEnO
0jTsMunKbEXZy72bh1FzXHMoiVjQGo9NVHk1o90o5JO0gs8nwNgqVEaQyz621FDm
kkq00IipyIOvJNl1ILgF/uOVKXpyZJeC2R50iFrEnS32ywqjdyE43mWqe51d1HX0
kjGiGOUEVENeQ0d9I7LHxyEgIkvx+zV7uLUTB/nVSHK6rk1vYqBeB4cuFXOWLme3
maHS6xf0fIW9lUh9S71+TN5O/jbKPjHIkFzbHluldG+TH8EPo+nQ9d/YmivlPXVR
8lMwJOiqXW5AbqRm5QrazI11EYoxZEPqzEErF0u8/6un4ysAkxWguoiw/vIuS1w8
mwAgp7WMML5t9hYEZjqC5/qCkU6KD5HiuqjjFp+qVee9LPPvhUxcTEsUsMmRno1F
9a+4s8sXYaq4qS5RS5oEwhOUytilbzNmQXANFTVeVKgsljzOXij03NCXKWRB86Ux
UtOwj4zQ8Py+boubI/kmnufgNdePJrIcbaeFJgt75r64CJNm0asz4hrndSkqf30M
uUbcPYa8Ls/PtJkGhs7Fwx40NEvxB62WGS+45qoOtCcKv5v2+pVnwKZr+I/cHZ7Z
XNyyByrxU1jr1Rrn0FfYgFg0qONA4tVWgchOSLwDNx5EaryR92b5bwslsSPgnIQC
bGtUKMVm0UNrJyxM0fRO2RuqzNxtg9fn1Lo5xGQBM89OUkwLmcRMTwHldpTUZlbm
LIElJ4octg+c1dvcrNU58D/DyAwswYNl3IMFOomj20tTvMZ5bIzMA5tNnjpTdY3f
M61urgKHjKz49+3BwteuIzBAkJSAr4d9mYI9TbtYHG2Z0xeS09HZBEIgF5h+dGo1
mkdOy5fTMSC7Q0zSd9mHNe/inj5AM1zSw3g/gtR4m7bfNZfGCmaaUsCIqM6Pkuk5
JhrZzHknzH/A6MCBWUmLOOAEHi9xscbOfWjnBlcJ0xFmopTvVmj6JSR/AxL6bIu0
16qEdQDiCm1gxNLTdERBzxZbaL2m361ePTFLZ6xUlpSyP60udM67b56EYq0jAMvE
YKykihq2QE5KHuXTXnq3grfSOX2GBzbY5DXFB5hbNQd+d7V9iXz5SEysjfJWI52q
vlau5yasEIYxqt65Hrl7Gct/bbAw4sRrCV9/dlqiVNad4CFGEpQ7dki4wtiRNxkd
SOoZMQxfZJKCdku2387H7Xqaj2L4MiMZWkfLadHyrDVGBpWMO/43npdRMQIDfOCc
CHBPJRqIkwezLlQ6yaXtrZC6LdGvslKc2efncOrvfVwKzcQsPVDZ6JRiq6rN1YBo
cMhbdhlLzf54eTtipjzup1qWGiZq1neJoZs/+KIiWJgjr0jp6Ae5aNLn1h5FG6M4
5Y5UwNWukDVaHjKYG2zDWWif0YGgupW/W0S9Pc5fpmYdWRIIedkOGNl+Q6bwPeDy
SG2Ryamoa4nI/30B9f3Uh328tQhufsae7dvGUtDUWfrLnd/fKWbQqwUFk5xzR2uv
4bsUVzowpN8GQQZWXxuQzVd7PuaVbkJhtT3kfulD95/jhVgk0leNWq3n1siSpvLL
0A+YNygKnfJw+rLsXAKP/G68UZuVeLt4WQCbWFuOKEC5OKoCdTZB/WsF8O8+umoi
6ZT15lCRqWXJFohrv/BxWKCxsH+LA7nNgGsCZTaFL4BT7aAX7TZAdeMeijjGv+j+
94TPYjnvt6sgzvekayeDbFOaWAsMKDrJTYLbG4c0cl3aCs3oX3VdMxFDHO13Z6+L
sx7lCRN9EGh9PtrU2xEzTwB20XbnApmlrGf7sXPp1LyVRdi9LkyfwFkAPX8ESIpd
nE8Cy0bWOlLOu67GC8pmdSiR4aHi4MN3H9khrlm6idbRuIECuuwBPdhJC5fHUsN7
czSlUHC+c4zIx55sy/OYLzo0qqGE+ME2xcQV9siH8EM2uuQ5nlg80l7RRNCx2pu7
rlQKPCmQoRmBSGfts39picvM4oo+66orL5YU4zUGG17zjV8pE4OXXZeKeppOK6Q+
McZwrstd5QinMu2xxSsS1o8LPWPMEU55/FyLGG1nxUL3XDAWa8/xcAxs5y3ZCAxk
V742pEvzp/9mQiaKMGfwmeqleO9gTQmlqaAUeC3uhlDBoYV79W/RIJOlC6OrofQ+
Bek/vuFWTo7XflGpBlAbKR3n05SiesCd4hH6gQ0VTJ4PfcohiQmCcG9Jkiel16wF
94VU03Vgy7lYeW06GLi3clxMS92ogQ6xTt6oOMsKSkHUjE8I6VQ7PRcia5rRBxrS
5yGWE85ZLN74f7tFbT/b76P5QwvazcILODTiqpmPn04JkR+Hc3ewXiqwLrV4jOnb
IicrjouKEQ8si6UcDcjEu6e08eJe1migWW2zC9aMsH4ScFRq8de3iq2Lz2xc08Zw
m2ZC8r2pxGMnnEwQYMe3nt3BHGK2INKUVo4IGkI3fDbZ3P1fVGis98s3Tq01zJTR
X01gRRltaJpIG2CGiFoZKohhr1yau9nWI7C3t0iSf/GG/mhAOq9puYqViTYfaAuN
4jv+5eFj9WEIlGkPMDeAj9vmhHp9GYb655MIFF6yfldo1l1vgx2Hv3gvSeV3zzmc
QmX5m0EyaQ7xwXcPQ2YoeeNfF4NiqyjJoKA4vq6pEUGjOreA8O9COH0vEDxSIxhT
BMxTn8TQr0wG8UXyqNdOTMY6mQXgVjLqXVQ1WDKlImc+dXvJoXCQUO+cV9rNt6yQ
jEvbFs22mbxTgnSxa/Tzt8L7Eg2+99QKPGtLDEKHOYuZB7bSWVyBE3XlkGFZzzVg
EuoBPQAWMMe/wT/jGsS6932fIFxjE3wF7E+pvMf9GG2EMtyj9m2mv54OBNdZP+mv
ymtkTs8RW9VRR+WTwcvE/3N4IH886KFW8qrHy4RGocF9vHK/wHo06bE3+k15uGeM
Q7DBHwo6MtvOMRDV5ic+o0ZCDKPzOWqrwwMK68Dj8+hCqbRZq1/Bua59XpOgOUTR
X4HqFGZSga3xX7jle8Nv8ZJ8neb6nFMojiyYkv1FstxgtncBMN3PmfJBx0yaZR+N
7JSO2sCatBHAwBqQPhFmG56Br1O7q59FfYxSwTnBOtXGV+u7zWE2xGtATq0zKWDl
rSGVNPVzuDCx+DY+N32Ll+K1ZPVK9jKnxxTC/P7tr2iQLaZK2i9yjoNL5nZsmq5g
ezLQ5H3RArXYgbb1Z9hk8qfQEdlqY4JWe6LBuRyq4W4Xcfw9rIC+aOYsSji4OOSn
kWfEDHq+VsVmraIDhojf2MAGfDWXZcvjFvz6x2TQLbNsNTBcLxwSmogfoHD9N97s
ZcjLFViw9v0+TlMYhgEJpzwz7VQGwyIkIxSM08L26TBxCNZhPqXstxDYl/TsLmWl
HO3fdyXWJjRNyCwTkK1g6nKu9LxYnNgBGJb/83zcH3uSi/QNLyEhj9PMXf+Snl1l
5GarwOWhzxHXT9iFLkSezFoeExVmaBKZ6doDV3o6icuBeRvkdY62mLFv+vA1PCdK
At6S/0wG98Vm2KftPWI6GX6muc2oMwzgJEBj10eV5dEkqe0pf50EeoYDZT6nr/eo
+rCd1s4gkZ9C3stRcApCATgBbkCA+ryDN/9odcy3yAMKY/sopYAVaQqLxeOZKdUx
ecxXEngfCxyfxpzMzFit/u7s9vhlNDMIKdvh/lm9GisYWqD3gwYPIP46B8Ok6dW8
zujv9y7ttk1jxN60MI4CxIzv9U+XjBfZY1K/GH9iyINvFPFlTK/Shh/5HrroOeQ+
ywlaqq0ZHW98Vec7WOfadhgOGmlihBI+HLr4XpOn0KvFEex2F+LQkrl4TqbTk4J+
ejGKKXcUKZaFrxADOB0AUPfOKsJ4phbKJxrxPVYcZtwxN4IU1HpuA/UaTFocE7eL
qHPhX24Zm/5yul2vwu7TRAVnhWQPOJ2xWfReDdT6Efzq7xRACSGfV6Ll7DOvdaC+
Q0HWxGVdiYBw30oQ0fSih5K0q9mO0byzaDB2TLGxIhaEU/Yu0/Sp2g+LZAHIrSaE
hIY5JUixMwEc2AjzDn/OGVQlLx53pHNuyzbUi0fmIj8Wbv90DJAXFJIfj84J2MWK
yVrytH2N6JenCiVjEP4sV7G+xtLb8gyze6PEoqCYPEYH7vL71u0t5U5xZjo5Pvwl
2seVfL3qcGqrUmPRL5qWn8tmQmEFCaIVD4l/0vN1uw0Gqw4w1n2jm9ZgaZ9GtPby
n/f677IxcjZeZs2KfayyVp4ZlPIq0L/9cH6yt1mQ0Vy2IAFK7YBpIRaX1T+B+Yeb
MfkphcziUuUYwrKdbIOQeaiuJcGPth5xTx7fUD2qMDaTpu0F0qertGLSJKJWyS6w
dMUC7bFFMLP4/+u2KM/awfLeBCjh0ieqTSzKmPMGnURuCldKz64VtMERzGtXuXEw
U7Kkq2lsa+PT1PylujdpG2HjpLwTpqLbMlIyQUqeucT/qDwJbYVX4uw4v9rsq2yz
KOoin1hIPedPTnMdWY3q7O/vLroR4Cfrb6ar2q8Te++wyHO5SBA+jRirfmLSI0Fh
hiR0D4WnQ6bryuVaDCN6d41K4m6dT6956GWtzfReY1xi1AJqbDToGHuDZoZGYI7e
nXr3xZKyYqig8OIY0m9nxM97iPq944ApgAzZUShXgA94GXJvzxe8CA7qyzCRihnm
Sv2yVxZ+aKJeZ6QF5iFMC8XNa3VS9/fhV6Ts/eKpeuCuaBAqgmzqxucnhp9jNMIi
XTySCA1G9KRKrUMBeCNd2J0TRzg2VPZnINz4zlsJ6iSNqBSXoWA6udfXtBvHmupR
Bft3KZEU4K3iFS2eRmMd5D7BIiyjLDFysDQtGOkK9JD/J8sSp7tGl+yBQ7tac7no
T8mxej/ItO47FQuKZ6o94ar7g/IZYKfySVroUX5EpSIYDI+m8V8aZ9cWov10Tccx
s/3STFGTzKQjoBL0ZIrN2igt5nMO1ekH/Dbhl5I1XgRKXze0QTMi3DZ9Wj0jgHzI
0omM6XYVjyEKSuwt6BwX09obDqIVm+cyIEdDGo/5xATF2AoSQoLFjfpeQZIjCpLG
QOSN1Q+Gg3kQT8gzXvhA2IxQOKQ6+VjClLgJeeGqBXZBLfiJFa2bVJKUHRXiKPgw
HdJzGLwRqgbtoHz/PA0IqPCuv8KsbkrJpCQP4LCdfjdIa0HfE/Qc3AuxwQTUKiTj
f4UYfu80Ox6yHT/xdL4elL/hXPwuygiarHexe320U/z2Q5vav/biva4IKdT40Oq5
jQNoDWWuWxxF5JeKt+bWO3o2kUtneTyoPEVi9Mwon8v6b0mELNojfUGdtZW4byk/
AwIyPU/KHKYKCroyb6y8gvGFUzVNGpVEG92WjCKoE4jSDYqSloOgObAHO3IkIJ6o
fDswR1mGIH3DEN1ZAKbfHY6cm2mVFSv24KZyrL5e5VVYGk18lkVQLLvarZOVWLe4
7kBiQm9vpJno31/uUgMo5JSQSZgkIkYVC7rhix4fLC+mlLGUNL5zKZe9ECe8WZPB
e8H55xSgfQaMD5eu8Dcgau1/Z8eqkIWhgxn0K6Auz3dZr3OZLtVXJTlEcDBmqDHu
yRdl751YUO8D/Lm5SLDgdCe2Emt7ZNUOKBjEuh1MPhRBdtgUSop07U14Kls+MWCs
SK255MLm15N2kpiZ+HKOg0wU8GjYsuomcDcY5qNCxODY7Kgarw/T1BhNC3P8ZJkC
WGF23XwoiHOm33Y2CZhPyAyF40zs+Bu+Xm8kmigSJnMPEdFnv9DIo8B6v0Zj14C8
4yFh4ZwMXLy4CWdlYEN8o9w9QhA+CmesQyamtAs279YGuUGSFT2qLf+SDt2866m/
xFbnhYx8evEjJ1kQmzKLxiaWy26H/nQ/YluI5vx1ms6JEOVxJzDxTBwzA/F9Imbd
KP1xSYxJ+C1asE1ksnM+Oie1TrthlCG5KM9UsvTPajFJOVeUpzjudipl2fkvQNP5
0Lf9EF2//tbaBcz2gKgeA5LLwZGANPd3I8prMGzi+wNA+pej2YHoAxEiy4oCNH5Y
c9dHIaE0pnuNqFhAO5X9KUAwzx9NKvfoue+fIlUAQ67zK4bXPPypyqONIre0jmhh
iVu9Z0nCJTV/g7IJWFfBtKS3NZz/ErD6N+r/kNWS4hf9Lb6BJkYQ1YeWhl0SKkb1
OV07ffMcYFVFzXyRSc94x+Dq6GSLVwNxIK6P+cNsM3d9A/jVnNPLkcr4tHw0UjCG
iSqBUI/UNw6jV4ScbJIbMN+yQ8hXLNntJokosQcESKblsXmKch/6GUEI9SerAtr2
eW6ofd6lcC3UhaC6Oq8VjUCESYmTShHW5rqGygoO2TbxSFoEgROohqRzzuXXDoF8
IhEeE9dDEnP34lEy55N7z5uSkDX01ZbU5eYXmccs5a2X2a1bG6i/Ws7udipdkItW
tYu70zEbxBXzEst71SW6QKG0peQxmI42HiWTvkDVHXeNFaCT/cU3zvJCbW5tCfp6
Ki+AM5cxQ5Ko03034vzZtWrrfQKUo8gze5tN/1nkKBCF3gm8/tqv3OY/S5qlpMyI
aMrRkJRBPSzwDdgbHEvQvKvAcSuSPVBOoDChu2RUq3APF1zzLvbFSwcn+wVIDHFi
53rRqT9blLJLywi0pK3hnbtkWNr6syKBefu8z9BVikVm/TNmxKhePI6kacWgbWMr
s+2si+W37fTE/YCKkd+s5DtoJN84iHSFCT/7I7KsO4nB1Kw1GINtdTd2dn+1GHf6
TeNfvrXFreC3bVWW4IB2e00NPdi7t2sooqT3yBvoV5WhYF5jJ9iBFSQ8ttL+8EGi
pMUijgkmf0Ctb9iA+h+jdG88PRB8iIPtzq1Yknx69IBuMqygIA0z5WuoVxhJGL4T
QO7Waup3cpLTAuIglY79gEYjmulhs/EYbhFf8O9RcczUQuIdoA53LiFE/0YGA9JN
KCKBN48Q4zXZMq8NyZgWDNAuJp6HDcqBnrMNAdUoVUVODEJRrJqAzfvfRUi7tmuV
DZV2mtY9e015aD0IcWCQG7tf+CCpLyeajCzMv6tZRZjws+uB6xM1ygGCqKZn8po9
94XfABLwMEqFIeS1ecnm4phRobrFKDCWYMdmfPet7CM1myi3UI+JnMWp2A0tcxXp
0GXKbfFlhsqGdhs1LNv0hQSRGsRhrjhIdshLm+wEfcHY5KqVEyFKce2q/ADBLR6D
LIiLCa4NRD/cffEQ9oUuDVtnbbYsWilr3c8EK+uPU7FGPN578onSaPi0//xsqy3N
0lcokw29bxj9MBvDCHaxowgJ7yqvtXI+TdxD49pqxsrztl3uKVvnfBJO4MTe2/ka
OP/PCVvfTNV0Z6bcxTb3sWlhq5Sb904A6mS1khlhM6MRP2XxaB5krsJLMFtDwcR4
DQvGj5zaAEQhX+rYcEyOoUEYohMBDqBhoeVMdLIj8b6lCdiXwPwT3kMQYbD2aXka
O1dXHAAyCL+31X0wfKcllMk4Hc5ADYFEog+SJJ6ZLqaoUB1Th08BHXiCT5Gr4twv
z3ZP/y0RwJR2fT8JExCS+UrNah8KX2S5H/MWlDDh5/ETAub13yLZqfETUcxvMwj0
pRWzIo6yEY+rf8ANxR0pS3eGwh7yIeUVuDcgbWHuhF8RJts/2gY4Udvk3jluut5r
jEQwZkvL7e0VtlXfJ2yMz4Fn0n+l1hhgO7Vz+CbBurzh0ujNTyHeBdZYVRpwgD88
qjwOzPr2M41WDWT9M4dnG4Tbar4SKD6IeB2I0Zo7zt+xZhjO/xVFdEr6XNHSJUGv
mr765OEhUCo1kxg9EYeMeQCe3unjduQyKtvFKQ/8SKtyhUK1nWIJL/c9PaQwRy4Q
GEMhkJmaOga1v6sFCUsccEbNxuzi6wA9EjcsHnBPj3Ap3kix5QJP+vfjmFUyY/s8
bmAuD5dkxIhAj7lHssNpFGmx4kLr7rtkwe05FoMo+y4eR2FZQhLW27+FcE3Rysul
Sye1wbWcLF1Ejhzs/OI7QOAzNGUu2+Dl4jHIWch3qoVkzrEzfF37G5wwUi9hAFa0
MVJfgJhUIGfeJyxp4M2LaWp29blzWN/u4j2jYaADrbGyUEmfwF+dFEhVmwrd4XHw
4yTW8PvodvCDAMW2zRlHueP2Nv0gaPL5lRefqvOSBJ7pFTh5ZefrokUo4hjrbA2J
+Oen7l18Q2+IZV6pZFMyoXJBFIN7quSchKy+ymV7GJtl5i3JV6NVbQb1xkwGBy86
/N7MoGJ+LIOHtO+JDxLj74ziDRLnXZ1F4brofOnyJs8Pg3EzTbpYGhpmnPTPIH5G
/RtdDoVEbIiW3omn9P8+JKoshDeLUl2fYxeWyCuGMWkqlLDBe/+e9AaLQ5n6kkoA
DBd6/780fNdpFrIOHFBCQyer8lUQF3i07TRPuuaYRgengdDfQdU4gRyGbtpjSOK6
PE0N5jZUDcLKhI2fUEWI7sYDpSap8jhcPXumNVEldGfHZk/fJwF5A0etKc5a/16P
70LR6Hl+eu6wr5uUIItnCY7/DCuZwan0Aaq1u8kuotb3vKheuxaZLn6uTu6uDFgU
Ev+9CgQ0P3uUyJ0jYc2b0o98Ka/2wMewhFaRB5LLTiiICJtx8h99w4Ljufo3lvl/
GGopTmIByROiv/bfbsRp1c/A706NGiXCZQzRpM4AvkOzZHUaGkWvbysASC65XY0h
Q/FNNDMz2jZd/s+MJlJhJ1dkUW4UUfr4qvLksPbnOqdogD2HVeLdP2erNL64ADA8
TK7yis2QR95NQLfVQh+7tJH5ZpIRqeJj/dAZTVovy1aJVBixcY+EduD0UNQ8re1h
WpxMGIgPixvNpy50vWrEwfPIN/MHLPxg7p7kkn0Y0+C1dOwkUEned8tvl7zv1i0y
VOXS3cqXmEb+PuZNFN7NdDclB81zWQmPT1SafHNOS9fBUsspStWcZwR/ErqdZnmN
LVcP2xgVvw3GKNyX2BoKK8S3krpmhoU1xgv0nQB+lPkxDsIG8k7Kt4KixLQn49Hd
bVbtVdwLYhES48VyjJeV0K+No3PzFpuQBP3xY39xO+oYYM1RoaD0TNXV1THACvGq
NOVfWWRTNueEmblhmnWUwxXpl8pXPK9gPlV/Su+2DgoY72rJb1J+DTdsWk5Q2xQk
wv+bQnuxLAC63QuwXhhNuK6sm5uUl4tPqrzK+e3wUUUxWT30uIvV8UwTODyZWa2F
KqmI0gz5ZFfBntP6+1PTlMqF9cazOBgiIRmlaXZML0wqJ9FBlt5l4qm/NOulmC4T
wVFgQx0lOXtTKtDiO5xaSrDGsisqLkTAPmHbBgThg1xgyVYRLSv6rzVydSB+uhYy
H1cyxVBgn+SRtDzEl0PnD5dwDCBsskwRP3/13RhKzRlNM4PCzvnccUsvbODpBJ6x
6vwXX7Tyf18pVMAryOQk9qCgTBIf8MF37CfmvnTsZDadmB3KfQuOLHPOYIXnRG81
RVbRuyH7VM+7mrOwi5O7VyK8CgVOvKWl3w5eXiOll2r0EZw1yIZ7IbJnUCxsElwd
p4FJqFjBJof8SKQsFzWgrWamzZxb46jw8WcdF9oc0mWnBgCflFXJm2oMwX3JJ5dc
SstIbkHtMRqlZq2xlucQ+LPoppLGqauX6szLxr7J09Q2i6FJEo2wR57jwzvtw4Ib
kY1u7Plgjf3zcowZ2B68YPq2GymxJg2hdip+U27c7jU1Zo/t0T4HeltKHjpog+Y9
GbvpsINwdxaVcf0rXc4yJpFqWDta7tGWLe4/oOW+SoDyfe2l0ZwvSFRI1MvxKHs6
xAXal7tFlCZ7/cyxnRyeQnwRNdi9Are37n11ydlHYVzjU+NsQw84uiyI4OzF7wjv
6Z0WwN9otThNk2LfhIgihzdls5N1sV/zh6NGwbohnafQ1OlnXgfb7Dkwq7Mw5XJb
aP9T9GAVtY6BCzR8+aKLKrH+x8yQrTEFbEr8LLY+gw9qtSpd8nq1XTtxlrfbtKwm
OSPSnjewb8XEcbCeNvoXoZQLmutJQMHaK/hMiUNl8GFtcnCxV9py+dlGlr/qOudQ
SAt56hIYfAiaFPsf0yiRVPtaY+OeYnGaZI7eMbvDHOo7HT5e5BSLJjY03gDoleQf
xnnAYjxsVgOS6DWnlTzCTl/YgWlgXxV0joKhrEJ2n3EK9/Hi3Ehf54KYBg3ZS2j0
A0KTnc3TIdKPTSD1KREf8Nsm4MfTGdF4dfrShJ6zqzmhrmgyPNJ/gAtUKcVrmnmc
0vl2qakemGiFv3eNGBAYyq6Dzd+2iCHztgBT0rPtGkpMAYYNdg7cAO/wGRFB/zMG
CCqGoi5AOUDKuF3/vkkxS7hSscUb0gkQ9yPbpAL8jwDqIVYq0htybh1IZqHDFxwA
Txkti0NS55hOMF78e4a/JVm0ETAsl/troU8boQxYPSQfobJxWAEdF0w/MbGqkjP/
Gq+3f0G/UyyWS3X2y3CAYWmOE7baamjYKPByZgvjinEGCy7217IlISzfwBHsOnRv
GTGG8zs/0CuOaHuSfeS/uZI+y7RDg9se/h8GfLjnbtxKQj1KXbanPTHNOm8fZeFE
uS3DBtVjCTtUEb1XQkqGXwkYrQ0l1gjMN70KeyfV00BMABhieRFJocvKybq7VZoi
N91S7k46KOOYx+CcXQu0H/Gc0qZB8/j2b/ymLV81D5jZR9Znq9aCsrgD8KKGK53E
wVzMGEBjzQGByvWWdh9B2CUHSFhLGt77h/GEkPtwR+dhHJLoR3fZXsgesliRtDRD
XpZjHgXuPgueChVM2mNyzSXnQ4aJVwAkf9tzGz/i2AaDqp/wfBSIn6JXUQf/BTsY
In3hOjTumFjn2tZWsWyMP3zCwkbvNG9Ha7wzpKHqB5b+a35N9mggKhrZKep5lcYg
1Jhv8suhBkgt8Gy4fRwJ3xtvBdMuxIxv+TTReeRb9AyEt/H0BetbSiuKkBaP4hZB
2F1V9CdLdxg7RktpoUXnPboKQ8n4Sspf6A+AF5UyrUnt0n00VsPJ+XzY565m3Qvn
nGyBTgLZ7/guUA12l0wsZHyLjkz1BhJpOnS54jK22c43kFN/viFpb1HkTx1uzOGj
PiedwBgYj2x3VErtzJjQheMmPfD7QsxhHhTKAfmsrKRZZWcXDPGVYuNc0LlO3uQY
XD9mTX/XeL3vRHg9/x5rfyec0/xzPsnWA5okmwZNBKdTFj1GZa4K0H0EthujbYb5
DY7QSOURdEYhm9C/EBO270xErcfk7VarzwAEtzvc0yojoSQhHls5yvtcuy4lsROD
alercUqOUCHlYvKEPFUEAk/RYnn3ON2kpwl4Ew+OkGEGdPCCUe03BNVxSI96snVj
cUH8xkE8iDr+3sp6/MaX9ENkTIDkraFtZjqmZzC6bxi+kS/pQw7c7uFfems+HblV
cacnJNGEADBkrGSTrepyHxtnMU+ZpWyPXSKnNsH8mXkHT5WdNsQq4noz08IYCCcl
lev/GFR++aOT4FIuw+8bPRtzrrT0IY8Iyp7mVt1qq1ExG18bIQrJtw0jmGtAsHhV
HPppgi6FLye6LMJWZj6pqcvuej+bZ0cZbEt7XNOJB/WT7AXakY3/tw5p5P45tvqa
r/tVVTUbBoMkC2v/TxPcS94ODqXl7QZFj/Kgz73PmJyaeTYq8dSfRg3umS9/1Fpt
gwd9HsyJVcA9z4eI0zeb/SXmTrk5Cl0UwGN+9iGl8BQThjeQSYi4IuBXnHIjhpVA
bRHnpiY206NI6qAd9Jr57V/ef5Utr0yREE4Dqfm8MOYleUatc/JO4JA8lIvZezoO
U2XTRxqWaHPdCYZSExedJ0EmcARSwjUVp9/3dWdJvxRx66srPq7NkVNDGJ+fr19V
9n0+jfqVAkmSR65fobuI3ulxgK6vvmnB8kHrcwnZ2Uxnogbw7fR4vshYDL72yYRq
AIeraQjPFfOUChUJrLNiQWCtG8DM+NDrwzWwJNXpArXki39gznxfQXwTXyi2dZfv
qnuEi6YVt1ne6aWq7a5aYKvd/le2aDzLl6rGXbgG92OzIXzkWTFFUkoa6yuL5+cb
Ti3P9D7ePbq5ZUte7oFlWBh9FKQcFNrJQYZgKnokyrY17HuQtKrtdifMg3jhjBff
HoQ2FbI1DwSz2e+ALAV+ARpO235m9oF+JOtKIrLeyKOJA0Uqu/fimd0bkhPEWrlo
w1OjnTmK9sQLG+hYT9dhUWtW25enX//T8t69xX/onAIcgj/2HYD24LqwEllMig3U
TkR7k0YoaLZDNEfASiiBk6Xg8CAgbwuWQQCZDIm8nfXnpGDcdE5FYkzcg7XZRIVP
7CA23/LXMZSNYN++BtiBXk8ki//yMWRjA76iCW/R/1tInfqEKRTMp8dhZigl8rFt
Dl8rTYoXLWkE6cK+EeIQs+XX5h9G4+D6DSDNUQb7da39Qz72CWOEtlBXRsgabDIA
QBjPfX796Zs5KF7XfgeG/g3LnQworbzOVwgLqampG592zfM0CdVo1HO0ksule03L
dL66wKVE0UbfOzDjIcAxWNJ9cHb8VbO7cOcN3PPMdKUBWISVzefwjFNq+zYK/QCe
ELdJvQcRTgnQdNNyZf+NycuPZKY8P1LFwjzwbG9Na2QbFY8FFEC2TJPl82I9FGe2
5Cys/XvFENCp8Nwrp5k+0AODjqhXem8PuewbEDrGBhqt+y3eqBVdH57YCOOKLKSE
2y9Nb+5syaKOrm/Ab6zPqSxxmUNNCjeSsH3FIbVzmm/wtwkmtMnXprXrGEvaNGy3
mgvEMDvfCOnzU/mB43sdWmpRn225oDouor0QBuGkvAMYI/zVK26SPJzc2w2MLJQm
zx1Ei1gmNVrk8vlo/Zna4hXzpRu0u1yq9+0uH5KAX16Xj0S3zghnBVoSwlqZHUdc
u4cAFc3SGZQdqIBfVtZLTI+WG93iJXtOHbJ56gY41AyCuI9+HmYZJ8dICIOIr64k
DPqLmMdy9YAf1WAT/j3m3YAV/MnIrbNbItAC4uNLPQTd6m0b8TwLccDQKxmZ2NVS
lVnoenJbV3b501QeYsfb+7v1uyZycTHHmUeX/Ule0GiMZ/u1jBmCu2Csfx0bofUm
6yK+oqUzfiWLoQkRFZENqm9ddN3PS4fKdOS8Mxl1SZnjPycyP7j+X/Rgg8hCaAM1
LqPLeNQOBSNn7xOMUb/c+Z+XD/AJNnJDjDIeX5Hfp4Hq48QxGDNMInGVlTe985f7
Jh9Hydoft7cojFXPbWTG0B5IQHPWGmXbGAYzpVpWFqcy/QuiiJUZNqOF56zffzKx
DbUgzlUkrWXQ4V58mcsyTjCCr3JmAFAUOJ9mIMkVG8Vubux2sEnstJhqDurZFwKN
LMzKSHs53Qi/42shwtz0CAATiTsZiH0TR5ZNJE27rf5BYk+aIX7EsGauu4WF9am2
4o0aob5+UxmTQd7HYSF4PpnfgMYqEQMCetMp2EpQYXdZdZ3jcj2b+ICuPqDebAfG
c6Mv+N/BvPwFkDB7MDAjfqCPrr4wYQFhgfOAkCvLg9L+ulcfJeEVstde+dP6FGK+
3/WYJnmQjpnvQ4sZZrb7d90SLHbblSTPUh44cwHsndd0oGuV0ugrTntUZBIhuB0m
s7ezQ5QTk1imHKYonk9EEODGn9Ol/BliQPnxYfaPFv5BMeQi0H3UFJauZsWZgWDU
6h7305pTdInk2HkOHXfYZPDvXcgHkHntJVo9NVoMXva6i5zUJ/SF94f3NHEkyAMe
ndnR2a7YQ+zKmDnCRrafLPHm6wfQ4pgHHOXsOWDcYr3jxFsVT+/hQ04dmbJsS1ue
Z3V9HU/TOsDJYdWWc8TyAsd0ojdUusbsjJ84QMuDTTlDqTGceWK647CCFf4sJNh/
0rQMWGlue8l7JFwQ3PMjZBVdD6cZ4gyKrWKmyGCptchXd3IHmUqm8XIJmCuM3Q/I
OVmbJsJzDN0pZ0Jx0259qHnnC+BCbFCzFvskvJDwb5mH0ruqWFthG3mHkpDUmIyG
sBKu1pJF6+lxbQ+6kxAdya2uOYbZ58nbw5MSVzOmh+PeGa42cHwvgEynEPiBkXg/
99ZaF2oUTWTscD3grczXjeOsG9GHH+s6E4MwwcmRSNWUjw9n/D/fOTencShVy1la
FQG68hq4OILr21PcBh2GddtJEB48jwjl/r/MHDpCSGLXydVzwLjhpijPpzVisPuN
7mEEAjDYrtXMgKB9xEI4axJuy13Jeb8IRg3xs8ALcL8xG21xp9s5+QHAgvluk8ab
J6G8FyQjwj6+LV0e0HvyyJ23tZW65g1EQvhYli/WloRZhlnHscX6kOJU5mFVadsn
MfkCtiZhCyeZhnWteSsJgB0hydXc5NYgdqhGkQnxLuQFKp5+LU9Vpy+66/FgjH7/
eAR65/n9tMVXbyIVIqsSSZCwK3Kx2rKOmbNqf7nnjQRJ1acDbw9LVSIFDY9VXekX
TqYYOkftAYfPG4zY6zXLth6eLMKdkoKL08pohrgX995Ha3nxu6Hgoj7HuOJDXHMv
O0ZdJLAIrMQWpV8MWuulCfZ7EBOu5I39sftQRaAnEcjdkSOqB6eiTd5ZGkHbpMbP
NxDZs1UiTTXMtwx1NFguPcBGUc0mk6MshaFCcV2NB2FQNG/yra17k2zP+6xOIma1
BwEk0lSaV0hM2VO6lxILyeTN9cQqcpKelLehMb1v1ANb3sxk1wxPV/PN3URhAGog
Pk2y/GxcJCY6h7UFI4iJDLs0QEmEJnj+OSy/nU6uYsfv0L6Leu7ydTmWm9CkeSKG
UbKF58izbOwaCf4LaesJRWD/vj0017MtVwDhKGx7N6f5tYuk9ocxyM4MKhzFRGpG
O9B7frZR6JuCGu4xUiWn9ffHeFnrumMQK5Nur4+pgf15OBN3kXQVJGtprO5UeesM
iRBHCykJtaeyZHz4+nCUWCROMydlD553CjGp2ZAAY6n9nsVHNUzRjLOm+N1xzoTi
Emv0Fd4pce2l7DLJPuiWsX33VeEHNLwpUn7fWNeJLmtvvTLw8fqHawAt1wHbQkDT
ZJPkWoCVHNn0/9T8gAsusPFPTElhsWgYIJFtTxOgpv3bGGLFwkHtvRGG81BjB7fI
SZCxP+JOcIsKo1bRyf7/PxFja/gjVarMtz4dvCvRpZAgppGpR1yY23S+EoZGYTfY
RYP8DFHTX5lMBfPdbLRRmHPDh3EIEEFtqEzzfDNlosJ+z1aDhqz6u/jMEQNFqtc8
W5go8g9i/tmei6LYQumKNsoOyRtX3Djkz3fIYpqK83iUJRB0mgqOOx+3JNPyNvNa
29UPllHfPsGCSK5JsBWiW7ed3UOhN/JESjULPlXlA25tWeD503KHktBIIcwWPn1s
jlvOwN+97Am82f5NdDL7hXkb9YDaT44LfEjih7zLewmFpNxWY7+cIhvqEuc5g85b
Rw8VdLz2GB4GtO7OLrGZJ+b37YlwanAXaoazdyvVJgN9+eeEjnoGJLpbuYOnXNud
gc99LBHAq+y0B7w2VO7X4/8v5SL735JPesb9ayEOitjU2k511iyb66sLkM1IWo/V
CvFJnChkEtamumt69ljc8FVSM4dLBm5kV2H5VYqeHcFt3G9pvpDmfvQDZDTGk3ND
1POrjly0eTkJufsvqzY/4e+Y9J9GUp8VAJ3gkMKnt0XPj3IfBzUYZxLNbZ993VeA
sJBeiL2gW/N5IEhKqH8MHwIIbJN+B3iOqcGAZra6LQYHPLd0p7Sqi3TniPTBLpPl
25xn3XhrefT971O5Iv0qwquIIP9I/ovKUnxTjYEkIaJpKuJ4iBBN01y9Uovm6TmU
iOAnZcf68Qh0t3BoUlZTL/ES3HO0NPPp4CiaTgcXR4l08eVDuJCPhUOcVLolrC6Q
ZdghEWUL9uo4+1qgYvAVzZCk3PaNFXFini25CGVUYeqP+Q0gUDAEAoSKMYkk0f3L
ZMw93tkoPcHd8W+4w/tz6x0zUCuH3bCooX/QgJ0VtME4Azd8alTw33FYPfzK6lHd
lrbM6ptBju88MsVya6mqPBMUxVCROg5kz/ItQalY9UR+BjMzENUMPrW6pzplE7U7
8nVrOBGCi3DhExEMSq1l8aCfWb4ZpXPM4BSbXIWAXwLO2LqzfYRp+eExcjMjzOFq
sbgeVQ3FT8poSemFfETSjTJRT0S02PofH9F/fAnyPcQeSAazZ+4WTjqrzMKd3f6Z
pL/rSBynutALiug1rG2TJ09GNFa93w8rIIvGVJDea+XDBYOiZO8Xq3e6xcduk9wW
wJZpfVWa+YBQH8nNXdIAtUQxBMI0Kyf3+2wjuXAcVFUiCcaqXmU1SN0fBMFATHBq
bMrxPG3bFIa0LU0ESQSjm6I9a2yGP1o1QgOHOz8Sax0xn3B6BhnfCjg4n3cbiIKR
qlIItvdeDGbOhugmlpsgQLWGMJYRaTwSZnpsp20JqRER8mOdXwA2fx7i4o2ju+iq
IJDZ+Kbz05bBW47hqNK/pyN84pRVWlFerj3F6WAxsyq+AYT/qcE6Wgks+4ipuwQ/
T7PL1PwCqsgud9X+GKvqoSsY3xe5f8zNmuTWf8ip0unVnRkLbLgFyMBhIuMII/zg
3vIDAhp36lGzG5gvrCtplSGupKfvi3Ra3uoKynwfVlvrakz1m0iH45NNHm8cmXHA
FT9mdfcXwr067Fa8kb2Tacya44zYsXtCgu31n4ho0m+qxYOVz1NxZ2aUBTjXDzTu
1LuJP4fGNsqsdhrg11Z5iMPtuZG5bwO3enyOwaswHc/kakcTKXRRM+iaBpatBI4l
aqEMpFIKXtkhayoRMHZNJUHitcrfJo8h17nmP3nqfXl9R7eqn7aFj+alLyz5kfac
x1PdgyXKOcrVqGSrjaZizjd8Qh6e69tRi010033bYRcw8smQXOUeMKTMtApD8wdL
o16RQV2VSR0DITnj6iUkob2aCG1kFUnAvVfT4dxVnhIzU9pSRB76oTQSqS0jdSmS
LmAcOzxJRi1FtgeEvLSz8MM19nYbyLCgmhlN45wVNboz1YTFZJhssF4AslJiyPSz
gzlo8djt6kn5WkxNZTf+92r7oqUWygsLev3ZLF3ju+JaGLB9gV0zwmnY6H/ccP3p
QsuTrCgIbzwB/nzd+o5T/Il1jzVh7G/GVoa/jTohHiQ8RqzyTg8FEP1pRWjlZgs4
JdXJtt8GkbBD5udlg12tHFLKCpNxaql4WkOQ3fb2vBafIZSRtTS5HT6T0TM6rONO
oh+pnX2WOO2yeeXPTVMqCAOlAf6RdZTxnGu441+ZG6JvDCv6/CQ1jb5+fuwCp87A
Xef62srK4ylhDIESwBHTwfefW2PM9xdcyhPGqA2J6aioWXDUdBTg24PJe6zU6YvT
y6uGN9K4fyHIw1yNTDcMJ+b0O3ObJiUkZNf3yIL5EmeLJh9jwFp0AII5JX8YQnPO
1mWMHSFmONtaxYqkVfmizgPwogQ3kxwWFu1doKB51qpfyShApFyPQVKukeE8p/tW
MU7daD3pF6tu9PApRwY3KDXOzldabbXGj+LWG+ndqpxfYV+BlKjN7EpFCtwyIvsL
c0x/vGp02znndcCe+PrRboSUargB6RmESr4vjPERft/0Huwv6hkAwFUAHPSkC1F8
4gtjeVkZYvn7U3+9dLbwB98fLXKKSEGfuaC7D94rygsVFhU5iVPs77cEHIO+SPOK
74V2QbbvQtTroZCfQNEDnyjGnLdwVgnU8Rhrc4OagQxl7QjxCLtckTG1CiMsmZEP
Rw13mRpploWfHYWOQOp9cdgNOb5+8+rBRUyTiIkzLim2Gso3KzGnYHTthzaxsI+W
8BOwzONKpyp7xvyNNMAi4h/3nnVCLuwAf5OEBb6Ecl4EPra/BchvF6BXqUrRRVfA
QP7/isJi4JoODWDnBVf0fS6nDd4YgU2/YsbwzM1wyaqt61kfh0xnzdie1XlCYPyc
qWpWHugm8L5JaYbq38C/23lUs62SUifDhVIVzDvRzHfKtqnN5ooLPOwv7xEM0eH3
+kDC36I0K118W/IHcqaMvaPVJ6XC4uyUXDM9BQrGyL+28JtTVuhrUeXubO7Liim1
juIFsbeujSlWAXH9fgk6GBd+YPw7lqbyzR+GHCH/jXyWbHpLKcvraqStPc7PkAgP
RNmODy2mRZQu4t3KqYqC9P1Oslz5z5T5JGclezsO6hJDgAXErz+LoVqCNWpCNvSd
W/q3Bw/t9gtpRazrWUxgjRO8QOUib1jYvA7SYgsTMDfrIHhpgTvpv/9FE/vXRoyP
2y2bw78Q4jIwSqJQAkk3cLF9gKDkDGSmFd1Zm51F2655Pn4Plvhr41S6RSkd92iM
O9VGNFeKbZNpaI/s/TBWdcF5NtKLWc5QgwnK1w9iBRiTaVatis8OvPBSdpFYbmSn
TRZV4OEgCeJmmH/SFI3cOYx5vp1wpNCbq3yvseof/pEX8vYZNgdzGXLpCK6L9IFj
PT3mCI6brDltwOzf83g8V49khCtHv3sbscpoaKCjgUjMHEm6Jg0hk5JIOAJcwJHB
83+ZaB8qx00e+wX09An75QJmrkPbZ5wSVCxNUu0I0O6OD3PF5jCKwIuaE76441MX
jwr2i0y9vqoIQeDNIrYtw+E/KUVdHt9dUUdF7s42ZblGGWtnk4xS00F4tMQZE/So
UhNYUCfZUtDaa4me4XUNoUYic/TTcos+7GjHizwiZNFs2THMp0JkLMwFl764iaCX
5LGIuxME0bbOkOg+t5Q3tRh36gBwVzHHgzmRS3DR6Yij0D+4cLr30BkwaJ4f/GZ+
7wLt9wvafHL8N/d37nfyHij24dj1rUfIwBRG5eO+LPWEyuYI6EcXl33kHdiSD3zL
n3hJg7/HSxnqd/SQbGWHk5jiDA4TjGH9w7GtoFdMSrTJfw3y9POqY6w8rT6/Irlv
I0+kEhPNoeDadpFQUHaLvoVnYt5wZ2VfdaOJhiRcq6dbqygZhI/gMSSxZT9+uxMp
CRXMID+LtT4cxFrOljqXadewwk6TB+jaZ5nj5XXpe1Pdi7tTaVrRgcfhBJGOWSfk
lmF2BTI3VfrJXnAtBHsM/zM46A2updA1lmS1ZtrvLjArxHHyx7R/0gdb/AYdcKrw
xXjFIQXZtoDCQxE9d4qmby+OJ08UffGyzhNYjJqjxGcAw8D4W3G5j/ssp+l5IbCu
i7mO+Jt8J4jK8bkvecrN8TYZSaFJZY+aE1aFLbknRb52Cnpf520sXRkystmATe12
XLlDdqtCAJlhnnsTWn6JKjwG9RGN5ZVOOeo9snh8sZNj8QTy0X+W3exvclFGb5AN
qxgBedeLUzG5gbu22zeEqrdshJrqGBIsSi2LFwlV4ab9C0kNSuqgNuXZq+EzDRiz
hfwJ8g/u4CzUBDDpVTBZnVx6zJGkbgwyUne2KmVvPXSSocTXCbgCl5j1iTkj4d66
uGKL5eMZveuWYChv+lozjg9I7ENkzVEPd/2x7QaRic/vqFQ/tyvIfEl41iINuOem
Wo4bg+B5FC+UY4/MAWntxyyYazzA676TDV4sqnrB+/4gLhIgeqHXHPMZVI3yvT4/
kIxDTJtxJ/H1Y4Swd8OwQV7eaJowr/dWIymmDNcnsiyTZcDWjHRiqAzCeAqAIDRq
0ZTwttV8YbHFkqPlkDjVRKtVOFVzO4HfCEE5BYX7QCsj8tas8gm4fqbdvTJe/K/E
GBIee7dRua8fXqVjcvR7FU504elMY8pxIRKmMxcrIEEk/OE35oiyXijtQpxqtUbf
PREViIpqD3m+hYm/aTfmbZKIIHGylxh/gjJZvzryLQgWP48TMoXnWGPnigwe/w28
w5Vx53f5cwkfdsVqdT4crpSIf3q4uE82GeeMLqfEEXEQQlH43zw6lGQcyywkcXH8
wnIfEv3OT4/OuexwghSLKQllx24xuoR4P9fjgD6dpeSg9UHW21qX1+4BV5NLPvHR
2Org7rec4FszRU5u4C44YBplG/rGnSr1HDKzhJRTPq/CWQjqwU3TRstFoIMfTc8h
sy6WwWezNd6EzXOfsaWTzgQchI1gqToz2LZRoxmhtyQ2+1C9LLp5CxHnSNUreN5t
V+pJMhApfYTjTbkaoh2zO7/i4NXJl/rOwHgHTaoLNuAK1V91dJTcPRNRqZyc34nQ
Srbvg00pcgugO4tOs8iCvWS9ZAhi87HRp8M6EqCrl7o15P7fZGL97e+EqRrLjj2H
wkOATgF8+xUF02d8Q0Zw5l68x9k9laswBiHz4KHiYhta2ORuMA02f1ReG8tb0ovT
gMLMn7ekYrB9vOWtsZdV7UStClYN9Bhn7K/VXx3ludHjsM6A/wiiLf5KJXDkzo3S
WmKCa03g5fNy49JlujbXuMcuo1s1J2+xBV0ipKUWdQCWPTS/3gOdeWlIKIxLKiKM
4/unVSAl9bnEXc2+31bON20bNlPlOgPzTEQyJFkQP0AKkZXZQiS9eepkSAgdJDVw
SKYfuPSU3xQmxyDd9W/te9O6kC/Ua9aa0H5oPB3CC8PgUjiFHZXJFzv5XtRQ/8Xt
xXHX/hF1hrgY+Ov9Gj+XnA+9FqvllHppRXxwdIitIpa9xDQ04sefWSfFs1c0P1ZD
IqkovwI5X/Xeat2U8vbqGzTVm4//qCj1jjiWglAg/9SbZ7L69WnB5AgCeoOvRHS8
kzEbT0dM7i1s7nao6Y9t4pJfUIl+j8KUJnRpiM/jq/N6IvTQULJSRvC7DtsgEamr
J19JLzhhq3zIdczCEz78jV4WzLKfvH/Fx0d+4RW3G2CIFhrQmLU4ey3xBX+QDFG7
0lr6diVy8LlLSkLBZalMO/nu0IHVlQJ/i5AK47H/G92MIfunIIlOx7bjqFGU9JEM
CYLzsSiEmcVGQk4FIU36EQHkAvmgr+ilLkqH9fuNX0008/Ae1drznyWaXNAq6gBz
GVb+x/FIA7ZPBK/ZexF/iPFhDn93VP6+4qgVa8QYfACPf0T5fRKggwSRSyMPwAMc
PUPPrCws9Xw5mjInRgt9zGRtBKBJ0tZr/ukYsP/1vrToy4SFEGwjjzd/zppk+l+j
JU8xSeitkVYPWkY1qmOKRsHi9JS78Ushl3p4pMAhJuh4crPEde9fcS91AUTv3VIT
HclZj0xT7O/Dt8aUTBDvf8adx1V2JLBYBJTSv/1rwCFD0lqIzKayFFHSl06oaYVK
k/TOWCcx3JVMUkMtNqWmXgViBtFdWyDTXO+ov0gl1HWTzUsRuxXA5WjFAm/pv0JN
7GfCdMlo5I4maOX+NLvS81zsII5oOqIhff8aavkKqt85Rbd+4+3xIyG2jO6ugSdy
l+s8ZKAwU9od+CX0JyU2WDgH5mrHqrJAEH2U3MHBQIBQJ7SjxYhdDhAW7QMu1CHS
YHstp/ns8BqQB82uQk2ydgS6Hgk7NHodz/maRcSDhJNCatqoYcDOslYIkNh2wJQh
ZZ8yZP5N4Ns8+lYli9et60cMGT6X9Qp1t1ChKswp1pd5AbMPXiVjtWcFu0fqASbk
/PAgaUqq96l/fDtBkqSSHQEH1nEV3DOc5H51UKK2IFHXkGkpvBmx9kQWQI7fq1sv
kPtKLD53dAJe4xwk9wj3oVmsgm9S2NsIDLZ2SqYDUQcrWjYrvikYvR5lGR0oHwo0
jd9ORXa8dePazTS49Oi+b2Kswh83aqZ0QYR2QR/Lc4+qmNCVD/PJ2cu8JhKfGvPg
TULgiJ+/fwgPduupu6lI+feWkw9hP4wBGQPWzRcE/V33J+tcBugpum3cLigfkJij
8WlSv82Bm8BE7ztfRfPuYcAasMWPz3PTBM/jSyKeKMdP3QfMBglblVKqdMNLq9A7
u6s0EnqQ0w8sdlBNNhSCXwYASLeS9eEsXp6wGdP4itevQK+bSN/59svkvDzmCpDL
na24M1idtXuTCVj7mc+vF2F8JoyjSv7peXGYdvRK0n0dNUMGSLKjCKs/FYVDtuMn
86zo/Da5kmpgIz+QAGlEUQdII1x0MDKQQkqab2MUO+lQtLdK4yRXjiYPXQKuLPbh
mgxPICrKirnQyrZdmEOWEsYrbQdvDQwaICqMu+SJr06xJRR04hUdwOAC6wDhM4m4
eBNT1WlLS9/qFSw8KmjpSxyxnqR5HEig2/RR9hnwxb6zdq5IZrVT1AGbu7cmkONn
dr1rG71qiuJ2E3Lwq1H3iwG5Dsr5pfJZ+EiRpd6QkwaDs6etm6j/huy85/R7DNPL
qx8H+LGA9xCtoTrnXRqvKXcRCtYpptdOY1YQsqtV4eVo81ury4MEBpwc65U/MZ3w
AG3LsN9wdGFwlvVOJDD/qAHVL+eLkTlwv2TgFTKnOqNwqoW9BjlVLaBV+aZtLIv7
CzkgEOMLzdClM/BSsew+4XcAov7Fc+yw/3OWEcMIeW+N5yBsH5UHHOqGmxYDpd0z
rpMV8i5r75/BI8I8v5RGAktvr56WkCSMdVyIlzLrePPb264ouFDtB4RxJ0lSxVO/
eg/gKky5ntdpEfrxNmv2cf5Cy8zfQcrU7Sg+Gjkct/VCdnr2ZGxlolpslQlFwK5s
2Bv1Rq2PMw3oafyczpvEYdrb4QuydUkf0vA+3WoEG4h80/gR8yECkUQ/ZjLVqvni
2+2eiAo4T0D40ikpTscOt7ssp/o51mgPZHfX9gwSHZ7C5z9cPWQM97H1O0x0QNoh
xVVXuPa32JG7HKAmtpZyAN2YqyX6gpEWKqOyQItCDEXySoTdVhploiK45gJguKUK
1hFfSvtsXmevNyPZc6GR/TbkS/q5PpqD2sRy1ND6dD3D+3uLEo/aOwxOz95DrTv1
vVOA2twW8tx5jjHILSqYbwoRcNn2IQV7WOhWMRtetpACQgrqkA0d+jQhiy7nv7jB
38A47+FxBmb1sUmPYKr1AyAqQ7vxlSk/exJ23Sry32D4OVI9FRbUeUO9kQ1gDtDZ
XV4RznD9p4QfroqgWe5kennHe7mVC15VZUZGGhWk5ha99qsVOCSrr4y0qdFJtmqy
zsBOIWZ0PBP5//OnPdqxlXE2Asd7hie7DajSnrhY9uwBz1N7m47/DlBdlGFBjUQo
dqa7yzpLOhb9x/WeozAyMLudwW+EQnnqontaH9/gC+CMKkW0wNsVXLeSQqyuZycE
Pjy/5h3GSQKp/Gn86K458rB7f7dpfpWUFcKHkCVvaprJTu8potIsxspDmw6zABZC
hxd6NkmIV5XhrulxZ2RHRRJSQ3zGqYd1fG+YbIAAbRt0VQmz0dcDO/EtCO0/Jii/
Cm0PWDqk4W4ZHNhTOizwCu3gq2XSl0Fvy5O5HebAl/he1kbCLBVaawQgPNo/8fGR
SlES7Stu3oRVws9fHel/tr24zlg5domytfRicsO8StFGI0ZvNR+fe9zBSi9jb38D
Zg+mTmq02UBR6T09KM5rXHA6oDm7lQw5FVJzeIx+FYe6+tuI38ul4xSo2zqOyICa
t07+dk09EB7AdJzIU0mH156qtTgWVpSdST7fuiSd4jPmwAcYI1Y+Fr/nApStIfU4
1RjMj+uBQcm0IoZ2bcOJVdw8oRtUis9S0jn/asawYXARb6xdIuVUEVG9uTH3LZug
m6I5FH6KPLX1l0qVl5xtuzom/AwxQ9ojY5cayTBAFvIsHlxZmHYLGQ9mtuClJJTl
qse4HX4XyQO3RK/fkzoK/4q0xZLnUBrC1A6zsa+paPPLALwsx0dCg7qInbEW1JpK
/u32nF/M5iWfLNATwFV7g/CR9qaEoEbFuqTN94UgPKJVenDwOlTaE30atPkjT2l4
9qvUCzlorTsFdUANYpHYi5c9CzCQy3++HEvmofQqwsawhIYdgNeHCY3LrMtGRSbI
7aFeRIEjpUMOe5mgZcgEC9RhNkkMGPwxonUDvBPR10RP07i1d1axCIWxWrTny2R6
fAC08qMLk+MGtNo35Et3DH3ySM5GaAK6S+bhDJWdOZW1TY0NF+LhNHW7aa/hd+kM
bDrGv+iFuWqjlpYslVWJSLdivgXWMEBm9kGLzlyoZ4sLZSVk37Cyyry2/RreWz7/
9io7f6SRl+u4Tp+xfdeup1SM0S8y7NHcz9YR36g06Voeagd/B/lEVlzKeGIufZ4E
K0BzkrChcoj7bvZ9oYXlkG0mVqND2g7twMH3HMI0x/T6ZQabg3r+akhbrNOftyR0
O5IEekfzc9Ndt5XQkmd3tSvSdriUp/KEpCmhbE96fhJPGfz+Lih6gHmIiwf/pQD7
dAdZsbAMwxDyD/eNwHf4TPndGiTl/lwoJy4nknSBhDmffcQ7qS+YoAm/nCJ2HgCs
DKOZ3LlqxYUWJEV8XT5DqOru69I5adVHnMA+RTU6xl7BxkSFgz6lOP6159QK3EWB
RjgB8groEIpowOaiFM1/QTvESBE9FuOXobFnEzuq5vEYwBxl5mte1p7Frc5Yg7Qy
TvA6rsSlt7S52TShAIEHetZ9Ne5fOBjvrUKjBLrLYF3NE+m0tJ7o3ny/+ssnRCyp
fK4xHSRLt/Gb+YIK0wWcWQwoIwMIBeoMFxWvXJsqryv+sas5KqPbkgSBtPzUeEgj
kqJFKbmz5q6ZZmNxQCKBMuH9AtgOkXHfHYn5FRSqnP2ynuXMf5Vxh5qkoHTdZH3C
0/NQuyu0a4GnmbBQLRO3Jbjx3fChbeizYeudi4gyrBJrRrL+jpFhBkycVDrpaeKO
i0Y9t/qQnuSPPsE5fDl7yHHIKFbZicN3TPEX97nbxPhNVbYDdvcqXTZLFVXBhy8P
9Wg8pV7bG/hxWSQd+jBocj4F2SlbeRdOXhwVu+ho1jN8hziWSDWW/06p6Tj5Mx3M
NdC94tkZaWEC0xfKCZNRfNBKpr1mSQbAMrqBR26A27EYgrVr8QH6hZXTaPafPLfr
u6NHMFr3bWNRxAxazKWs/xGfsh7jx+zFLiV+MMZYCBUw+2Nv4zf06jsH7UZ7Ae8z
xGyRC2Cg2wdwe9wjFv1PHIEbDL/ZMFT2EoemM+0lSgqT7Lf2K+5J9/mn8kpzKfQ6
ZqVrl/I2FdBT0kQD2O8aS7TjLzzVqyG48/m5NvOkZVYMGvCkzimQDs0Gcwd0ONEp
9eVj92GWC7I+k94WGw/Uy6LUpDLHf7gZgvOXMzlp/X9cyBHCk/qa3PTUHlyhUgXU
GN9WFTeUGFLHjCMk4/126DkC000QwIs6qhds+PqD7AxBRvQsa4NUpqW6Po/DW9PU
HKDxFJf/WzA/xbbA/mCbHkfRaYc0H7NVPtLKXjvGkkKaQvSvQQPLIGFMgjeD/sCz
fwxYe7KFA1xSVg0VeRAgXMACmW5o4bJi8lj/nejBVKk7qhAureVm+ygTKQMD8fyA
+G+chJOgZkn/pZE1P6SCz1PxfylAAR1bmOP1vNadkP3KPgOzzb8wvpLoXxndjCxp
BiPkh1fjkjH1nYarDmEIrb9dnBBMq37hzaMq83rjXAy42m2Qff+XOZfImGb/9bsx
wEkEfkTdxKNPCqAXX3BzU7dE1kpi7I2z9QjaoLXRduouLXQIgiLy69oDpUTgT51e
pDrz1Hf/8r11AshExrjsTUstGVu+AeXWg6dPYS2Jno6OudFSxVqYRTkvbmmo9ucC
UNsXk3aWTvOiCZMznNFC1d3xQZXGfOY7H6QNojbTQbTOYLAJknBO4O4mLbXZxJmu
G4nFJ9JhtYrhPKr1O+f68drAVUdb3F7bbV2QnCN7EZnSOXKtk6RIdAN/zqGSTNjK
1cr1CwPXw6+lRlm8PGlpe+sTlWeylnikB+W1f4HZC+DLIJqBJ/yI05v20ZiNgnW5
he40rEqtSZaEoABw4j9CxsGdAxc1ntx2/GRdv3hpYBHVWcg29WvzxqJX50YuehDN
3lZ8t7O/nlDcodZtKd5cJ/JGmvZdyRuwX8D4FNlTzVzxC2sv5Bz2VLJOgKFtvQ21
r8XZ6jAdrdGPWAouKuGem0o207hTdQ4hn2YT1qJmSXJnvk3yufqtCSFat06IhjJZ
6usHEULra080bKdSEJDR4fCBvT6cKzVeLI5haYvnTcELCx6oC/cTaGsvT4k1fnsu
S2rSIXn4M5ZOIYwd6+qMkIVlV1YMDyorLoNGhZcFD1teKEtFObl03nxl6xOPWM0i
dVnWdAJxV1fPn44RMqE8mo8nPexXxvi4hJ2TvP19RaOp0nHEsIaQQWPSkrYhZZVb
tWnkSTkd+LIqzSKRORiDxotlZqTQOBNcj9xo8l+NtY1BDmyoOEH1/7tPtkrDJScc
6np2T3z1wmG7/M6iAaH97nCXmuPBh2h/wQfQSFsIOTtwUoDP1XMBgFlms1jF8qHt
lsz8wdx5bB/Nc4j2nFAhO+XIiBf8F8JonyMkxAXil/QLvpOWIxt9E0rmA7/UX3XL
YntGR8nzcyKwwZdh5VZXiFjKsc3uZvDCrzlm5ItHPEZK+7LYm2yQTryMA443H/3M
rRq64f3FIea79MJ7dTgQscZYWF0kvYLvf3Zn51DWsVKvwJjEuL/BjbG6nP3hLexu
ZOWbri69/Jp2q0YE/O+GUIkmrfclm0gdaK9xYkg7E6daqS+vt0Utv9CJN+U1gJE6
2sU5pv+GusfE4huiRAyUhlIKr09DuHrXkgIqN6gSbrO5PVy3xFIB65wCtU2Cn3Z1
vK67PE96eKaspclanLJLnRjPsMRS7EHKAUZvtaePrDmi+8mVAj5b/891/lupUzJG
EHclNXoqwNvbuQt4YVnW2cyufoCwTZCJrCuIJIfOd2q+OdL8C1VZ2vK5aNMHWy3o
DpIzO9uBZfWSCJHuSs6RKMgctrG3ZntnICNEuCiuhatx4nZJPqkxJpSZa/2DHDuE
RxHFViaR9tOjdgJrEOZ2EmUZ5EyG1mPkMjUq1OyQF2ZAZmkOgWGj7LhMT3FUBBAk
/qQW/rO+V599VH/xZUmph2eRvy7lFpU+LjmNjuffLUXQ8iir8QkEP6bUq0IuAhRt
lkpvHasOkt/aCdF4G2qu/zpH2+OFo5tPgpWzFbiz2aroCdtUt9ZDHyejY/yjMyJw
gbtQFptE4SFCulHi3opO023jI/gK2RBRHUXKTO0OLZ0zjnuBKRavqhhHRmrXfAxV
oqmTJ5qK8QyETEiXnaJNY6xtQAmhf8JiAc1Nq4HgezhXHEZRZNSVe/nskmbyL2gq
KoLWHQujt+QXLJNUd9b6bNuG3LUdLIF1L4fDL1Krzwr7KYqneDWxdOmBA4mto8E6
WU5p5U3sGn0rQ1Ib/rFZvvE2x//GTz7IMMNKmwUNyzcn5waFPf+UAktAzjMAMIQD
UImOTKUiukG4xa03T14/rIiXRJQyomlIXx/1iyrWM9Ocob+7VnWEV4I3l1gh6AgR
2qahUjxxqAbp5WPn0Wbho0n+QK31FpvoSwDdmjZCQ5bdeX49EsGsry+yEb+qbCRn
PyK/rrnpT+T/+KzvV2ja0WQUEprg6llZoGYVY/nVrPRl8a28Dw5Y9SNokR7di7oH
FQf3XHCpJwiABLXmt0pGWA0hcbdvKgiDrVrtfBuhYHqiVkeakXaZJ3QCYwjZlG5g
OCZ1lx+0EoGv9dGZtHMowyQz3UVfGOpTBFhGOSLA1NV1A4X0Kk+QrVbLSiMPQmD9
IIukVu0Mmd8YVoBUK2SJxQ89CHUBnY2ly1NmriCldvLSeUwrXC6WG03EO9gyuwRU
Ws1vjg0YbSc9hrOmhB2hUrHuHYPi9er1xnClnT1/9eeXZFGnyIhrcIX/WPXyeeew
e3H5tKIkbex3DjOfDUiYOHMnbnrXetwK2RSLirNG31ybdlW6HQ2d9rFRAuLmEgp7
9tehgx2VguWNqULnrAN1x7FI69acZIuD0UHj6ZmusNB6otVSrMNTTIQP2wi+5k3P
oJbE6glq2TgCNJ1trXwv6fYpd/m6VKiH9BmQNdeMiCzzs/vqHAyZ5ROj4W2Xf/xL
O9hZUPfD6+hVFiG4b/SKGcqQZG6z1t0yVNKJ++wnoO3hzUnmDjsy8/NOBcPLeXqP
fUYZbUmsLcoKSEJUwlAw0qtBvN3WCffwP6TrZEHI4Z/XqaaskatuO+3Cplvedoap
PAA6PRgFHUa3dRUAyd1YcYBdj7nYThq70Bnd7j1fRbPRUSKCiU8C5WKVvZnkng2N
IWbMEDqYrr8kx5XECJAA+hy2lhzGGSKGx/aMAiR1sD71GfHeiGk24pxGjeP5Sfyh
riyFeYDK/X6xjnN6P6g6vLlRF3x4L7YJhT/BEUmVNclusd0UgaIm29Q4lOBhpN7T
CD+cUGn0hp8DWFmzQhF6LG7DCg486fQY24WZD24gia6nFVCkYos54NE3sXssRnXm
DlEY4Bcj7cys4LK02sN2Sr72U2hPhAy/8xnTNBxCoMorhheX8ivLJy9thMaJmmWB
T6vvF+UYwCg2bxgGh/DMjFLukG353yrvSaIHYxskB6kAX9joVShtsflPUji7zU5D
tvKXOW1VUDqAcOiBJcHy+H3pa60Cqem3peCDXuO/lmInQudNL0OFLExEUy6ZS3i9
4BhL99v2/HGuho+ZJ6xloziSLCUIgKohcO9IEpFPz4XSeaSH1K5Fr7cYF/j3uSt4
UMFZQFVEzp1zpJzUm2aNBvCVBbBW1fLSVIp8I5+HHMDQHO1ZuS0u9jhHqvsZ8Qgx
ZEm6+zRS7u9jqgOuZUallkezQE8eisEhANWLEAx7bhZ3U0wYqYSP+GEkTmcK40Fn
Y2PcXt2jG8rrZfnNljNZFu4U9Y4ziwM1T1cPWlrZGDr2ExwKOMl4/VotISBk53/p
f/rcavVWmWWGxrLynwtREqhZEHwcp/EGOsAOM5LpDcoOIusPurSgFMthaDpPyxJE
y9qdcBUsd+SnA2K1zvdPAt8i34/5J0rZV96xqmkC/X3sv+MDIIniw0fhZeKWjT83
e2OMCd07rhHOW5LG7q8eh4X2as6vcI5u/cXsuqcjFrQ4qcdIqMahpV3xBm712/LC
+9SeO+Ne1siRht7y7Borbgj/Fka+koo9TgkxPHIfdFpJUpO8hpM8rjWLgxG4kncv
I1MHGDa8QEQ8JFRTrUpf+HO4ZCXbWXyi90UVDz/eQiR0Vs3+AdViCXwHbWaIC5Mp
O1t5dmKU1MjH77gbpontIWVqlz1rehun6zfapJVk9t+pJOzzbsy9ZTUdUwyLM2/6
9zkGUlMZPr23Ait5fa4gsSnXtdYCmDQomsJzSP5Cca283LfjmsJ/UMUmltz7JbKJ
laYySdnoJ45H81qMohS+sFXYldlc1qvRtMTaJvtqvNzOgszYbBxcYkc56q3rc2dB
fQFnDTkNmRIZRtV7JrLQhxmUoKTy96T5JSNkOd1jWHibynfVLNVtlm6O5CRDQ5px
YNzHCOB6Gloq3cu2Kr/YK6THH0FFlxkrhSdn3MgnEeHh6zikK7A6DzA4cT/aRuJX
PiRSAd1kUep6iZOrl2EwbJwndm6UeijYRx+fTTXGyZZB2zQlkSwStcSCozICBrN/
KdH4Hv4trCk6h14m6b3zi+eYC+w4Sipf0Vj2eXXiY+C+9k1cAH202pJ6Wo6DdGrw
ikaFv0Ia31RHLqIvcXEivlRrKqcEqpz6iEQndJWGlcrG67azLp+hMPlFUM43ZsBN
DtK8c1Dqqk7adWumhjlfulHch+o6C+UN7x0YUORXa7MKG1jAHd6mZT0Tz4cBteha
tZKG02naHuBShcQj+a24IeGDVoDF76wXCcmgV7xcMA+Rh2f9zPbT63cCQQdJLUCm
ooUd2WkJNKlo7NAlgFQLaDsFfqMc5b0z/4T/HkNDSI6FqGMfGzj9emxaplROBUL9
oFnL+Y0dOz6niTdr08sAezXpu06qiNmDgKGdZLtZgb3xpD+4wcvqzgFU3m/MlcB5
x3pbvu1+wMlM08fD4kC+uLV2FOQMGxDyUenEEnSc1t2T6cn1H4epuAHP+ueENeWQ
3XVRt4hqH/0zMuY0OnzE/YFFZrHNbgmxW8byPidlj4aDWBWavNoH27J5Pesuajes
jw+epyUC1eeUH2Jtkk9F/mphbYIruQCvn/9mHFFeJdlpAMZrwi6ZmLXm5hOif8YU
Xl5W2wJkh1K4nt381rplDQwprC1nSBRStkif8eAUr/SMmB60dPTw9+SmpOAuWYvN
eiogG2ZGk+Zfc5vGqE16ufgscHovgBOd7FPpVKRRXyYZKs+4yM1jboAF7z9RS2yo
bjK10EDcMngPMdOTbbufwZw07pwzbYOIKiDrnZbE84U5BZvYhONzXyDheRc0PX9T
KkBe8at7PMMO1UBFZXqt11wzGbh1GZujNlPZ0OJC5l5QN1y7LgivkIiPR8DZSXH1
ovNS7E1UKqR2lKJCIjvsvKUgl7esI33106EDDhMCG2uI+7USz57hd7f60uTjoLNs
1DOSlfUl3M1Y/mrBz1PijWsRV00y9xxOcoQ5do3JbFgE+NTrObmqoWS1GIEd2oNN
cgcqDSaYpfJXCj3d3d5f8EXuvwTyYwjEpATdk0TQIJhM5+w8TCRBncnEKVxtLazN
gE8SSbvuclFYUZwH0gLYNKuMWoyFm2LBdKd+xi/sPvtJgNCwDdU5YJBHFqIkLT8I
3uZg7nPKfFwjHwklC77Pad78zE4BqLNNU7XSFQZ0d194i+EgV8xr9YsSLgtT1vjS
OObNsaKcZ0awZN/9qCtldKF1bXmuKnLURsbc2Ben6hwhBdqFqeBI+Sj/azWBNAYF
TD3m3oEmqjZr7GFH7LN8lZ3WA29pas/NARFd1TREirxv5ii8kLMfOoiQCDA5zmMW
gfq5RPwlA1tYDhjbOA+/PYlJWodp1HO8lUK234oAZLHqXrz2iY/UmTmVtOqakVjO
aD4weq3dSOtUm5gEL5Cu+gisEtgmuYDL1VR4hnaCTbE3Mlxgl6bC4KK0QnwYWuhZ
vygDkHynYSo6c0IzmnDoc/AJN8qSMjueRZSSc66ilrrhxUPLMkcjeQZgQ+GgCJfZ
cRKCOLc1wAedjp79J/La2wLif2rPepZL6cLU91jq3sWaO+o+NrgSRu6JBMVxZ4Xg
DRirZkxthpA3hn7c4KB464EKxy2yT2h7/pPSzQ2zXS5FSn23qpqLsFpG93kdeMQS
T5D5+enP5tdjRN0XfYfG5IRtyyGRF/RSvXTNGGyZHZbYnkGImH2csXFvEtmigWo3
OlrPVtOOEOo6sLNyt/1XpU5mPnwxDstQmww+EAqMkF5an2/K+E2RvA5fH2GYvcx3
eRfJra+XaSZB/i2Dv2DkstKOHzHUZJjHaQoMABtQPPUkNHxmWvu89vaq7Q22i642
8a/Au4y8Bd9Fn8kYuznVXY4end41AWNlXNVlaEVEKd6N8l7VI+XxseOuYLAkWnPi
D6up4P7Ug6UFYEDjOVlw4NAoAFrNgk0j99d11crGB4pWLccZBp6syuq+juwGX+cW
Ikf4ZKmLRKuZsjv+bXeIOUpzhPi56vxAWRaQeTJgUkKF0Od2v+bhu6BbOhng3M1j
dLh//sALgEGMV3cX9hGlmOmHSmPP3DoHyxeeTPIpMLNEIQcU6t9x0DPGD+BeQYqp
N5l4deW351HbrMVS0Ikruq8+ZkSkTLvcN4w5+6d3fkQkVIqPhI3Xf9ttcR4Wpsmd
XNp1Hu3nhe6eXF6dEVHrcUfquL8tVG4vfWbUaRjq2v+HDBN1/wZYMvAdNOefNZ0I
l2Ap6vaKB2JdmA8c1NIl3fCDIi5Lq5Rcx19983Yn0yAnWmGgBi4JtMKLywPYT9kL
pRcw0e69st6NC3X/lHkOQdpVJ7E7Z2pTdZWhD7Q/UQ+M54ClzLYSbxdn/2AL1c0h
iSM/C+3BYsEqj+M2zPO57Rob5olXzn1KvHFwsPz9w0UwkHS33SHxEZU78dDNrByf
XNzpkfxpGu4CueOlY6cO0/zBYvqicGoe15YvB849xtRt/z+BVJy3PwfrhcmyK/jo
sjlAehzVhngvYvcOFbLqfI8ldYbcR9qkggp5SpbaidaXGY4QH9eNx4dm0V+DeGKT
jsOIv1R2d7zq1AU/E5p1hxdwEjGxohf4beLmqxDW7Wg92Y0thMOyhzFboU7GCPdi
BNm3CO4J9WUcThXw3YjitCiFBFonkce29OBW1rKx1D3nIw28G0LUH/igoOnKGO4L
YwOK78xhvbnsshXGLqTeEabAF8A4+aSxzjXrdjsXyWUN7TA9sobFXiShPXJyhNNh
oZe3awaQ0LMtXmxiHHNoFJ1wYcaJf6+QSoWH1uHZKupG1tmM4w+jq3Illjlbc1c7
UTxTzLuKJ3pPagKsGy/oizQSl/J0WrUc/W7/anZ/rY587Im2KmQBoq6Sw18b6474
q4jzBxQsWqFnQhbIOAmrOwW36c3FXjlqcDvEjqdj0HVKlpBvinq8436/ja/zGStM
HMEEI0oJagTgonkd9q/DRi34r1tDXTVitoe1uOqp4/WFw4WSWJRqVzcgNqx43FQ0
ueGzuJY+xo6Cmf+cxBVGoRw0iv7DROhfkqs/cnAwx5zncMTWv5ynjIv1Hj0WC8Vq
HjuFq6bBqfOO3Nj8nBfM0qYuM5haxv9Pj5qwyrBHNpxaDBFPY3cGGH9zEs7jZfPu
01sg9Di6KKnznD5539eXwugDM3tI9pPmEIyvRObVrwxJtcV5+l6nMptF1kqRjjRr
+F4ou6eUQHHHQo6xKVUmTOaD2TuBXMNgh2DXvUHyg8jsSqcqT3nKKRT7Yrf7AieQ
f+d8RP7xfATzvK/EGRBTwTaBBw+1UevgyS/b25ayKEyiJmObvy6J5hn6l+XtnxIh
saWsYGhjMqqyRV27LN/IxtRpheUx/us2FRGHmenOTp2wzbqLgud8NaSKosrzk/7r
dOzKr6aF7fMLgwDbgFVbLZLfrH2TjjmBYrB671Osewl8Rw7GUR1gSW/jksAfo4AO
2ei4SQhSA9DaF7aYNPfwatHn/SQ75i8f+3n31R4GIgXMVeV4Nu72EAnIVbe0XeI2
LnE1nx8AyvCLV9BbVcAsSVNlGVK0A50l4hNa2WEjU93a3JeXB7qTu+fV7ctjx2Vf
BMatZL6DsYyqjFhFr2BHV4BKwKAGIg0OWeiRbM0s6VNAm+aAJq5iV2JPZmSn2DBj
y9TX5GoZIQrHjmAKyFaKFyhCXflYzxUlt/CAugQjHpLSm1nx3oS6uVme8oAtCH4d
ZCpNlu4QTRgOsAIneNbkIY7RJh5CiPY8aX7ycdEqZJ8bIF4st1Tmk/Uo6OCs9vzY
d1l8n0s4DT1vSyXNLxc8xp6tFAHbhPLs6uNGTKFKC1lItNFlEq1j5OpstZDvH+EI
PwLssWxCK7e8bIclrMjtBxJmymXYPAituJvim+KcgI4mvSTu4GTxoAOXeNTdTpyB
Yo2lu4ykWPjj6h0OqL6gwERLPSTzAuZPrEP6KPXFNznVlY4nou1J6NoB3FgHd3wT
Oe4tDY9MA9DEVQpyiaV9AazYiDDlewtQa9ZDBZoSFpvDXGAsjFHCojAgnBOrwFNl
QYvg+peLaNtL/4SFA5rJNAWXuRgN+4DOvtBSLdNQE6sBnnw2Ge3bZl121WSNdnI/
klwrff1YM3fIiNmE+xawtpd9R6FuBxQKwWdmsaWFvOw2lYxImRLaokxCpPZCChiN
wWMJ0zmeNqfaPzRI+VdCe4MxGy7PoVVHZxuzP2919KbH77wT3d4s3FwVoJEDQnuo
PvxPa8NtaIm0aWyhYbaLV8o6rMUDnIFiYKzlIIuXwSc/tATGAi1k1LUDzE9y4izk
JcVmXZcYcdDpak1wUAK/TQS8Jn9XZO53CqCqXJo3SFxX5PuD5UG1rG1vMbkRJYMA
cFEzZYVKhft6+7gmXU2gJsXY9PRCA2Lr7dWlSqddiXrmdGGtLMu2k9wFAg7DtaJS
Lg1j6Ax7jG+JY4jefcZ7xOEXUchnfoPigz0t1pw78hcU8FhUjDDVs2zVkdsuJrp1
e7V5xMf0mQPD/H0dPOt1theraxJao3bZYYuAFLTqqBowfe1qwVLrsExq1k06jVit
arw+7oga9wyKduOaZB2DsBNS4aOhuX4oGjGUcks+uA1K2dpFpyxADSomBNuHHk94
mDi7tuS8yUEh0BlM9QfOVHfwp78vRHOxZhI7xt8bcWnpp1bbvyvVCzPGzfNZM8QB
esVhDNpJXtlM4c7VJ5TS/0foAVTDMByGuq4pdVYM7XvkdYX2RXMoa/LvDevqP4s3
lZdu4zC6pBpi8YICDSwypEO7oTynBbGTcEmu2bCnNPPNB7rcGIQh+uWX2MZlw7vo
5SJ4ffKOB/AjXDqXnoswt5gUxN8t5C4Cce3I+Foho3HoYVBzdVkChtA0SM8pXoCQ
mx1ZB7NuLU8ojkRpP2urpsPDCS2yf0axzSCxFtZA15WPP9nNHHlJEJPTpZjWrASg
Q8chNrtDVfnYGmmWSoNfFYMbUJg1BhEoxSsI4mWcgwVe5cpPlsk4iAX60KdDC1mD
EmbmlEeyUAUjeq0UjRLxf6Bw7nskMN49u/ukcMZDScbQVL14s8ZcygeFjg6awPBN
n/VbYg99Wzb/ykb5/ExO3PYNxSJZjOIjCytXvT12IiDcHODS81bAoKNQPizy4ICB
bO+kM+veQAGMpMMMu2l03L/bN+DKHGQ5XHeOqbkCqeUqql+ty5wD3IaC8uYN4NHY
7eoRzvXOwH1F4No+LnC0s8h2+HEBLHxtLVCKjapetJaQHM+uhlyEwTNpf2P/dwYK
P3AX8AqUbcTwmpE4D9u/Dycv6aPZvukDn+vvOpRu2ZkAoGzYzepUTkaac0UdhQKY
Zx4LkkDcAI5tFyT9rRFduJDU3YxF4UTBUGcCbjeUBtlo2k3uGWL8fuiJFCqL1HGB
7IRxUBeSsQcNOKfKR9NL5BlAU9UFIt4Rbhin3NzX713qYZel4ykM69j1EW0dqG7A
5My+pt1mW0B/5hnewNYYz9aXEHKdFh5iHeRrv1+94vlhGLS1dM9XoW0SA4PH4nkW
DSr/eOU4R14mWcXQAK7ZOD7MQwiik+enlvTtR6Ryoyex2TZZf8VD6iuJWE8ulNkQ
OsqILPGG2csec6UfGhINpH2SXvDR/eUPtxxr46yqJGxDH+8+O7HSf0+YFgT/OedJ
yk2wLUqm9F6wmu535wzYCd1O1c9lT2I3RVtu1QNGlSeok4v5uVIs5Zd0W7X0xItH
4pOtWqo/PJlTFBJKVdfsBnhQOTXfO/tsOoeTt1t78znGchidwkZALvAZiTYv2Csb
9pDzYh8Bcz68i4QDrplcF5sdYs+D0SqjYxQMoGP02ohbkxEGg8qSvCKYykc985wp
XCBmGGzczsKito5PGtvlprNiVJFsmCLDCppTRbczFfKuLn61uzHFpex4ODmbOGYJ
qEPZQ1Onb2u3+Rm0UHLzQysCB51dgxHU4BJC6ZlqHiKRE1ytInh7ymqaDUxlbsQh
/zKyceniki8OpWxGg1Az2fmaz1pxA+6k/ToIDH3GvQpKYXUyFwuRDRuuulC1oA58
08yFAeijJKqMCo/uZuds2vhY4K709MN0vyFKMkm8sj8I43jss5zEMddT032NKXx+
SCiI4VEibSSgLJj+xoOw8KBnP3HWsoZeJJXfwOhI5A/jRxv/4EBeMOC/RDHqyOGu
mcUpUmbkR4SAaPwQyoJA1BarywDMlDbCfTOhUIykL9u0pDflI72/B+s7Ky4myoeu
720oDfESIk7tSPuEIJNB1Luc4LVXfHCFTr3m33gdIAqxraeTAGB2NyaJvwOqcpre
2KmT6os6FTIDRixNkmTuAiZhLptXnO8XIgmYaurQKkyvE1WSw74f3/8SP4EqrrFg
SLVHN+5ZTWq9I1YcwrFkarvte2xb9h87mAHnt8YF/VPQNPY85ehFwhvOBBElkDH9
gtBmr3JKImHNDdZIwhEZdKd5CaDEGRhLHqGCUpzVGcUvOCDwEYGL8LvH0JMjPpWO
Zumj+ZFSOLHYntw6s4LhIdhSavApGyJVdE/sey/dYLTpOYSAxq2SXh86kfUiGd67
HGnUvBw+MqdWw3o/xbfLwTz+5f5hs7qHjexc2A9v4Tp5InJHul3S6uMG4UeeCZJ0
l/RftSgaXmNBrZ79ovtc0IesgOZsOqyONH0ATqgfTkHGUxrVsBBffx8WQV2fC0+j
69CwlIoaM2LvoppoH2E4WL4sR1uOyk46TQIU5RE06Ib6JEPIbQNe0QqSV4PZcmLG
StgTRiTVC29PWNF+QotkCK47Lfg1lRjJcdLGXNEv7JYQq7W3/mYnXIC3sCI0qcGQ
5xT3sWbMRZkK1Ysm98sYk3oZslZBLhFqfmEe6/uLsrxRDFcFtLDy/1QxITqN20nT
GDw5ANG8CDcEAfb/eG+OG6crp6iuSUtaVNuyzzwJBAlXqtY2tUVhj4ZwIp+WLaWu
6llX2wuIUFOOq8OPtVo7k5spS9gi+zjaoaTmsezhG6Eh6powWRv8nX5izmm4TvAw
xdvuXFkJzSSTOFkbyn+VN66DJoXYLL/QJtirAsdHHaj9EoQWdajzDIcfwzYX87Eg
PNSKYQr1fcXEAL/Oyi+zZduQch+kGWcjxEutq3JHxKE7YCyFVzCjKLm2yJ6gBrsX
nf/B+Kdcpu7NVROHN/ZKp2GkR1SGNyGqDcICb3OMU1sD93VkjW/ZMoM8tq86d3hn
ArXTc3JoC53kXAMaqhoLnVlJvzbVHb1c1x+HitO4V4LcRm8xPyyikwdUzF8hlYly
BYNJupbc1MwZKryH6n6IMmdA3drp/Kv0hhapW5Z9oqoF0oinkYqMvcK+ubVWfDFa
2SFf+7wdEb1tOQa34QOTbacTmD08CwQPBKbYlVMhzbYGv7aeBckzCYkUqAzPqLqA
yWTMR4sdatfaqgNGDDxCxY2dXbENK8nFYU02V84VX4fIb6ffLhKmozEFkFcN160n
Fq4dYeUhgs8y4RnuYmYmmTjyVIQfJXLm/XFQDRrWI0Y2knGS5bmTI7Kz4kYhGryA
6iXi6jeCgc5Z/Exdz+2O1BrAIRzjYoA2cSUFbV/qevzDF2RI1p2Mv+0a17E3GOE/
IZXXq4JFddo0DV4Du8+ZqOYa/lsTJuCwUxcw8qKpYZm3E8FNjKffGed791cb9z76
dibg67A4mfHD7rKz3aS9WRIUQdFaftTnB1yU63r5RKZAaSrCIkx5d5R3pyBO3s5x
tNFDUe1vbj5gtqlcsUYD2tQ4mwOQ/bK2rzd9PwqcG8ele3rcdID5kotyPoSd297f
vEFYuNmVnQkmBFFUQX09dSF7Lrncmb8SOV4RxGqOBUn5FSiuXgmHij1ZEYgqN7LA
FyWfHGatlXyTjBGBUVsiQcWVyHvIGqL+vTS570TOmGmXbo/9ejqw3nL3qpqzUzBa
/oS6nZA4oyCE34HQqTUuOlf7fCFhfwLUCxvV1x1rIN6pgSvl6vX5d42bd04wFOuz
MQuOVppMs/mY82oMU9VsOBYTmDUzf4Uznj0ydvCacJG+CENXA4fYrvavq5a8oWiS
hCNmU1NrotK4BetuK34mgJCo34ivN+MQCRpWVckFtAQqXRzXtbMGE/H7toOWY6hQ
vxsdqHjKo4ksz5qVHXu6+pzgojmZA+TCs6Pt31xlkjhsBbldebEWJInxhI7gAqKf
rGuJvDaKmHNT2O+sxrJ73FznEOhjDlkrKLRl5iM7CkEfSvMCejlieZpChFsRUHqk
Ko6y5IZFJmbYjTbbO6Wx/JSEKKWy3dwXsJemmejVW/tuHaZw8QemmgTFpTYno3X7
9ga11Yc3dHcgYh5Ui/yzG26yPYwn7bpphT0wL2q2H/OeD3CFVVV2MnR3xnQsySiD
+f5GV5nvXkuHpFL06haQW04J8gPd2U1MFHvb2iFkDyzC1T6B8fQt68/hn4gomC7A
OMjV61o03cZqxjPbOUpyT+QA/w83oBAnJDIBRdOS2aVqp2iRaFw917wXLaZAc2/L
vJ/iml5ojVVY/ReM7Y6SrumSZ/lbP8vUONWsO5x9ZozE9gqqJz3ZP6v7Y/0AYPz6
qqOTzaBoIgLQVKf2j0OdjXoeLHNeEy9/8JQeRusxJp1F2totCja5IYkFqIU8wXEq
F8tVu59zrdZXHLVqlzIlr1ITNv/X1XEUMevhc4mKP47J24oKohXnGnQyZ9rKIw+q
YxUIUSm1AT1VYzPJDU6TILMEyAxqyXwl+7/4XkvKRGAw9r583Jd6JSl2R5MTqV3h
VkE0Z8lHZrIIOQOWgMiEPLCEpFNmPJEkyV9lMuTcrRJF2cvNnFpS6lUUqlLC1CoD
vkKtfzArIAVHWftZq+fbs4BbrLlyzTj0jueHzPPiLyzFMYPRLrxEaiFZn+I9iB55
fsJ7CcAsM/CpFBimiiV5643SyNxSDOIzUYmN9GRRg6s8uxph0x9Pey2BFt/AbenQ
vOs8eHeSDE4+mOOhWeDgtU7Fn28sDS7wZBshnsAqVUVIn8AGRduYt1IL8pnUwNTn
uRblLUeUIG5Wbp1zIgkT1UEP5D0TlFcjO0lQ3YTYPgve5/g0GtITRCLNoZ+vrA8w
U/+/h9XDCpPX6O4yEnmVrRFLNSOjfhTHaT1BBLh82QScd4ysv5QFr/Modd6ixU3U
C7P+skC8NCWim9WxzMlAyBb+EQZxNDOLBgDIgqF4vNY+7Hq/5FTSO8hvu1/IhgzK
oGfAP3GqAPAvXlxe5huGkk75wX3kX7Bg5GUQLJfo2O9bGPpU0QaxalY/SWeHovVC
kb5YxnBUCOjVRrJoITGdf/bZtM29dG3F6vzajmBGVY5fdHI+G8w35+v0OsfjK26D
9SuXm/FxtsLx35gZ/04Uar6uQqMNGMO0pFiHmJG4wLeAWlrtV40TOBWEcTWK9LB4
ruyzXfqsYztlhXiH72zQ6CDY1rrA0zGw4l+zVSlk0LFmhOkOAFL9DOlhLAYcfRtq
nq5Iwqv2H8lo2t1DVXGVQjM3YXpTPeh2h8ZmYhh7aniGviCluC5jtriug8o+XZnT
wMisJZU7FL8QYqMC/wYBBtCh4391O8vMpo7LJE4afhWLVOVuAZKLqfGEdk9vlk9o
U60xTvClqyf9aEm90spBsQ0mq8PpbRLTg/fPDVCDUqmg3zdqReRF89O0DPz1IkJ9
AETPCzmMGQYv5T7b6GBTvmp6JPeN32f2/CoB7YCxIfSq4ZKVyxbuGfFLW6rW/dYk
+JlXtoymaYHV9hB2HPcBPPz3USE9PVVYVA5NbieucJsK393KgKdejRBFVCpOUgDj
qqIWYApPnczxJXgw9I/ADoz78Aol8fDXNFa/013LOIPg/9Dn3jZY4uGvNp0hpuiU
74S2OEx8HjkFf9yhaBlVoi/lo6YGzBEAAR+JBa4qytAFA/hmyqLD7gGvveT1Sx6C
VCLVceDre91j8fjsqkRfdjGlNPp8UcqoNmH/dQ3YzbrYWcBW8VLh+iuediv8IO57
mllWkry/pV5fY7Ol9XnwUHE8afIEjucY8tPFbUE/sjM3U70MjkfL24kYZxiOz8sg
jvxzH4qM5XcQT96jAOlTumYNR9Zll5s8vWycnozS2o2dCY/eahliE98oH8mFaDoG
htTDg496emqIvtv4mkzSDTJdXyP5ubuTxrTqkrwI3+gPWUq6K0ay8MtyJYhXdeH+
qT53rNO4yhDcq3tZwgSefs/RfEpA+5SdNP2z0kJHkbjHFSHp+uHD4xr2Slaq/bIK
lh2qw+pgFs0nI0j+bKkqQE23fbwPvGRbyKp15fOlidI7nTlpP9ABGEfWCAHCdwEN
CiOERKxe9h3cmSfJIJ09N4p55usSXglZm2R9uNeEaE/J/DVNXNRdvQRG32lyw1e3
aW9H5keGcXKPoq0if1+Jidq/LWGLbJ0JsHOVLmo9cBKf/xcwo+dth3WLgjalSHH3
Gld44+UH8nSwdayokHZgArKW21jiFGxXz7ny+0RJ7dOgktd59h4fQMgWu5UtRJfA
K5ip/jqu+ZzGzp+sm81hwIL61VCbv0pUxJcNwUB3kE0uC1zqAOWNipMcJLMY/43u
SZJZmZT6frKyiZ4J5bnamftEWG0YP97HoRan7++k6bDH5/szbbqnttixrm3CrCL2
yuEw9H3OvjRucn8cKMR9iHyEozRjNJOaH50p+v6IzTCVpqcvSiQE88uBw0MNKxTV
FziO9KlTxSzJlHxIlsXXA+LC9jEDOIfzZVEx9jEL1CGPDEa53PMdbi0YXcykH6gT
ZrEp423itLOmqhyyGQNyofoXsIogrGJ6CczliyStpeK8uUgCbYaGRu6XC0LSkYXc
rvsaCA7sChI92YT/lfbWasqbU78r38B5E3Z7DB+dgVk58fuWrfvpQAhN9PiEbTf0
m2f6xl3b74r6o5+mtTlRQRTBO7Jl9UxhJOvGHM9Pmt3+4vmW1UYcKatP90uLpXkc
nFHUiNPwYsqo+HucSFWHN/CFNCAe4uzlGunM0Xs6egO0HhtwNKgYHLvyVyzmhiiF
DjYX8os5GhHnyNnF3artOmPAYapzAyv54g5BiQYynB+I4M4NAKSI17UyYihiBAwO
EsgaknLqYzcdXKapZgz/gnk9ryZnfvfEfZIvY3hvgogR6Emz5+zqXejxXwKtkrn1
zuV4yA7AloxWD9LQW3o9om2klrMtxPoWw2fOcHLgbC9gjFHJwYtdoOhRCYWA5x+o
GnhX0pZ5gV9NnF22ahhzJDJe9KR0KwYLm2iiOQTwd01VqhZeQkNIQYqiBNq81oFj
Jlus7h7ilZBF7tcqu4b/QaMum7n8pSvoxp9XEh5Dyn3CkEjPxL6H1x/jRWzvAIBH
7nJHSz7lqdxU/A1eL/B0hiyYOv02Mm6AsOR12m5SYOC9k8S12h7vJfx5iIJq+QZj
`protect END_PROTECTED
