`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dW6ddK9loPzWF4vzcP8iBv5haERKJlqqGHwLNbPI2AHfFFvFtQrwNw6DOwaqx9Tm
wflGXLmrOlwbJoFeqKogUPs5kId3oQwxatUtDcdqN4+T/z27/G5T+9EGnUo2eDwo
2NyfktGarJg/FC9oLKREbF1m11I+wPl07EcW9wQ3hGT37Y3iZ1SA93hgwvQn3P+D
DWaRWNH+InyaHeaVgpp4gA3emwZ7X34zWzc42sE6CSDlBLtyh7o3aIR9oSGbhivR
ABrAaqvXyfkvXSOuL5LHC2lurPlM5ZMHiI0p4X5TdaEw0S3ZhoaWGfY2RLqVsc9j
PNhaASZMU/rmiKFwZ5b1QN7tLGEaMJwmXhfUHFuFNWSAFSh3wTlE5k9Lfgsm1M9m
mkYQw5idgYKgwRLlqhWovtRNMu1y4n94Ra2JSxxG2ZjSYateGMX+wSWwZovhmnkW
rau1BfdjwuksK64U5jnrVNX8pLRQr3IF65vzZI3jaBs4ze7+a85c5cUpfa4vK7zC
J35+2AvZ9nNiTpk7FPSoh77wQym4kIp2tMinIYDwdpc8aTTQR2zH3aMc6qL263R1
GRh+Ldl47h5716C8nIhhzQap76S3hJ7ZgVHxYZ3O03/5YlE5F0gHZSXmoGMpHTaP
tvTcF3mN/ztj8kJHwv/tUc+RoNDo5S3NVxSloc+APZdQ7sBQXtD85Zjst7iqTwfO
NpUnuE2gSXI2GtLwD1hvLfnsqBDyKs8Nt/PBLu4Eb3bzVf4UQEKSofqvHJwLQzVl
+uLc3q/FZfB46GVHtEPm+ouV0vsBksrUK/VWt++XKpWpCGBRh6OIzemmtFaXcBS3
tb/DSSI/3+/kPc/q8JOEN64+C8U65D/imiF+Ue1LSR+e5PtZZUKyqughGKb0QYRQ
ZYhCrZP3OjoLNrTEC/7xMl9Z717vNDqlYMatDPIwX7YnzWkdVmjUszwIalLxVbhH
OU02/enrcNnZAVeUfN3t1SXG33fb3sRop01xWvmc6ameznZZQgPTOeiqV0lklGoo
0XYU40d5CXgbIqpbwDviHpKg+G2Zn3zo6IRJtp/CooM7msjwgnMsTnq25Fxxs3/v
`protect END_PROTECTED
