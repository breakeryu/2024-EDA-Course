`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mA8vvyqxmiivhpkFVVB209wknC/E8ofzu786n6lX18+Y4g46S/XYqX9K/khAFc4g
g4n/Dkqh3kIkSYhm4fiWp3N7OaJ2NaeKqxCl508xk9Skea+ENQy4vNe12q9kFw/8
FZy0VPB6lL9cRZZgHe7WwXwO0HoUctMyW1C50LFD3b7iNVJUIwdmli6IVyFRTg63
GywbceCzHH+c6GoflgTI/hxOop/+qbwVjpzldfGtfqKU7XdPYukExzeodklsPnbu
tYmTFwOQrcWXC4Fn64okgKvHHEqL1aDTDBvXDBorNLFrswyV5gJtIjNIf1f1/F2D
LxcKdVeVAMYfCNkYgIleCshtDJSqrzjk4kh3LMSxufvlCvr/Sqfii20EhynmHssD
BAyvrpcti/sjZJd5SyRKjF3lKKd/wCaDmmKfLf4OJnunWd1mYCia+7BJuHLrI7TT
saSW8sPE9fkEQZo1WFkXlMjDT2MzuR5+jw/Aj/u0ySzbuxdFEqd51QPXeHfPbfbk
Ye9q1TGZWmSXbpaffF8lzEpKyFUAJEMj8r/yRqxIIbtguAfwxQB3BRprLw2O8pBk
XC7NGqHgezCu1VLbfbeaeXpuKCrN0DBeevg70E21GBH4Has2+iHGoAJKou/eVjAV
rcdsXs4D8JImw6nRRTa776WCJ6jqGuP78N02ZhFRVzYUvuHVfOEMnvSPO1Vnm06+
cWynkIQBfo1frwLtV+Y7duxgI87PbfHqo53Z4wmvcg8UesD9WBqzGMEj/k1p71NJ
WGgPBLD+WkIoFHLOsPmyhJk85drSHffrihdkGfMnAJpM+Y2BewG9p5ORM+kjoBjn
gWXzl8/aS+Zhr2C+/DfHLLRtvTtshz34SO6jkzBgyxy7AvYG1ex28ympa1TUtj3L
W81xKuH8CkmdqJsPZW7s1MfRSrlS5hHF3TYeeW6WU64iWF7N/YmEMff4LmNBG+83
b+c4hhPVpc/UEy1Q1Z+7SrvnP9hExTFKd21moe/Mgh23QcUYIsEp+3i0vOGKqYxl
vczPUref9vt7WUgNU4LLiZPomNsKIsC3Fkbg2YgH29PgZn+fQ0yCmTd0XyREuPnT
PfdRW5tJpRJqs6LQfDXbW30XUWMlbS0YWbCZc8DD1Lefu/KRvAVPLCfmAONJwXRM
e+fNvx+D8srZrag/y8cUtALasnqvjV5L8BQ+08lV5AoKcHE5O/P9zmh0CxCiNGjQ
cEQSRwkgbP4TK/IpBsBcuRkRANwNZkyDpDx/O25QqGZlJ4Jdwbd1/bx3aN1+DUml
iD0LFDPCrIQRrHCCOiKU44mMB33Eiui8NYZl2dJ//K46nYi+f8k31hDp8TG3Xttb
6Xo8XV7X9Y3k7CaQkqvIRDiBF2HJJMD5UBmCkzkP7DNLK/SkgMLN0zM8ij2/+kTl
ww4vOpikZx5SYOcm1CcuNUIKeRR4qE/YBb9ODX3WqKzowTMlpyzHTXkT+OQChjY9
kZhF5UXHQ3XF4gWBTkyGg4P5J+VN8rlYSOfTQtIKZ0M=
`protect END_PROTECTED
