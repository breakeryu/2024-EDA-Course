`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOflGpklg2oc3s0aySp1yfMfl9dR5PEufM57okFe0sBaN5bEJXwEauIRvGvGMgJT
OUqrMj7CWRCHkV6swxTjSDTj/3acWLSAbarUD48P+Cu2uMDBnCc7dBC3xzI+iIZz
/Ny9YHTRjmqAR6RmOuuUqEXRi9R6gcFb8AsDCtZPI9daJt7ZK/reHFe8ae7/at4E
gM4MdqscLa1pkmLsvUmecwrbL2bLTg2HZv9VCqL8GGOSUG3JdKy0hXx9+3RGO7Uw
XLSvDlOnxsunQkIfetqjvTmaq04Z9C4lq+6NPSAioD2v6QgwMxxtwYNAcp3SYofI
+Et8xuy/rbFTyWHfuceK8ciO91flVFN2LRlCIIVH4bqdsG3EaKr8eR7NgrB3FvpU
A1Bvi9dGZA8CrdJgZEr0Zng5v1sK+IRa8KXWuy/5Qk5c1//VffWtd2wsIVPNUFeR
QY+hnp+nPmXy4QJAwvWcXehaQ7gkwUR/N7LvYHrTpt5A1D/X4c+qbJziTVZwGR6r
Ap9qrnPgDftStmvP+COLMB8u5P3zk7WxOf81/eedkHyQumd5cm3QUpAi7PQDKafV
cAry5iBgXtY6ilQNFiB+pd4rzHHwKyBeCBXsi9XM6vmjpGsvhTmAXAAXyL8ZdkMA
Zvot6TCVys8fSmWa9xkYyeh6eGkwgGvNX/mRXGqqyl1OSeHKpMpyn4opay6zLdim
0ovwpCbj5Ejdbeb1oXYpAC9OwMGypIMcUm5/HtiCU7v1SpmazdCfdujQZWbCLMyR
Kx/hm5H1HlUY9h25RZPjdup1c/NVExjJDDzmKueCJ1MDffqM32nWQxjhm8SAfq1e
xzcs0KXObttnkVUIgAM1i8YGIekryiul8iVrf+RxwtkXTScnhks/hU6xG/hSPa81
Z8ZA1X7XJHVPxu58XrlzlRAHDp+b/9GqrsTnz6dfNN/bnVHyah2UHPTBvM6Nauxy
EGPD5iomEj+U4zw4ebXhYOwcBhA/PxUjCBAmXG86iJy02EIcGcRGSjRskF80nKYu
q5Zz6PLSKBsDJyiiy8V3FFFlXHns/4OD+JSoMroJ4BaqjCoG9GHAIDqiuqbrAnqz
dB/Gqs960Pd1X1HYw8KcWsEiGO8CC7P/zQ5Ic7Wrc9xAn+wRiTD5fCFoa2stbJpW
Zd47grEzPix+M6ZLPKBBErMwgYAhiIbO2mr6gOLzOUPXNHjrRxJygf6zRNSV3qNG
d+0LsjAPPGVWRylEUWIuyBKzH3kLfNvACT5N/CR3y/nTTxROH3UQGlBQxQgrf9vu
JdwQA9Fm4xlJcZWopzpyD0uSFW8cKiU4+F6OaPAuBJr83ICj19E9mML+BB6EyCk9
leMRJGr9AFhwsxtbIYRiLj1QRtiOSxvPi4MGgq3qx7zqCo/qbiDbIqxVPIv/GpCd
smPnZ+YBzN113EoBN2kbyDNPPzueNSjl1lzyJ2cvOVaQY+IGWdVZodrWYiHjLFvg
RV5B/BEAasZXca/O0Jiph8R1ndJNVmV7InfZu5LfIf3IUCyU9CsiZKUBv9BlHWov
oMERsbqtcqGV+EkBKJQsPtQUuxHR8La7kPPLVndfjc8=
`protect END_PROTECTED
