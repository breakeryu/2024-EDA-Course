`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QSez7G//YeF+7oTcR/GhNySW/rfM8OtVfuVXed5qgjqI84sztFRN+zV+5z9wAGln
ZF1Q/RjVdpFcojPDrmwgLLjAyR5kXum/3arjKfJHv9mIHi4rlDbjnn0vveWfdPBn
RBigLshvL3UBt0EXOJ+vQUgVniarwIsgR2n/W04HZezg+Xmm+BtrtaHXSEENulq2
55/DVbQRSKmc9y0uKgv87SGlG4Hb36lAp4b2xbywltYc5UpVPnRsW/SGCZoYgDXj
/oHvmhe7I9RIGasaLpV4RqhHBJB0g89G6sYAj/YPvcHdA5yfH18X+LWg4eLc8u0q
xY/ZIad3fKGYNW8hKx+IkQpcLgLTKsO69x5sM1VCcNxC4HTI7wFiQJjwhv39miJE
iSjwZVfhn1iyN3eSFDIbwgL7mVwDcgYQROqtS0O0h2AhP+72kXk79Qure86TkrRh
Y/nIbiCFI5fcarUgRXNpGy0zRivNHCgAoCVN2JviPAvntsarZ7mDan8NIIiy+QRd
hgNXx57rVMmEq15muRKhCTUVbuKwI4Bs1LOaorIBHlUa5YqHzY24s4TF7GQghZnp
PQZdkwavyL1Ep0wljy1BfbmQaiL5wAaCWKRnNX2WKjc++qW4/yGBJpV5n8zrgmgy
2GnFkppRXMUPfR0sFArBD0wJ1VpjVqPgbnDdGfz5Pvf5nSSMlgkdrgdnU6vQbaPq
x7G5juxUQjqkU2fFpTkvF9uHUxy/ATuMe9xLZInsmK4gtIqO7YqB9tzipuBr99l3
9QN4I73B7bu3NSn9KW9O7Mdov4YriCf1TxL2ikFtv7wET3kWBSQGlzYD3KbgnZTG
3jJxlLytewc/ETcIh3MB180JdwgHpvAeK2iNxSqh74NiUyzmBXixx1hc1Ab44I7b
eSDoAUyDSbkOPE6AwP0Rs7NORnbAXvNFLMbRxJCMqOtjyzpTBxHtQkO113YLbvp4
fEhJw7fIAOmYl5q3cPIg3j+1mVtNk5v+mvTYWL4edHvnsCodtzBZvJGLU2rPS//4
+4KcJ7aTJBkTXpzVfL9fcnYqW/7uotJN13vFkyncOr6ko//VBoxcpueMGTlykxfi
x58KAdROIGE01Vt7PByEcuh/UgS7sAq6F2V8IDsFIZN+YyCxg3HxQBo7CiU/PbPd
ObDN3v9KtZBseM7O3eEgaZBXoNhkv4LIcA4lcmShf58uPp7Rzy5kYPv3wo+OJf6I
dtwI/4O+AjKgweUx4yumz6yGwO4PmbV6eCFI+6HZUTbSef9ce6UhIu2F8/b/gedM
zGWTzxg0pg1gTBsdHBLmRz/UwOxi3NcHP5JZbfYSm92/Y62ezTDv4qk+qPWRrjRv
c11L+sVOR6F1ayhFCoVzJV2tC8bkxD8qQW98Io18HmEeM2FrIlTx9GfxhUKpWpSc
/31urpf0HA3aUFkqXPQHS6c4BX1HKZYuus55abIS2oJczOu9x5f8PXyDIMV1q7TA
9A1ArYZ0Wl+T24++ki6mjSkGkXogW5FahPwr1akVX7PZlOwkQ3fa7feNlEVm5YaF
jbwocSKSByrCG5zrFfNVLMovHk+wVYnky5uhw8MhsdDgIR5/Gy4YqE6+Ak050OVp
D7loRSev50jFVb+gnhb9/zrTGr8kkdLTYZet+yaL6B7+SJsHTZ3PpeKVAdjiC6PO
2yi093i8qEqqn1rns0ePJYnvT8JC1XAolXzjBQl/erBU2q0T1lROpPR4G3COBLob
sBG1z6F+oLoqck+qY8+v0FL04cMvAf6sOBNSJ8FaJTo1GCUVENGqINpd7eFOp1nN
aT9x263msTsAWSifF0Q3F4OqHHfFc/+mDVztQ+zBdLKZZ8GmMclqXKXHfGYJ7yJb
ghLSTJo/ErUD3stgr6qShjQ5V+6rDzWq5hQdjxhurOn6m4JMZO0PxwV+7qw1KE9c
2EmHeYkoibRFbbSN2RfapVKmdB/TNTLtLGpNiwE5N9mtgjRd7HpqRl8qltZFiLGT
3NtxhFJwdSlk/IwEUOAan/dconD/YLovz6rNT2cKHvaRiNiXSCqQGl4dNPsrS/rV
P8nOzBVg6n8OZSapEkDQvwSLk+a10+XV1DHRJYgospt1BqKPBf04cI2JaRaPYJzN
Stgbi1pltCH4MqIFRSQ+xiwNhyv6C+gxt7QVdTxD2yTmzO30yhedkJyAU6IF4uHg
Qlt4chUgLw/J9bIqblSepbzKOv8dXR+gUN/2WcehV2jHBxBoa8oXJC0dszuOACkr
E5NNsZDAIzeKxMx11mIDOoUeQcm/imTMEXUxKdncWxmKL6P9t3HIQSpjIC/bZNSK
ykj6xmC0hTLylMdocUMFOREpLzUno2xvpsyL9RyGEy0e5l9fYGUJPa4F51xGLqUE
WJ3lpNnwaRNPThF0GIP5SZMr+EkKuQ3rcHMzZN+XT9K9N6uWQdo69zTBKhOtERf5
LkDcZOzpThS3a2FKr2KT7HQGUR7yWkn6P3D/yHpgDqjF9EKonWUvAWSr0Et73fYf
JlPxmqMoxAufeSVMAmx7+oq8z2m44eovbx4Bt9fA7sFfcPzyKNEBQRZkqSIrHI5Q
gUFUmTd434JB9v1VDI/c8JN6vfm/68kaC9xAK/BEeEyY3XboVsv28P5gFn46qZ/0
YeogQEAKM50zEvenJu6V+PLSo9s5/crJkU+4uVgujg1ute8J0X/FNOUMjAhPWBSp
SQ6cmBas/2VFC4ZOvwF85Z6o3MJrGxQJXrKb/8lqYHGe1eTtriNZi82cZtPhxX/c
VDxNL1vxUSQ4dKDz8z0PNxZj3lPcBr8t0Z8CmcSIi37ocAe4C4yi2X8vYqbJ4qdg
SumpeZNU1o/HLwoL2tGxUPDvMSL8L7i2/IHUuqB6QB0vAr7YU9NuwxEm0MjCSnNZ
h6PZ02pbolXnEIkJkMGboeNiANuBTMu2TqxZq4sSMW/pcOXfIDJwvL5GQOba9QPU
rWOcdLUESdfx/XnsUowA9si34eLpjbXMxHrlAavR7Jv8NSYh779irbql1N7Qthoa
9nLxawzf//aJhgmd+PENvP88D+nC3E0MBDtdCCOmbkNg65NKoRexRWVFiRUjo/nT
lPYHb26m/jy+rxUSdstwdmjxnZqHpKWF4hVtlsKBXs/72ecSbwKE4XeP/nz7OAxi
PFLvEPTryVukhgtUPcZmhteJ8LdAx38czg/yKrNUcY5EOSM1opFv9aiMBRSgjbbe
MmNdV7Cyl6T5oDaqesoylHZ3eER3ltPTpqW/5Q55vleCJmQd2XM5d4yRhstVwRTQ
QTUnGCdsLJtFRTriGaQgrW6yNgX9kCY14ZSNbXA2zbswj0FxcitcPthaneupWUIW
yUfwVnw7zIwcTxerp9u8yGb5fK4ybOcoh4H4F0rJdFkanHdQePzF3TXW2w1JpIZ6
VMKnwUQYXgn6+BtfK6xsh9Hi9XMmb4wyHGiHKFeZvwyyNxabypTraVAYRX/wy1YX
RwlosNUn/VoKp5JQ229RDWmMQxgz39LZX4E9ASRBWMgOTiE/3Tc2Qh44Zm10WqmG
/KrYGEsmqHFr4XhKCSXLhqdvFMJFu/GB3bN8Z4Pn1U3Ss5R1MiJzBfaIpoiR5cyE
FauwWQdsEH7PYRAD6L7j+qbD9lmbfx5lxJF6k0QdjEhs+w/uZ0lfQqOyErak1O/o
kAja4u88TZnexMzs7EJlFlxsFpkISEZXYVdD2MZQZCkqkb9nWOCWp8X8E7FyoVnI
YI1Fus+0UTtEZ+Itq39hU+f0Th9JPgqBuooYcw7EnV7WYBibj4JYzjxrN9rpUZAD
0kGhIR6p+fuWGYsnLS1JEreeKNqtzxlyua8dLGknmwqA8biuYrDvvLhNkSnSaQsm
JcxLs+7XnNexOlt1FyembkDWOqRz3CxK0uBGMr4icm8y57jUv/78UCwLcOCor2vN
hTx6mm4NyfJNx0eeN0AB+9yHdSYljmpkT7AAvnZ/ll4VtmBy9AGRULE02Ea3RO8T
tCw9jvHn/yUnaH/8Fk/tPPndIjKkUKYasAc6XjZMKuM0Huj1GjSFBCqLVL+BI+V/
TyjQfMWSrbtnoDVAorTXSS+xjLgY/F0pkydGvqWDb736M/D+JnxnukcXBjpU9FHx
fMraTP4rj2iJ5btbjQKvO/j+om1gRQ1WNCk9aMTYaziRCA4CKB90lUh69cps7yda
ltcuvQju4LsT8WscEkM4DCx//hNGFjAb4vw44AUIrCAphqzG297Y+EQ1lSLf8vsE
IOw44ymoLwCohGaB+tDAG+8XpGGBFj+IlErChYWr03Vu4HI2gVvC7RGApNCzkzsX
Ki7/xFWg/tND91hjXI3zLQnX8kZdshwK+HyDtWZbUcAzcD4Aps89s5rg3RvkiH0o
bA5ljSUq1HeVBRfGt9EdI9c7JUh6r7tqtz0p9/lOBqM9I4z8Y6cK787VGOU/1jF4
jH9us2PgRfCJzmfj6kycOQtTN0JOWWBbML3uXwqB296ntxt3khxPJc6ppXnQ3FQV
+rTfaXmsBUmd40TRwsgTiQ2z2ymecnG28FcBg1wDgt5ocZ57SThv+1sqhzqNcEw8
B7n98/jDuEYh6LidAEY2uzp6jczyoyFeVe1vsgKCCrCGJAR3vbKqZNyoyKyx44Tt
pgnVsKHuiMmaaSZrpxchNcU/UPik4j8FywOB7BKejpfs43FTAcrRYJP3FxUbOuAb
ECjEzMhhS5Hiam2glduh2LVwSyuvAW9sdxPMvV09NZpk9RPk1cKeASSazcKP/z+C
aX843rH5fyS8rzs3hM5AgUoJl2+TN+9Pli6QaKlNruTSLAxlsgNfCgWDt5ksgC28
nSrOS+L4mv90yyHC/wLEiiGwrwD6KrTxqH/+1y6tSDW3Z++V36NWfEDZpMnlJDVK
/RtlNIklK4MeFZV+kiqmvhfjFIDNHqBuO/xNoAmStK/qcIN6mTdaaHBMmamll4kn
cKEBbx25KWWsCSZBOXt9gVW66W1w+26CUtKJFbzx7FkylTCsGO6KgTy3kGx5fdiA
VBMwItG+Pfvj/Z60rZ6JNvXxK0GASv2GnhMZTMhdgqG4vBYtM7WOQlJtFI42AIZA
diq6o+YhTM/B9dtnq2XK3Tlq6FWZPBFoEQ5ks3XqScvt8vCQ/9lT0UNyZmn99Myl
ehtWNhgAZtomWljDdORqrXAkG2Lg5rFZCHtrLdb4O49aiZ/YLNmf2TkwyyBIo2fe
unpDKLviLy6mJTTeOt9Vz2blEbfe3HM+imrMOfawZx/pKkJHNi+5WMPIauInbDCU
wqPBtNfN8UPLHVaERf9/SLvSTmBtGSlRnZau+5dy7BubBBQzcY6rdSsDVwiZddDl
NrPVtpZ0BBqMyQ22qXqFE1tQvHl+wTJ0VYT4xRfgjQIyLjdSMSR7r3ggL0XI60rT
sMLdI/g2lWxnltu8nGLl3nnGZClQ8ZHecnVeakKnNUOkBnsDQRMspf3TcZ7nOOkf
lAtLF6m8RoGtYpiTMflTrVNlOAUQe+WmQcukFiumSjXkuJJOBm584S8ajPssrEiQ
tI+tgB7TxZb2G7zIeXXADdiaHvZWGMvnsDea11Zb5DvzNt1OJ11ngERCIAGEhwVi
nIa24bd00wKrfUpgzkd4cO4rmnnCusY7Cx9pqJKa1sVKIbRy/j0syqpJaXHcgc4V
EvEn8mb8qYWKXjAYUlF4Lw==
`protect END_PROTECTED
