`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yUmInCQWsyhhBOlyZjLocZJDS5d+hENHdAqjkjYbH8Nws4DX2s1v0npbR1x/Q4cX
0WyAbThD/K6a9/M5dUkba+odx5ize16xUsC71NMAPWXnSRisBZYEq/adCBsJPYj0
Gsp+fqAzK/2FtTxKBZ2IsJqLfRiImBtvAje3YwD9HekrUteGCYO1ZxqhRF+CoGsj
VwqTgonictv3V2zBBSX8k2pvtQC6HizFYbr45SK9fYmLBHPNvhsXfItb6Dw5N0LM
sbWxYHdXY3RK6SyMuw3q09hmaAbMLOheLrslXJtcrNt//r18Jsf+75+kWOqJbCAa
VtxsP/bTJVcsZqkGuagj6ExkQJcEZZzyWvT7q3W/arKvTKm5sEbV5ljm4PGXWa4O
RZkv9cOdPml5v5NPJD6xmObOnCv2KmPyZZxRFiOUPL60rS/qOftXqfjML+c4YG68
18Womyhh1LW2ewzt/bnKb1yZxAovNKRGElnY/WT+ZhC2Eyx6A7BkyBJJQBJo2Y2o
33vsgdAADwoHrfs8Effli3qSo6/iCS/qkKEJrHSyDxHQsifR1LsVL3HMGTCsVZou
msQhC4VXfgEK7/VAXlZRfuv2xiRcKUVRe2iRtVNqLf0asdziSJR94VPLxAVtInlH
RPVx6N3ogUY8XArEVLFdmmGdXP5TT8o+slVDrBYCcWqsNGco45cyM1T41YIZJUmL
lMz5lWo8aW/MmooBwSiZypmHcyJVCcDwQtjyyLZlXYqaFx7TvAY8/yg33L8jaFTh
tyVH/6nLI0oeb6vNs4hsUUjAGaos/BydAE5cusm8Ti0cBt9tvzSXGwwBvDTM76ep
mn+dxwPjKy6GWk3P34kkc4jvvjOwuzcNywMdXyN/2lQtx5k4R0jZvD9niSABgwXo
vtL1Mn2K07z82k2Dm+f2mOYdPUghOHlldX+qJZL3T0c5YWo7VWJhp42XNWw8UdV2
iuHS5YUHxhVfeNeqTELcbCl7YPh2+qdYpYq17Vuo9RZXas/+R+J2tVsOd1uywDty
kwONBcn3cH0IzfbLVsLRevMSH5r0M4iJtZIwy5YMVMSQhXTs02yS4MGgRVhdVm4x
ljDZUoaj78jf57IlZxiAllD7sFs4Xo+szTL2GkZdnx5bK62vWjBfZuErgCe+keOu
jjiI+Kjts7fvcM59OakghoaQHVMZD8YoeiCqO4dkMqaJ7R4NskEmqYP1VntJSjRb
X1ZQPLXsPBE8j0GybIlern9W9wrNPi4vAkXowPQ+6r+Jeu5gWivxpe/qxCcF5EH4
32Y+FHXdmPLn0tVozYwFioa+8jMIAU9Wr3GPbDcU+vgJ0HDPu+Gj8RJ+CWV4VnTg
izoqshsa5JKYlZKhgV/6IkHoY+/Xfxv00KBPoMyfO9uIRTM7LTJk8MJNPR82etST
6m9s4OlmtgVKD0Gn9+yGXrDX1NCcmuikXJWNhSOwhrxjBgWs98dQO8gJfipryqLw
LKRp4ZaOdC+tbR2BicoxFn+lS8F+LB/0IlsxItmrJ55z+Gz2zJpobHaNDVUcVElf
AKZtQ8jN2bjNp7uZfiLQBZGzZ6jghrh+Uhn+YmdXQHoxcKgoojYVFVFf7VJK5HWm
ICcH1Cnf/JTB18Wa+at2UknIVZk57vUL8lnqNsdr/btDGwsPEUd3MMG6Y7ZZxmpD
jySAEp5Urg2YL5g/9oGbyHSNRpqMw1rnotbARfGrzSoYQEZmC52qvpttvualoCKX
I4hap7uGaLAlSuSDfWVFRBHcg2pleu49qhfV/QlzkeZo9wwJkGnC98KfIdualTbx
sJx1R28Kh7q5mtZNEPXwRcsdoIzCKLuQ5Ui+c8grJ5aH8RWZSFfcVQZK39+CuopR
kpa2FSx/tEAhIDTrjoFT4nO07iGYLog9t39K89u5+jvFZvTUZ+c4N0pCdpR9GiV6
dBhFhuE98vqH5pVI49bKqKFvEWDRv8dSzSowV3hrZFJ7AyG3wRGN9lh1OvQ9IMrh
uXGhGOKom9gl+ENfNGAg62/2AOvwo32ooOJhA25RwE8Dq9CxLZLfY9g8Kz59lOFH
h2j7IV5vHzFWi7V8BSVFOq9rw7DQJmtJInWi3CxktfnsS711imtC+eppKO7lTpDO
EmkSDvuRpBopBvvm+YixTbHbajCYhtDz8dB3UKi5fuksHeWZYgPaSfsXiy6qLhGX
8L/t4p9C78azr4ODZLTRDOT97EKSwm7iRf2SmJ9F4yfhiEThcC2iQUFkdQe/eZR3
ixGLV7HNuhq4ZvxrmTK2TmfuFeGeV0awrTnNiy6Lgm1o+OLjnfLkXo90Lpow6hd7
NXsIPhTBPi0qXtHs0ezIX+jj5D09lASG3IytPph9tTrrq+wazbE74zx+MVYLsQ85
FYLO1HKLleJPD4Q3Vd7lNw==
`protect END_PROTECTED
