`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjO7xesLdOfXdFXudO5F1Tkbguyt8EP66APDxdFgb6R8i7tgYPXP/MjiHmoHJDU2
xTJRFtummKE3lyZnxdsg03sit3yB4LOBLehK1eSZqFgu8GjTyKjq4CnNAUf0uWE2
4qnvBvjvB2oLrpUonD4ZI+6aMUIfcRnGZXE9r1niDkKeU9GHxPNjX4wwVF/D/kdG
RH5Mxz7ca6yWiYgA9VL5lT+WfYdlR2TXHiHAqkTn4sNBXHuN2ES9KvdCXq1waIzv
6ijPqnAuyHv3NIGqsp4nF7J6I5CY1sqGrN4i25yQhDSAO/SSlVEtdyR6/sITmhex
xMX8PONBk4Ee4Pnw1kv2pJkn+Lr1Tar6bnkJQENoxUMbg50hiXHEL06tE+m4CdQk
85opHCVoeWVlkTD3niwjwPp6tMrp+HOiL5vSwFlT8zG513+PDpQl3s1gy21IRSNv
XAcw3bB8z33gsrBe6x/375W1whPlx/1zVghSj0zjaDDAXG6Ty6Kp3M8cAtDGB2Fc
9S0xPcB7opimtWObFpuduPm5YQiuYqSiFXPAPCv9jWi2Bywl5X0aeqBhm0rwGmIG
rFxSUAJPVGjV+xzBEdnJRhY08+LJ6sqC4z033rEjlMlnA25U3ZtIizI9pLEdLVUa
Q8DGUAIk//a4CDjNdiYQH/tJSEjkQahszSyHXZJNh2JZqEAb8Q+c35cmLKdNPLw9
1UOqmIuyyhtX/PddLoJ7rQVhti5zzQNiL+BZbvV7lngF8UPJHuCmnwKNQxFmgmtQ
aCiNzq0Az45rq2RWyrrIi6DJQilFnHVhbpl6XETZJKmfhO7Xo6c/2bH7l8SfI/nk
GeqHgo7qp5mFW+OzFeLDZOEjnLcIuSFQSNtSQMSSdyqHJP+AhGc8PqmjGHGrUIO6
jXlOuOPuFLCY1i7oY4S8Mk2DNw1VQ1tEfxugX4HoXNKQc6rOKAr54CHO41beSJL9
AmdhTCZfFHZjgmTfDCKwofUFyQWj39BP2fH3WMhgz75ZWpqJ0MKAySV6U4ajGizh
6koDazAITtIOj2Lxgwd2ZzInP5V66JWi+bqXGBJS8sYQiCYdw07WZxzIWyJSFRQj
z506UY27YWB0vIso/EzX3p0r7g7rYVFoiZbf4b/r9F09fExi83FeM6Q9I1QHSNLX
Q/76K5mzEgQHhl58GoNpzVQoPmB5ss/4h2HDh+WFd5Y9+W+2gvebNnTn04odt6Gk
7C6RLY5yt4PbWvbPXwQmLkoOPNbwe6DMA1Fi7U7l1ySalzHmKEOH3T9RR7ckvh1d
ztrpz3C0H4V+X7r6JdsmcDTefRoepFFHRmpcxPMuoHiYi9zblHoE4ww3C1+No6Zv
ll3CT1AwtqYK497BXEyopU6G6+yolJoRhpLnMa7SJpDcLqWQax9byjullTIQvjFn
tpYnHHgKQhSTvBaVC4K35cOrfQIR3UlrTNcvFGVK/dYcyXezKjUVrZ4jiA7yi2qZ
Vr0UxMbQ043b1todskG0Ta+hJoyVZypNGgn0C6+wnhRrevSzh+vdeKRMKD7uvlwl
nMGPD67X/nXfBEre5mi6Mx0L/u6Sh24banlBFNPgR8/YHJA+i1Aj5LJGIX+Mbowr
ss+1DNG66adQaT+UdJRpumk7vAq8SBg5eHi1GQX9D1xvx1ZcRoSGKzt2LC6mKzld
5R5eoKZNEWn2v+H19NlBdOZjqL9iFh5c4xhH1/3LJPzewsHbTY1Lj4QWxbrC5K7O
w8aVDNybvq91V60+KP3dVc4e4JN1sQKA7W15VDvRqM4QgWzM1pd4xn3s+jZdrcFp
R9XV9eOyEgM2mdTMeDHHOlkLi4H9YIyMZ+LxAffbWlPB1diWZaPyLfrcbDRlFlCj
b4Jpyz/4HnV4mce8VsqOTxHm7KHdTWI4fazGdhWsyFCdArNniiLzWiwcNESw2CMV
CynMJ4usIZx5ekItd7CPEwD6xz1wengYMdZ97Oi3l8crZGkW09amtbmXfQOuNfhZ
c9RrJXkehU4e+SCiXMuTrXSxnaEe0EJDMbsjtmtzRPjzv9vU9VssRdaVVrf4X6Ko
eIjknXebdzrj7owFu04Ob79TWLNsm8Dm3e9WJTaR02zPf0PDgolJfM/7Q6vrc3NE
H5n079YjfVxn3R99A/I7hlEyBFP4wtcIO6x/AxBSAf0kyoWWV0f+AGgJqvVJTuDr
zLmVCeRw4h8H2kL9N+quyEdcevwJumb9HbG9hMd8HErn9AEBdZGBlJO8hKHRrqT7
OSvQOzrDQQXxCqXqHwSh0VIKWDlc9ZRd8XmcXPEYVk105S1t0u/Td8KfOF1pGeOg
AlHPJJsT4llpSWElfHWhoKlnCqsv6HuT0JqSu7TmhFhKvIQB34NMuM1gta9ozh0M
wQwiVQhM2oExlvJb+ayp3CftpIzUaSMk09j7um7CdFBMRt9Ho/xkeMBH6No+rKgH
ou0VE9BjbrTDNm05HbFywVb1bG0jAcn4MdVH1+jknDYOZWtp4/jvojlyaXk9IIWi
BrhZKTt8eqTlPA5xPQ0msaYPAHUyiQzbdg/v/KIeodHSeWhQFnScI46AABZnQROs
zACE2So2noQtWHVbPhQWKnnpHccxr7G0w0l+RXAnY57TcEagbltX7NK1IWUhoo3q
KtnYq/txCCTY3gV/xFn/5qaEse6QbzeVj6d+6dQZmsw6JTMwe6uAUei1WKBJH7Je
hWxJwbmW5fX4pgZVyCbeRUVwF8t7boAIY7JVC0nds5tnUEDJ9RsiSMKQ+dpCjr2m
vX6rO/sl4r9c7kMqWz8+dCoGrRgZ2BGuPz5A+gWjCF5co/VBLZWknls4q9ugOe+/
OsEMqUPtOfZb1nO4Ht6tjX0cRp8tnDg2JOiiNjV4jnLt+n41XpU/l4wdEGoTNiRa
MmzcPomBNEzOEtEn+GyyiXSa2Fm4ki4iAjVcRKmvRoVc635h4QSBsa35UECdEFnG
k97IV+8y7CA6kWm3T8iUBlIMFcUDIEeLd2WGKUlWt/KMSh+ms6uL/6baG1mX+XAP
Si4j+HDDnGwAmlBBEGaTSNI9LHe8nnHOpy/UmwN0R6qkv/jXDoZlL1ZDTYwGuEqv
Fe9ymeIS6kw/1Ztq6j+pGna2n+wRXVohFCMiXcKEePhe31lxIDX/JxS7lu77k+ZV
hoCpfFEZmK0xbNoJFhvcNMhrJE86OMyHrn7maesIWYwjIPOc5kz8vtau01LvfhyM
z6Wpgh4DuoziAy4GOw6uMMOYMquKTtyRFtiGYMqvVeti2aozIlmJTYcgwg7KylLL
yDvxJfXmy9hysN2I6GkHatUMO35FQK4CHeXlbkpqavhaCUE4fu2tBMyQ6kKxTs88
vk7j7+ex+P/YxEAFBdwv+DoLwjvq7S8JLF2faw8bwFwoC925HF4yzTYgUeKecKgB
wJUzfc2GxAMvuQJDbUF8nc/DmpLr7jfivtvL7aPSorpwLp4JF3KLEJhgtpXwim+M
AsvyjI4XaMutK6zHUEjHXqlwhGIvr4TdXigCxvXbHBlR/xuYesRJJ3Bu6dnuV1Il
BMlJfcDBnzq0aGfgaCE1w2zimJ0dXz5eKzvjUx+VAEIaT/vMY9vhAOZTKmfSKnxg
pmWvbr01vLuBvBu5vIBMaosHboCys/XdZmmmEhQSuIoOB/o3sDpzOO8FC+aAPGcv
eDXJtfD9AMTrPJ4VTKCj5IjFurFepp7uThNQK56s3c6iZaHKyLWJwPn6Ja2eWSvQ
8LGC3NTxYznC00rU6AHvVB+xQR1NWEcQZw94gCaxQaU0XKz/swUs4Sj2t58gQ1g6
sQOwpOq6/KWR2GT30UUQ5I2YWkUVSjY1DcBWhKQP8NnzP07Kc4SBhklD4jTZ8KI7
YQBCX3Lpv6w+ixHS/h0gZtSltVH87auhpQ01AFX+nsQEYm9W7eGKn1X+q1OQPMqB
6EXNdHTElNcaTCsN/aIL1+kk2TwTUFIJNP1exRuXAm6zYVD7026FW6NsE3yKhHjI
B8VvOrvKQX3V/knZkY50azYNL2eK33WE7jMgzZfL3zYUV0nNOqGE0Iq48HjUZCs6
/SLhGyiiHLN+9JD63Lrl/jU8Z3nqY3JSZwBGCXpwny689tlzb57T0cBaTGMIYuwU
hS93V/J8NHVf0zUgVZxvTJ22ZV2zZ+z+bVA8JFZCZos1nV5DbId06l+0M+QaJhZu
IFhU/fXOvR6mV4LnlbkbXhy0hZwCEnBMpStlhgFyJyJIm75SBHENEVC8uIKw/08z
k3etctYBoiZNkb9xGKt7VIUCoZ8s4tjE+oXTYg4yr2uf0iYrI3E5vOzn8uSk7Mym
AGAten32S2S4z+9YL8RYVZgrrQ1kk1r/+vBSQE8sWydthF/Acm4rDV4aeAb++B9I
06iPU7NJSTJv4m9GS9LbOCgWer9sL0WxNddl+VtTC6LwPbwxk9cb9zVY3mUnZG3b
7YBijRn6OvGxkU70mxlrvUHkhfrITnMDy7Hr8Vx2GTEjG43JAfv8nqcICfvyJ6Fz
cN7gWAdnMIKYMVpEo97nrSDFlpqtVi0aeAk4psYJVfZNY1QCAmfdGkEnH5KqtmD2
mH09D4XjZ7h347i5YTihSaoJIEWbLqaWZiE6EDPN7v2t5GDF5u6OYfxtuP0ZcWcJ
P8xCmK6R2qtoI+8uI150t66WgghsvBgaChGmu1vSfVSyQK6HuwuhhHISdN9Cn1Ts
fetXglOL9FVBA46CTRx14ZC4VNkJngvtxIDC4zmiGwWGSWN6F98JPuciVXom8voR
hcRR2ekcZhKu1QimZg6cx1TEbKMNNXd0Egmub4kAH4efoUJ6khR9YjNiHdvgakVf
H6kvwa2Is8dSRwnCcNd4pbHb6MkQkrId5YANcpmyEJyYDygGHfT1njhgBOfwoi60
VLBbIjjOXQkBY3sy7fuQ1u4ycyhiXDTanmDV87scaS4HyEoNx8vhfHMwZDw4LPrm
iejdS1gQ7z7rO2jLDtCGImKWAsgqQVAxmzeGpRQp9fNM12KcrXMlZLWVks0AE2Ko
R6DiHwC8BHwODJ9JngE3NJIJWlDVBwdSyjUxEk4S5O1SYgnAOAn9/AiruyfEatYO
qPX44AnzfLM8qK/Y5HTsLcduQUBqq6Y5NfPx6AsleT8B51DyL1kT5QnTKt4lgUjg
wh5D3ZOvFK8i1deloNBNw3rm45ssVlF3bSlnRCJjPRncek8dbf1AKqQwlsK82V08
cqSGA0wJquAUWq9w0cnz09jR7+BmSAqyDwDHAawNxNPSI92670D89f/fM5cyUxTC
/+JSDFYpyhfP4QWh8/DUywAoWHMbOSPCZitVj6f3Msd1vgx9qfHlR+3Q4wEOtC2Z
czwCMEOdn6rpRVlFQEFUGCkjFF4wQPsibQra/ByMVR6p5MF9k224sLB4pbf2ZWyg
ZrW6yIRoF+MC3vUw+o+69UkJoVb8Jshx7w6h1CkyPB/qyvuuxohkRZC3UtQdBGri
a6dmMI9we6BNuf2RsBnP681ZMs60r7w3IECaH0nPdQFB5EJy3CjkDnIK8G6LYf3a
EqCSWUPf3jEA758ADJjrmrKiFiY3zFZURWYPBaqu9mVBY+VDh27Ufk4V/42BQYmo
KgzmbaG3wjF6VlsPPkGOq/msXoLymBdlIedSLGjoJv53LtSZysJVtOthS6V9ly+c
qguKsZTnltko34q1haN5Sf87ZJ0ufZDdTkooBCE+Jm7aSSNe+X7u9LJ5amly+eYC
/wLFVlBndhCQaCy9qTRIF65gof5kMrSEe/VDo+oW3bHB37i0b9f9E3u7BL5fTM2f
3CnNJd2POWV3SWegnJxyaffhTqSY5NEqP5525lTXS3hWqjhI8JZCq8WfzaTO0c29
Sv4xll6YKiFwKR1mvK+J1tuNdpsMSMlirZ8nvX3Hg28HLYS8ABSrpXUUwHWjPfQ9
ORNqaFMHFd9Vd2Po3pzPx46oVsappx4m/fXupyfU7dxNnK+6iCb1/0Fo/9kLqB3x
D3zV50JMftfzShszl21tDlhaHQ2ATSQNxkgC/RmZmRRQViJThB849hfHx1PxFgJu
kJeklRKFkPIn0nQMnChQ0VAft9CACduD0RQF+vSWlnE3Nx8bJBixTGCbXBBedGQH
eVBpe3v9//7ELdRL/Z+zsrLvcjTxtShStnU044JA7uKA6vGzIiMWEGSHc0BN9m4u
14kLzliZVj80NCzjCtY2Z/YIXueqUuZuCOjsvVeoyecOP8dKHAlZJVJuZt0Qjoa2
hn2y3ujV0zvDI4MW6QFmfVD6nO+G1Yy4DMaEcueM9WkMT2qa+jap3Wj0qz1Ob5Bs
XaCQvvRoRpkpJTt3laWYZD2eLzuM3lNSxapFCCR2GFZ862nGL/lTHCgQ0oKbn3lm
qBB6xnH7jSFq4zOAi3j2XMhOjbY8KAyEmeQFI7X4A6nrW3p5I8wcMI3q4tVwrNAV
mUKlaqWBupMopKqbomKHS6kqdL+vr82tMFuzl7xe6eg2qvr0YE7bcFOgqgGCrbLV
9nUC/hpaqenhoDTrEIkSuZLq+x1iZC7b97thfDmJmInfxD+aMWqrEoYvQ+HALDNs
D8GTgiabJf+XSyHdjmFkqrhYZ41nLWLdK5vjbmt+TpKXe/i/6+446dqfwX6eem1g
sXhtJgjp7PWJ4zZOiTArc55MOHyBVoOf4ejfQN8bR9Cd6hhEyAClk18nz1lFcPec
E5rcw+zAud406UOuDRLXsAyeW3qIEzvLh8c6eyNULuGwee5K/tsj3vtBs2eniJLm
J6yc47xzlblhM1Q1ZjsoS1yH76asZ9AkrjktkVDlZEbTARTHdCJGvV3NiSB7/tve
chIoCHyehRM6EnQCaVeTIXqOcukrXL7ExwbWvrbQyRHlUxyNrdZFevF47LHQjoe/
`protect END_PROTECTED
