`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hy60MsNsQb6gXFkxITtJtg2RuFCoBj2w40PXu6KWQ2mAgmjZjX/SpP9U7xRwDAD1
zjC//vFruqRYcpXaj29MGel21X9+kL5dojaZui9dmdPyVmwcOYzKLU7XbSpaGwop
B20xlFNgJCsXHP1HHz6Axiq4ar5bp40QjqjID9T3dCfyDFDOnaHVaasl4aWGiXSs
0KAJyn4HpK3hqcW6HoDso1TBZPmeL/Fn/Qsm4qX0/8+VoCYKa6Lc4u0kFDdR3YBP
a6z+Ae/mp3xYSs2c8/UrcZfqbWyDoeqMMDfWZSn9cW8hWhXeo9KCa/39G7qhhsxT
sqhJ8DngLK8xIZJWmxVrpCOjCbbHc3yX0Oskk+jweUx+oKKAmA/2C41h7XFIcsB8
Ir0xeLo0Z0b9bXbNJUWOMxq1bwikW7r4rYGXUJkkPNMyKIe+pPDqIsGzfNAcsVz5
7BGAtPxst9CmqwNWJC4CZoZtKTytzK2uC8SIwy9fLMWevdeaPYKE9aaWpw1j2Q2H
zEeBF0PayQZ2efbZREbFRrP4z+kFAeFTlftQWbOEpubijk/0THF6H5k10W3RHtcf
ygRfJApg9IGDl1Y4+T1mKY9cCkT6DF/vTFLwJq33mjyrGOTHQAscwBjlCNbhLcpm
Lnc/aXJfMwqVCqKpbSkAWw/C4pZaiqwGFrhvP+N4yTW3WqJW2UcX+ww+bbPPQcc9
xIV+mRGRlt0RrPCHkUo2cFIwK7St9AsiAbAYrxh4PxY/fmCYsJZeYstAhxPembSV
sVihiZRgHEUAIkm6jeLeeWKt7aBAuTRhTpczH7NLpwd7o/nFID6m/62JmmxmUzU3
mvnx4IXaNos6cUnRH+68zouYpT0xIKGGx1+Yc9ma++JYTvYnzlSavdyFeabcQIE6
86ZikQGiSuMOHTc60xfDVsnAgWhLnN2332AWRoZ3yO9erg8EHVHUbDp95WakvQ9F
OhwhojdMqcanwevozwV5ZcsJyKwUW/W7YstAKQBgUx6i3zfw3DOeAq9uN6/cHu6o
c2MPz6TPrdqhiDhaU/6bKBF3AA6kXPXooCEpbTOzyC9JlFRH9a3yRyhoeDCAB4aT
7RlZjusP7idTpMEkw4B91vUn4QwoJY+JRhvGP0omgYv4WmzDDJGT7OHmqARY705u
4F4tSVJWEutBs1IQtGqQQ4xOcZKJR1w/kue+F3b7U/LPHxG01F5Zm4AdHI/0ykKt
Bsqi1UoB16inBDqNiggem+HHFX82tH6HxBT5u3aS9jPignewkii9arBM4snPpQ5M
FvLzTvDXSLP1Hr50E2aCIH2SU2t8+VZd2toEbjbt6pEb2Y5Avr42qnUe5snFJkYZ
UjINcKnjVua4h+aSCyyckvZtlw8hkuBJFrPPWND44kEWMpaTHcy5F7yyqoht20B/
CggOKUZGy2WxSTLeQDRITK0LdX4CJJ2X+MkmrjEtBEsIXnbArD0RxN/m55s8R7cC
AsnrIqpfaU3dJn6B3xaNTqfZKjh24on1rNkE3HQGiqiTHEAQ8L0jSWE04L6IZaKw
Jfj4NEaLs44ORzp6/AZzYi401supTgEQCYm7D2JtfpNEGmEMLvtAK338jSpuIrFh
EyBTV/uJOkJc0ycbHaYpNn9gq1EQ428VZrLfb/YwOOS8Fo9vVz/EQsjr0LWakPAX
uRtKyZ9Kz8xca0fE1KVDHlsFSiBDu2x/0Xe4T1qzA9orRcBsdERo8k/T97sFD1Ra
ktC5E32iYO4+rIGmfPWn+QwBiS0pjk6LRex31q1YQ/elJ5miFss7lV/j6RjwsVvw
np7bOTkkbmP+JeSthdmrry/exFBW2qRuU8r76B1EpvX/R3aRwJorKBAEvC3txsfv
xg1TC87wt65uAzNEcoFrCxS3J5LVNv6/wFiCvjlGHAzbdx0eCriHV88PBKpPgrci
CMB5+Igh0mshpYLPp8atiYuh0QGSRrlc1dV7KxVdNjCZFuEas/a+tqcpwUTO4fKM
vvOzRL9jE966uriWx7WyMJN6UZdcA2ioyEUbCRrKwZE13zp1IcryscU+WuVX7yTR
OM8alw62u3kpXr8FVIIDGo3N0gHG9kF6DuUJOFEKgp4AJAm2xbunLhjzQ6NCh8Bf
2iDEJKoGECGwVhDBIUr/2RVx6gupEhgZ7ma+PPrmmYYdy1I2vzwWzrekL4fU6oYW
RH27T+UWWpH4rByrQAsP+FcMlRlnfFrVRKAU3XYOO2laY9fvq00Jq9AujgBMMB3a
vLCP1wxjBLrSGX+O2YIgb0EYG0xyPgkztsgzt7ctNpwjSgFUCuixWRhIRzBn5ZTM
jPlKu32sOyuuyEpw78hgwV09uqLF4LWhtfpK/IaZjNMRs7DUQp6mFdgDcRZVlbQY
JRolXLtKnYaGt6RKx8Xd5MPkoj9VFyfyx9L/6HFpB3yJt9MbfUJDouxhelCaNLAU
7FXsOX1pF9RoJLmDTTKyY9hLNnGTuc6L1j23J3hglRkiRitmmee3OV/QAQvvObeY
toKtvODqkH/lqC6hsrsers2sU8TS6MBXDnaMmrRknQocaSdCvbkGdzXEptu4aq2z
B1auu2OkjIb7iTHQvir7w4kGJApR4DeY7JGxl6BNpT2png9trXvwqwJNlmk+jff+
zBxq9Q2h6QBbfPBOX9d+tF4SYuQvCKKaUn7d/xrer6CEyxhQhXp5sgTx55EfpVl8
yWkfunoe8wkGkOu2bir2SJKuvGpUVdD4CQETY4kCJFKAuIcID/R54tyF1rDLgeog
Zy0vnXS6E8drKSQFqFJm7MjoUfiY8oFodSI60oiLErQhYITFuBO3/HjUGKYQ4RqV
oJ1HE9H52LbBaeSPZ5F+iEuA59epS6h4hsy/XA+RJ7RqWx67R79wlv/5ltztu+4t
IQTe+uUXcex21RFF+iM9FCmmH1LElHDvzExxeoIVo/R6vwaS1ruk01IExoJfh4jR
NOoLmn7v7ltpKyRxVulGl6jdVh3GOUmuUdgTVUvknJL0KVVoyAU4SNJnFoi98hQ9
WTCYuwMRIrlVICja58dk0/1Qe7xrS1Glr4qiuFn6bm834r9c8Ag2FgUVFcMWH6wt
dYo9uoMPHreynbXab+1mgLNHpj+Cd07j0Qc/5nz4CkAuQ++Utp9wqPEnhYOG32XI
pUbHzgD8K+lpyJkkR44lblg7QrMI39IUjC2Hr/dUcOPsCbc60YO3neH6YCDvIGsg
XYxEheELhT1CF49vMLU0JQfAEmTVLZdxpChwXnBDRJvw7uIUZPFfsTGq8hLqBtBN
b3ul4F38fNBP/w+PZ1n+GfqwQaF5MWa6oe6tElNnSBxGhnli1VMi7fgb8A4AlK4r
OaYkCXvYPaeNfUzB4RxaxeTEt+lSepIjeojm3V5ChCnBHsuxbpkkK0XGCADo2vvV
OuTIaWozAHVu5JcrF8eT0AoZymCvTPUMWk1N0LtyW99BypNMimIm6LHWsW/GxszY
1xvmhGpMKuqiVAMqXUi3ZFBsXXHCvUQJm+qPo2Oi8QA3waALBDeVRl93QDxXMgYL
Lkve+TRZHckXevMeHPCihxTKjcN2yRTeAoavC9FK1zJk4lXiVsnKOFsjyIFch7iC
FVAOG9XtQTwgpLs0P3nbmar45MZHRf4KAfQMJ2DKAKaZGQhuac6YOTXNqdrNy7tP
7YszH13/Ku6dSpPV8TRorjew44LkJNcMH+FsrI1ukvLCbgidEGbC0TtcilDkKUL9
rB/2I8CxdaSuZuZPv+EGkeiNviTqz1aW28lVpM8oPKRu3aI/FGZUqUMKvhfHNrwn
vEhPiFxUZae3AeXhEfqGM8LQjkVGEhWyYkTEWRS6ygQHcfciMzk46gg9+vd1CLPf
U+DXT2Ozu9g66Kyr20OlH0dSJF+rzMeJwjbJd9Sl5nXyOYdrHkuhKa9oo6DQFF1O
EuSOcsZR8peQs6LEeRVM7SjourCsU5ziFisFOv/4E1X5y2bJqqqJZm2EUkgoVoc4
VZ3srOByQd9ERthkMvEi8+fhBm2O1G55Uxz7vW9tX5rGw02N4nvehlQrn0zQz4CZ
9jDedjE4u4NGzja2O7qkrNkEI0XW0jGBSqFCgmy18oMsOZdnddgu9/mJ3UuEEuWe
AkVkEDVnX2iw/LMge60xkctA02sz+PT0SlNmMwbJrtLRXOCmA4Qxe1g6A2xtgn67
zCDxXTXfxJ9+VFJzQTsF7za3bGDXmgQD4yD9vNX+QYSbxeEFAX6ptjfm4wVU+zCX
rmcFrpvopHj/pSr6mE1kBR8weDQ16y0bGYmKtV/WUT3KRiFG1u8EIXhzPJRpYkCP
aJ2UZMFShpFnudM1z0tdxYlzysqw8oOng4TaU2wq731DYfGWrQJK9A3kGZVimG8Q
10G1Fhq7fm3LcntMvpqwfgAHEEGVWjXlULBXZfOtuWLGNkvvSx1++MdLTPitiFlV
7Y4yXJ3Gbw6OWxcleHzGYihxhgrOuIETTwfJTklSadMZh4mzUVsE9NetiL75a+Bj
T9231IoPuH35kqWfiY9TWvDSHglBG1Ku3l7BYBIlt5sab47ukV7SXFtG5vxY8feD
CP4ndyVEyfSek6JJWkTianoJTO+FSiwVEZ6qB5KhpEHMtqoRCfIvBHUfpTmq8gkU
Yoei1joMEipnBjEbW4TZQP3x4ucmxLdxB7+O33IhB1l178w3C9KA2Zk1nB4rNWBY
0+6LYFcWyXpIZWuzEpd0ulq03F+4DxaKPJx9amXPLzsSBreIfMB+Z+wrJ0sOi461
SI42xzK9KXRgu3Z2z9ibTg5QNLxoGacd1q8/hDZuUBrTnuKyU14YrNFjG3sGH5oR
VSVHn/lGv3nX6OJtn8OiU+o/u193aITjZX0I+3KJcEERmPNP+4RnC0KGzqb76NNA
ZM+T8LaMv2f0vi2hZzBs2l0w51x6SLf46Fx5fXs2IVZ9lRaIFerxh2kTddRVcfHt
c+pNZrswv73ifdCUs80Qm+943JnXoqIb/k/NrLMTvsByfNi8FgFFhAHJbbCteUSf
OamfscPPHseGEmmwX1uuCn4WLuxGJAJLJTaA2oMCrDz66ljZltZKfPmVf/NneTbI
6I9v75d9g01Jrry/NnfXN3I+qCpckaTrPE8VhaXRzhfIfSIIanU2y2Q6lhLBBPSn
7ltF6Hajl77jHoXdkFrVamVFivmMoEkoSS+P74XjTXCSvy8UanN9/Az1LbyBQ420
o8FyPEdCrroJEX9BJTyfS3gQA9tuIPGvusW9DRtlIQ41pbiYaZeCZ2Fy6Ig2rtgZ
eS6eSmrE37Jnb8q98ajTZ1MHdS81rmsBhWtTUMzn7FOFtbpaplJGEILtghh7OLT2
vSyZ/pWP/PpnxA5wP5NICJeMAy69at0/4b2JPgr7DDKlsMFyjWza8t8S1apLNG3U
NLMVeCx3i6jACNjt59AZWObRFgvpRCEb70VlXd2cGXBaBjwtJS7W7ykC3Elnttlh
VegKmNr6MqFRpqlTABUNDwDxwn5GlDaANNuQlagEAb3U4qO8JRL8Som+GY7tn4WI
fsTy87Wq8MGDqw5FkYwt32GmghyTZd4+9Y0e4O+cEdlR5KgonTOgaA5wQ0YmS50x
ef8Fka6R5Vlfi6sKirfMHLQiThnZ4325Ta3FDxli0/ybApYiPWBRo3cuZ+RFE7kH
SnCV/SJ2mn6e0NoSNa9WfewJJ5ue7snwrdOJb9SHVMdrXDQGf+oULyllibwygNd9
htbvFO+tcDNHmgBbSHxuqs/hxH1cauBKheTr93Oyl+dHQ1498RFrl5ZARtdG7//E
/uW1QWAwRvVN4PeaLQC3h2y58vJVZj+uTL/9AQJ3p61DNJnEXWqFIpucH+ptb/3L
DRrcbiA7XYt9fchNCnigb1N/VDrr7sVRQaDKTY3h2Amsnp750eTVNsc0dEVddUk7
Ybz3ZEVuy3CGyOeKUn0QWAERz/XqQfQYYzfxUCqUGfCaUNegRg/c1e5k1dwUqaOr
BqoP1s4le4xKBTF/H1QHSPLFpzTVHcfQatowbfQIwacQo+xU3JWSwz0Wngoll1in
iw1eLNZrnTaBeIWzoYalJC4C6jS3njKsisgcEGmd7g3X7r6KkDBAmjXVL74yzKtg
2QjpY3EJd7TX6R2MLbEISH2BVwWqx0Z/74x8vg6tk0KKF2sKN7Qto2Qe+MGom5Kx
mLx1L/93Nwn1BxgB6gP6qQ==
`protect END_PROTECTED
