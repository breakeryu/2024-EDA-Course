`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8Bf3Oy4spqGG21+9wk5Lv7WyTzAy+uJt1V2w/8z+kpneQ2mU+YdzSPvwbRZQOmQ
X0e+ygQ9PmMmR9s2tHeiqe2ORpHfwsIo0hr1MpnKFAZhQHhEsHe6EPY153Jcm2uW
FAfn/0sCIJ7/Ptgw3FpYH/aQ6gSPQbKgeAlIN0sFB5iMMjyqRaenwyqEYaZjiiym
Ze9xjOsykM3O66Wyex8FCc6/vF5qMBpEA0qXzP2NQH0SDanhJFdsiHRP6XYnMlPC
DOGGQacWabJ3EHBt2jshWJwPQfkmaQukQSSRc7/tOsXRVjWIwtOOsSMqullm8D8x
Q9PFP33aJ7tnAf1GFb6QPc5tKnOeMnuCRTZtWYRcd4OHhXOqx5hsP+G+XqxrK5DI
`protect END_PROTECTED
