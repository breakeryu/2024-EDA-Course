`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YdwxMRUQyeGjmE5GTOnPbXqzuK/JbJ5duEeTz+6Vb3+VzH5Zyi6rPsY2WffMI3h8
tHRDpniZFZWTKtXTk/29xZBJd79F6LCYd93q8wx6jflJvSOgy+9DXTYthImI3M8w
cxbQpnjvPR7OvoBU06tPxgUaD32cgf49ivyoo6Vj7IBL6Mftt51pQKN2HuA4HxWV
LNLxuaD843uHke8kk2ZzeZvTKTAqkNvBgOX8STjJap39eKB5tyV/epcU2e6rLGBG
bEGDLhFSXpA3Rh/4RflD2atMhkEzihR0ZDn/AWkhUw3JBuUyXTO+JGa5wRrY8JzP
bp/gv+u+sltda0LyFKWB643j6Ph6otoadn31+kdmnrBNxFyWSiBUOvVxYIwVfcFh
yXMP1gb10Zsy7wGKmgQNAgUfa6jcBwQfgoRI58ZKjRT1qDPi2QTW/DNNZQSKpHpg
mqWdeNXv5InptrCe77Pu/je9WBqOpZDf81Qx2THzdeqQ5iN1ZPQEOj8BrZUlwyZ8
+oeFc0EltRn8PeKofFIrucQjMDuVST8OozNyLFNB2T23UuVWPZjdtBLHXPoV6qRD
itwmNBjvGeFHmh3A/b5D4sN+Kvqc9/Z72Q6ubLJwIbHtHj4a0chhnDh76ym3w3uf
orkCazy2bt/DJ/eKdOnH03+R7x9c5E/MVllckvaQH11MymC7oV6pfhzBZaf53CCV
4e3ZXvA5JuYHEbWkZx23nC8/ZJmlWWnZrpBO63vuNPxxGfAdtGVezwh2Yuz4KfIQ
3gQrFc78dcCK0dFROYi0ojTNg03aZFQ9u0p4MyFL4mCqwXHd7/eugTg8F/w4L6H/
c/ePn23I+ih37fehkGncjm/uM1W6cGN8qSjabyVUZNBPEgcZLOUK+/a7PTGGmoX3
YtP4mmni3ngWGtIuwNfosuLpkUm+TOXCWZJPuyCD1EEfB6SNXzCcozd2lLXUEIEF
LP2MaMZZ/am1cw3zMUYv30R9dXSpzp37ihsNAgDxsMF5Z0jjzT76kbVGm6v6U1aT
Dnvyx3jj0+wwuclSpjHAiHGPRtkw6DiXTTGi61DtOc20r7e7tH2/yh8+GHBvu/83
oE6y9oyb5trzIKv+WDRcmMWP0nPuXJBIoJVs5JTJ+e71MEs4g9iRkT6rWhUtf64k
HLz2vsNRkfbCdyLvGjg1jGrDgSg0BdYiHC4yqaXQVI6virixtU4yb1JmaMdd/fNR
V+3JiVe4PoNUmeAmAV728hq8v5rwkvnwuDHyOBeJ0IY5b87qETLzAmInJTMGBL99
lTX7uK24C4+ytLRAv2aXf1vQCRPLBV6/+mFUkOxVC/PUb1DCRWy9hqy/fNstScIL
9G0axewOK5fKyY8ParRtE5Vawsv26cHxPa4c5S9M06D2rVH8WWcn+IZhIpI2ynU6
vBV5Yj0tDUemtwwjDye6BhbLa8UpIWNpVaYBVmUeBYor2OqQubgUSljGx6DDJC1F
XbJb6bzkgH6XJy3gIr2/AW+RYB0YIJv7rgi0bsam4zSXB+Sudv1HdYOR/BPwSX/g
BNEmGhtg852ujXUvfeVY16/URg5ZG8qx/qZIXKCoZ95w0VkxfKrSX+b/AT6Q357k
jXFyLsnTH+u4DPDk0gMg4buSMrE6SnXRRv+SqxpxGa3fsqbtDklz9NKI4uXXrkPz
tqwuhuA6oXjb4yiU8iPfBmEVpjlxBBr/JsCOp9XfV+5KYW8ueD8ajEDngcLC08Z6
OYVlk31GdBJfpWZVcUIDGiDm2TIoeWVUoGmRG/Mm1d+zFUZHVx3zilHvVYlTD8aC
JM/dlsW3D/0bEwPDVff/0g==
`protect END_PROTECTED
