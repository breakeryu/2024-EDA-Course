`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+Kbl5VJ9asiVXbp6/2tIS2JvOzfqQXiBtzJZ3qRdrfbmdz5FiLF4GpOpkpq7+5G
LDTnJvkbZCRMa+W8ICMgih+zKnXZBKIHFOTft3psiVSnJBsp0M/iBVfZhRk47Lhb
R60+PMVwnjt/rMsyQUksYye4ezBQFHHPzlevmR1XohuT6IxIyjJ1TQvg7J0dOodJ
k2MEasE0i6wk2vE267BX6VEkzeOMyRJEXdcF9sArRwOBrtBkHixx7cKMQ3DZih23
wpL4xPDGQyJYLkdhy0Vm4tqUFS79Yxp7EXfuhrkjX1m+WcfVMPMuIrxC/YNQ6ixz
EUxBbo/viTLIHru6POozC/4jFgNmMsUP7XHBsW+KhjQVbjE6UKv23nH+6c2GPnmd
POBACyTguV1SMksh/hTRIjd1yNteqAJzGlXd09SHnIYEMsayFyUHGky4iya3evrc
CNQjk+U1axqOBsLv44nvOWd0RTK+GMUh+apDy79dXxBqVgXIt5/sxDyH779N/zDr
+2wgj2yDvc5c3QDORVDScvkbiLNnDbt+H8N4+S93iwoAVW6mmizM4HKb4T4iR6D9
pVXfDkPDaIZ+4DKy6WH/vdmapaZp2ZViENdtkooHgJE0NPVBYESwSGB40mPxchOs
SIF1g2TR3sEg5AisxA3bdbtEiKwUZ7grgHsRHdkZgKpFIVLNT0oINXMfDKaISp12
P2fqusVbUhFdSLy9HzfdK1/0kmBUQaXU7hcDA2PPelokGj3McIxmBMm4Y8Sb6Km0
VG4dA25FmCJ17+2iO1SvkbdJbOHxOgTeLfXddlIZBoFXGsnRmETuzllk2qfaqwHT
PKvd8VJn1m9zY0gtBRKy6sNMaIBC5SncpyucIim/1kcI1cWUkUyEN7X0E6A4elYM
rrghtAIwL6HMYjKEjbBrN2i3w4Z+yvKS8wOw6I3JY1+mTv/x+tw1Lu4VRYxsNnRw
sUaEFTWPTX2VwSyIA3vu0TO71an3iVX4v4n1Cktk0Kkrx+BQ6AgMkZhaDwTp1kN+
RSa9Tvaq09/WU+d/OU4KSfFPIqnQkyYP++KguOfcuo0m5nMLeSv5N4gFNvG0sfWj
fm1xTZxvb8JLZ5gBxdoqXnppc4MQDz03owbXpR7bfNEb/ILEuF/KXx/KtABfhyhh
06b7zeUon6dxZEA3nIJCoGWit0p3ukdojHT4GR2iciRoxFVoQAU9lz1gOSMGYKR8
CCfbBNDtq+WL6fjBowhsIDQ6F+AfpD9ww+u1uIsNTPkh+q4EgSD+3xi5ZmDYBbLE
5LlR9SPvyt8YaL/Ih+5gD51GLbiTZUwIQ+jrAlor1kHFcQ45MUot8qjv2zBK/G5v
ho1YDj4VC7GtZ754oD0D2ZyWX3xuxlEqMOpQRPW51YQ/8AeVZhr/v2TTia/jIoUa
4I0tKy4n4o1WFPuAucewXaR/vw1qYdeDnA3uKZqY+WbwdzczUKQUAQEJQ/SZAHGB
Loj/WVw3bIhAPBq9yNyTfdOyDDxnVFbVnhYTVOmmFQqoVn5NUGBjsHUtpRDsM8vE
YkHMuiWQajI6tVOcHHLTrJ2p5qCQcY5MNZMsWtscNLxLjhbz5M9aa75aPgYFr+nF
Df5mc0nWr+ubIrvucDIxXswtfRujHLcVZ/hEnC0JGNIvx9THbEUOouwWbMyre3XR
fSWSNx4qgYMn1roOP9w3W8lKyPEIzgTUX12Jo8G2nFsaFj70g77WgyOKFXFTz4CH
cd/HeL5SkaFHcSQIRXkspMfzq7/fVG3nZOIqcNgdu/F+ydurRo/VGofrfXJqZAHL
8T9BmCwZ1N+kA2HKNZzLwn9xrbYp+jfahZ0Hgjj6fXbsc2Xr4m6aCsDS2Fu8kAZy
sLL++R9WZx/JJUYW0798lEmU4lYPiSGmeFx7dafYPmI5NgopZzkl2hTdSGCaJ+zQ
yuUzVWMAX9oAZRItS17fvjszTVRvqIUHA+7yVoJHT0GqtPc8NUyVI9J2s3cmYaH/
MdcoBIeCHs4PS+mWH3gQw32UrijB5M5y1uE0ti24ZcRiVwyMFN0xr5kr6IwQqe40
vABleLcdGe201aLkXu6UpvnsNFxICT+SEWnex42ZDY62EDXTNA3n38fhnuUAu4Co
h7KwImBsEt+dAq8bDW2cKsApzi91DYzsnYid7pEHyzc5KknK8kV0iGIFq9Bilo4f
PPJ3CWXivwhhAMUHPvhJO5d1K3j5v8TA2k61laiXYSSOKECpWD6hWPulqfVB/9vy
EkwbKLyHnBa9UMHb9uDSoWlb4QHH6ppSydllz/yTREM/jkFdH2ylppVVqK8xXK8O
oW2/WoF6T8h0h3xkQs1AjthW0Wc9RSe2zwJMQsCUnj9IlOMH3QojG5hpjD7z7+HK
usR272s6SpnW2fi35VrX4VhEaZsjJ8T2U5WllNj1url2oG/QvD3ZHKaS9Axhi777
uSOT4u3lIFhJkX0cPyN1CKi82ERIRohH8+S6okScky53v4r4x52N5UQ4z9aYU+gE
fsR0QkVLrWqg5wOpcCfgHlIkpIu9j6dXooc4INuVVehRGcqDDMbS2QJdB6FU2pf2
G9Ur1iXkSoso9+ajCep2v4V6GAV76EgVEJdJUP4G+PH8FsdEmaIVAwM1PCfDEL+b
YC8ArZrJrOOel8ZFLnmLV1+E2bNNBiMxnr/iJbl+dsj475wEP9KohofnRpsR3T9K
aUzARUVvtRVjk7/4U/Y0RAYsiNnPgFhg+tDTpwUg6bzMytnDWAfuJrL9u9aL5Bqv
lz/oiMcrp+k2l3huzcmUzRAun7TjThplTYZx5xr7atWmOpucWoAntCSLGW6rvNQh
CTTzIN4RqTmbPTN1+vu+AkwSSQv93BS2/p63jYlpV6Aw2/mXof+GAdHYqfKXViZy
wa9Z6eAF7S97PLJu0+2V97qvis5ESombGA6ded/nJrinSDch655Eo0Y/0CvL9lFD
Fvo4b0yqGL7aIyl6tuj2AD/61T+789Ky+P+TofUypeAQFitUxl31cLtXdYuj4P71
uEY+i9uOw7AW38jfg9na33URa070GlvQnCqjLgxhDqRUXvSCYW4yh5TSD4Q5A7Zv
Y+6paqMa8m9cQKKsMRphMVNUQij2NoQQiKsf6NN5GN6Cqla99S2fOk//Gs7eHuwr
CSEgq8VhAaN45+Mr9h7p9gyOLy3jEgJPk0Rne2AIqvYEnfWStWrZAWobiaKvNewh
AMElJ4kIx5U2GW/l0r1LzAKwBsnHRsR2e08sMLVWg9fB+TXPS+jseL/Fi3ammWHp
UdtEHNzJIAKQPht1LGjelD1Vpc2yHc04Z0dXJVC9JKY6IXUm0caqu3iLai3IUw0J
et0OdepYEvMb2YOfjfGpSb8oefZjbyzMf84cKNCNCusFiVDLd+jtXjKhtaQFvj3n
3bVAHAgQSVw2doeotn8EQK6x3z1bKPdDY6yc3gZjB/Rcp8dNyxfiaN5Jii2wBgsR
2itIjzXhgIZymCtUxfTtAO7iZS8j7pmgXQlg83cMnCY6iTdyzshsDs9d1og+/BD6
7sj92ZLDtWAUYEH3tAp57Mc6ZZ8AoU0ukM7uUSBmI9R3BKEFY31o43KnEOJ+8+i7
gSDYyysioHYvlTnEAcv6jEIVuhXpS567pVJkIuYm60pdhMjRtfUkXevU9DsHU7/C
RJxtY9hDde5mjp1l50Lbe+4Ttrq5XEOWdMazv7XTiJduPLZVmeCvctgEhwx9XobG
M1SHQ1dHLDzZsDtvqF540UBpVskdgAS1MfSudTO4krXFLMbFn9JVoEEY/bToIM02
Xs8MyHk6FJw3LRbn4zh4z+1X69+nx9Cpg0RbVDNjnJy1aKgluitDJMjAYOK74Z4P
2IoL5XxulP0eVjH0uv9vONyDDbe41huLLNdzcTjGkZe+xA3XNSxEJYIVXEEmHHa8
Tj2qy+ccEne00PPMfGufJT6gEuo1hY2t/tKYicWzdp1fxLo4OuqFI/PXM0smLqnW
MpnDeGcAnPA5wgEfTVxUPXKSxc0g2y1pvnxT93M9ETAWHZV0jZ5U4SHXFl7ufD8M
Bv5INPjCNohr4w3uDkAX+tc7v6Q/lLH5O9hz7PvqZA3H8w/kPBGBZYgxVbEXkGit
fFoN3Io/DzgEBnXaxud5bTmB2kldcaGJu2uaIwT818NbJ9MZveTgK/WN+jNJrVQ6
WaM4ETcNOKA3HInFrTOhEQMjnZ39By7YBSntanqo6RfyM9JQdEjQhQpGBhSInkAB
JqaZWEVsQSLNiJrEUze0jqLJtkP5tpgaYSh8SYlyV8wB6uI0IBTPDWzzdqaTLBxz
I4JPSnkKN8inQzoYPQ2lxUgmMglL7tZrhdlsoxtcVqnKGaoaUQBMNSeexZ7OMRlj
HY7PqSonb/TM21Wh8SwbdgTSchBjc1NuAW+pfsZgu5wtsOL5zhJotkDkntHRZPGn
Ohhw8U9ljHl5tqvuAEuFpzU/RnV1VRhHJC0yul5clHDmh1C5wMFsn5o8b0T80x0V
rQB9l7fjxCnNS1tH17z9ars7X5GPT0E7PhseLuLV+8lxOSR6Pr9zGMbfcsl9q4FI
R1x6rYj25r8fVqQD2c/VPXaPcS9cPY8BKBprd7feQNTkmvlFbtIIcHKXlOTQ21GZ
z8V2bqnzNLIMQz0rnxRxE47oG80gwOBh1zi3TWk6kAjciU7vZQBTW4Ghx5NfGjp0
3oJwPnyTTkfDV/m/L6Dxc264euLahTrR+oC/EPEUzrK9XcHSuHteoDGSjuhPREs4
GEAXJu5tlEv9XTbWlZSZAzNnDYGLjIV7wgJ0JUzf7ww/oSgSZ/ZLNexjVSJh6olu
fFNV2ipGOFY6fCidQs6rPEI6H/l7OBN8tK+eRD7tffCMzaqEDgEWUDA8BTtTKQre
2jaloaYP13JA2F1GedMH9Ux4MDPo0Ony9OpX1yT7HQGt2q5MTOecYEIspeQreIl3
dYRkx6QmlsssnIfu8j2BJP/wR/p8NrVwZEmx5bMVKasU/j/ww/x6hlUK1mCYIKxt
tPewYuWpi2K2D16rYcdi0uxZ6IJfC2zVe6XuMR2Eh7XaEDzXebvJbzWhlwZkxbwD
9dPyuqReFEslJQAKCidSMkae2sgsySMsBleT9sUGak2hVuZ7acxWuTPk/+ZIzYHz
llGo4rWtcNnPBQ7VYhg35behti4sm/sjxhms6fzr8u3sbXILSORSuS/IvpoRtu4I
pvUse3wRfQYtD4WLgzyLedooNgKWwKeaADcX0GLIMoKeiB66ctNreRlUFmhjdLXl
Erute3IpiPL5Upc6yjeJeijF2VUmxbAww/qTnGlz/CNNcclELYfxtDvuhZYKKgeW
/QTvkjc57IdaCc1mWzJkGr+bI562Lg80pYsMbgZCLSRgvKoVPr8/QDHXMHWmXC7F
1Vau5FBygudbJ13/gKWpU8nz4XmZEhe3kfnNSKcQKp/z7QbNdTdtTTh39lpRJdIN
md3D4N7TI07wzaz8HUud2GGqiHv3z3pb8AQ0ogUqafAthODCLDW+y8eB2j7zXEuj
ho2RWZwmmvOfv/8FGtw5BilKENWkB2ZSNmUg4jF+YtxbuKyjUv0X6okgg0GdntCZ
Zp5yKqsVR1t4IMR745FdRS+V63l4Arv9aqUPxL8nu8KwQuIJLLJH7Vu/Me1Hem9R
arBxxNq5Nv4MRF2q2VvGMA==
`protect END_PROTECTED
