`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmOwmoMw2BKaisUurSFbD6c99vzq4KRjiC8Kf2KXRyDCSpLcCKbZWTsyC1dQlD2S
V9l0m1+PW/rQM6hleSHQl6RAgaDy6Gi73lGNpaqcjo9cjUPTxZZISpE4AmFGUyto
qBVkyOz9JseGX+N2rucoEPT7qiXiG51XgPl5yLgXhFbzcICMe0E1ASYHn20btJv/
H7JeNQyB+UQ8xal8uEK/V/r7dLssH9PcueqUDAsV62NulbUDRfE6LJYNWdY3RmkD
g0AwMfs5ADlqPEvnUFdZ9xhQvnFYvyni9jxhgSGharn3icUElz7LeWv0oFj3c/pG
6SQUKXdhekcYI6RVOmPxZXsh84BFTNWLJUajhoTINuktOYP4iMzMrk2AsYViAoCy
GfaewhFB4fbANNNLIpLsC/iPUqQKr4SeGjUBwBiK4xDu5K/6UgTiaz1GIqLOz1Fq
sWvl125pATGDrPyubrTeccZLp9Djr91AmdmhQ7iDe6Q4GBwtKAgn4baCmsQ9kKoC
PETDyWfWa++QLjyArZjDbgsHpDuDPjxbod2mAEYQYMYn+eM+RydqVo3qOddXy+k+
5ZysyeIInREL3ELmnGjesx3u/ykACYI2lCy1TvFcPEzNAW6UUhB60LuINCcIFmkl
eW+A++WHS3xoSh/SnbiaKPAzj4TYIFOSQ3w7PRfs+gYAjHEdKRS31E3Es5cFjbCE
7dgqGxgbVLkT+vhcoFESK+j/A+66Jt8pEDD9yL2tqTpjeUMouoQmchZPMx7/Htng
ev53JEPjZrV5IgsaKTYFO1d6mJEiI+3CCbjvE2GNKqBz3jCnUB36j1JQy+O1pWd1
75toYQ7XzQ49FMoaJaN5AGRhgGYtCE7NNU5D4WvCjGFz6ic+c88blxJHBsuzil9o
PvJ3wCPJAT/TlK9+8hdQGmynj0lh1Z2gUL5EH0HV/uz5DGk7XUD8DImbDCxUM5qZ
TW8LCTdqLwmyHF7BMwV/3Nm6lWt0vRMPBrRgvfx0ylZjW7Oqpmg7/qsIVdp0/eEA
SSxouLSDMltgwZRAkQczx+82ZSQ0LdwJsOZNus+bd5KnCw9Tz1Z4Z7IjA52SyzwK
VtehfPL17HAPh+5YwtH/AwBfk5YAADX6pHIvr9knb0WxvDgFrLcVtt4t6TmDJ/9S
84kWDHaKKDAR0zox3W1zbXpL8I1cRo4RkBAOOeULZmFvD4FhOwVlWy83tx9y18Gw
80fOv/cIxX0e6C6IwRZPpXjpIfJ33UpKfjyUDYX/QMHuAX4IxzftmAaSkGL2PV4T
1mIQYyO/SuF452y9C6u9Rem9aY837CK5qcs7FQO8T0CFttCnB8GeKIGL0ewJhplb
sLRiPmzAFSRZpIXdHJXXuhUbbFQnQe+Wsn3JEOnNEj9YftDAO1iUnqU4OdP+kP7s
MBRUpdwBDGyrP9E3R5L+++JLap3MkKhF3uNZs08a3IxazhZ8CMAmUYdYrPqNWjg5
VRqJf+MWopx1kFzspJQ3ZTcyW0c8N4z4dAoBmxUDw8goOPufCCxTWIqCpa7bSTwO
GmnL8SgqMY8MbjNuyHXWbfqOAH87ybUrHN4nClu4o6P6A94C6EI9rLm2KgfUQDRA
BJUxnKf3LI5bz2zpiIgvyg/+cXJFi9ROp4kR2+gOk4YONtzJsq8g7dZSZ5idEg4K
s/rdAPLipWfL2+Om2TrgIYu08siJzJsfOJT7bWQwz44BUcdjXkO/Ibqp4Zc0fz2J
OEvNQhu0UYITOhMTMxgiK4+6ID4HbEyxTYEhghRa4wti92RfxZfRd65VRoFpD+F1
Xfn9tNkchi4dXQ6YRL1dru3Hq9jhgfMrKCpuk0onP8FytE2g2ajd4KCJqkx67rW3
8n5q2AsQhBM7zOCnna8GHG4vVeSRMWQGSH0bC+A8fx7lLo7Qes2xBmELmTsE3wP0
J8UI3Ex8KRgMf4oGYihPh7TFnPBP41VT07UhG8FffCUa4+dvQS657vnkPTjmC0TP
FqkA4o8uvneX5WjcD+ii3WLaGtMhghlLipNgHMi379SStilDqIf/bmCySf98MWu/
YjJFzCJW3wvvN9Vb+j64p+A1GtF0vOB013zb5ZlUUaa71/tZBjC2tw6QHjhcUj1C
ANOoKMuBuzvVsYHAn6u0PboIS3+QLK7SGGJa9mFqJE02yXumG5Zy8a2WpJkw/5z1
N5R/hwRxs2AXfT+5Fwc6ekJWpWZVBPx5iFebz7I/i40=
`protect END_PROTECTED
