`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5G4EFCmKolCVAbvs1jgB0exTtr+AmJ0BSr2FKZUgsw/Febg6h0iXPNUp2MDlFlJi
ffShyvhc7IcdB6llXXCTPPigNXFWOCZzUfc07EPHGgiaokmkAzD43iRiYBVZtKTg
cHzmUOkYQkkxoi2HuAFW1sxph7FdXNIwmkk7LRP54KsQK1qfmKQQLVupEREk8cli
cyFMyW9Ye22QKwHdtbYxw8mHvxvod7VhTX7G/b+ynuiA8kNm/VrLd1mkJ+ywPABf
SMIp1o8wdOogHcn7fC1/turayagvg+ohdg33iG8t+PHmlOlzCbvG/ivU4o8jdiai
PhROTdYOk0MG48m4vsjrdF8VhEbFiQj34wqbj6xraeA3yS4fpZT0XkAJ2/sl95sk
ZoGCze+ot6dctVwWBy6CtzLedfQXmiWtUgyutA8+0TTokQVyseY3bp8Afr3mTEWE
bzOp4orWysB5PgexHTFKCwvRpF6sZOyaRcmSEAAZ0umcppx+tbJaYsCxAfkppCbN
yzmR1U/ki/uNYP6saXe1b/yXjsC83qJVhxtsmzfD3S8NJ/cglD+A9YXDDbpPdp+w
GIiVwCdtitWPwTxZqSllZYtZAAlFqxRF2nBVJRQ+kjNLmnb9LWfft3TpmBmnP/c2
3+Akg8VGFOFDV/xcbR2XTcj3k+Uebj45ADChU8n0cI7jYFLAw9+RjHnfl6S2j82A
ZMBFh6p8i6QM2rY3eR7+ogrcXIL251n+NtGuWxLPBn9YJcgD8ZXk6ffOJ7CMTDDG
pnUpAROXGthxQXC518s0a8KPmCHOV748HUrTAYoclgw/BCgMHDrkNJEnvD7LQ92N
Tv/L9EVfNhiRm2NZA+vZ5NRCNSwFEk9ug++RY/FSpMMWjQOU2OIiDz+vgUr+fIy3
jpiM3vgPcenHnLoHAlOjorD5NiiDKWLhc2yQkXx7xAqYMTO/E40K5NYkKWIHv5zz
4RPpSC+F3jxwidu7J2LY9Mm9b9+56VrFY7VbZL0Lr32bUHYk3GCMawjTcszB2BaR
Ma5NUyb7VnfshD0azIN5+tWlAAWPDPb3i6Zh9xfLdYDo1ZPG/ePCrxYlEMgYj9w/
cLLWefHGs9XF8jOkdxdcwig+yrIEtoSpaPbmexHrzxnv/H+mMUznDg63XUfpRfE8
f6MJwraawqeJeSItHyGcG7xRpPIhf6qIQT8veytmdqa/pXSC6Znhnc7dZbHtzyff
KMWv74pc18iV8e05vPkMu2WoFtNOUfl0GCKObJW7HloJaa9tKBBlQm8x0sAggs7U
/8wLCXk0wgMM1cquHKXZFEPeSI2iov/YJ6B8KD/w5B8SFo/sDzs6HRWGfBgd6i/6
n6Bal/aSdlEmDUe1JPZKx9wbuUpsS9hyYd7wHcxapwOZokLSCuFFXs4DVDXaVPY9
1/rdhFa+9rFzkW60t+s7i5FmzjROQJZpXwNfE9dCDO83dlYOpY8xGygpXZxprufS
0Tc6W3KrbnIBu7ag/M+Uf++N48Padxy3DU/3RyYlq10VsMxhiZnI8SeKnXgym5oW
CLLX2qEmi7UdG1VKNhNiSvPGdWwt7zuP1cxxpA2zOmkSkCPnuFoAoJ/73rIzDaCl
sA0KUVfZbb9SuvTLAvxufmsiSN3H3mzrg4DnKM7Hb9whRdB35gPuCXzBhuFdL65u
rkqxAzMjqp4YuUqVWPakFfhiPGCcNmNFC0Jd16DQBeP0LQxmrL6Mz4ji8/a1wrGy
HSpe4aLhcb+40Xf2NCO79yPlNJuYL5rBoFtMvLFV9apqus6V/C5VQt8NoGcgFIo8
qAfXuiizdZykDhyWGT7JHU7pepVhvvwl4Dde0kpAw4uGD26AxbURF7OIm3MMlXL+
Uw8VlZCcqZCr4/QSSEIYd7yCE1qpQyJlJGYJGoHkrBjxEK3sX7psbQ7/2u1WwC6k
j6IAX/nhRdM2zEC9iEegyw==
`protect END_PROTECTED
