`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drLwa2WSmjVmkpCA+HRurTggKLXmt0ZU7sUk9T87iE8JRQYqF0VjQCQ0iS8TBGiM
fKmfumvMnPSRP3CH7Ax+7gr2WK0mYhIIh+L3G7LHfynySO9peWX0P/UIUv7Px/Na
W7sngwko2xW0blRmMgIAUJNMKoBB7TERr9vSognKxIKUXn0QKSNAICczJtzQpIbZ
hpG9RWTJ7EeExdRQgGCT/liPnHWo/DgARfnbPS0L7dFgYeZUrk7ksWUJ9TiY2Ayc
oO0nTchUAScIEUEVGo+1Uip4059ohoJsajXDT73b5yhGNAYMhBiGd501qqL+qOqQ
ijP7DGCTz2eD0C+FdWj91lFSQOHT4JiMKJlMCSEuDLhbENyqqqI1Z8gkM16B7V5t
O0oT9PGZnOVOcJgr6d2Jh/0H2j74AYIMAsEUGLQmAI2+wqzHLXz3YRB2pvfbNPoy
SDF7AcAEEq/Bh5uh4W6HqWkEFGZQCpc0tLynAnm+g2zJxHG4at6Qw2Z6bC1gUqKB
AAg/iIk8H53spyo5MS/4CSnuVlBum0WaSr5DKCZy0XKJxsVxIei/pmA2jH60jDjF
ecI/bB7rfQ8cZvqsowF5uz9xW8MSX6YYiRqO+i1eEXoY5AlgqCPF7QBxTWwYUm3a
NRT2HHlXJHxm+Ho716aTRrOYqEOxCQ9t32olxBmwYaTLGEUVRQsEFcEfZ0D26kkR
5+SRXbthCO3MkmUVnNpUtBIF6hTEOh83dQotffsD3hRuAHDRLlDqRymPD7jw37os
TCO78a4/JsBC2S2jx27CKNVUtkDsHRRxI8S1bRGfP9NGgsGYO9SYZFQXj08w45y3
WoOiMA4yn+l0grJ/Vk5w8S69tDEL8qE8STe2gxfMKZn3UrrlmM7lmSqCEt5Y7x7v
vjVzPje8C6UUWtJFVWH0GdzjBkrFGyiw51yBequInmaBpdz6nRoQNRSfDbvWCK1s
vHomKxZa3/npSuXolyPStu6iSct3CuXxqdAxg6uvWs47LWe8d/fRLcp7ay7HJOWE
mOXfJ8yW1m5djlT01XCQGGEQdfpep5xZW6I77VQ0NXH353IDZbUmjwMnGZsDzpBn
b9jxihgJpMJdonhAyyfwa/ZvFK0uHtrJzmF+bqQsilqCUFJeoLNRHiUMIeaHn5FI
aFrApTzLi8cLov1FTJKPZVHN6Di7F2CT6Gqrz3hbS4iyfPXSD1hKZwFIeXSaZnGS
Zrc8TlVbLEuipi6rn37xskdQGhadt87i2TVrzOGLA9T8jStqZYxmEktTLf8kSxzK
X7sZMzdNOLD4iGyjlA/tvhxgTCusveHsuyTKdcmxEl4c23f07uMAkyvsyxD3nqsc
RQlZZLYVMxnJga+5ytdNQlI3qaLSyhPh88nbqwyxvv4owomC3oHLowkZrT/YWJDl
zGnCGRo0gaPzrdwrf7vJDJCRwRXInjkE0wX96C4EXxnXZHpOtg61Dgylc1159EN9
5o2bvAtYMmukWPkBQ9czoYaHFFd+iPSkCRZW906BodVfb8Bvx0bqgHdezYO720Zx
CI8S60bWWAcQ/OhUXvhfGGJ+xYqSMO4zQWyzPHhJts08nr0j0lBzl8wQhsUvpXV6
4cMbOHprhi9LU7qUJnBYPUPF/9P5/fF7MlbG0H1+FbA4hl2nn1Rt9jYk3bmTG56a
80DizsYGOB+EOWxdg+ulS+yxpC8SAOZ+xXDPlT8pnuBasBPlFY8R1XDV8R1HGUY2
Omw68K6pP7/D3WeUOWrwoWr29v+kEq1yZjPeF+8VR0+pDX7Z076afdVosIhOHmVx
pEgCZ+YkYJ3FKBkUT+etguC4EzL78x0MNhfR6T3NvbNO5p6GNzEOR5FTHSF3eZvf
syUujZWQZCARgmTzLazLTscSeoSQk340tdSQ8fRwCsWN/6rA1fv1H5V7RJn6j0Dg
TXPL38Cej9JeCNajd9VYxIX5nVxuUKlf32lLuEZL/I/rgdkecrUToC8dPzy50+L1
IXSAiz7+UvDcvIFssdLfxvPfSzJHVBYmuWPxN3hcJhyyos/pkTZHmipGmGNmT/8s
fMeXR66P/uo1EKf9CODSwSyXQVTHJdCFuv7UJIREQsYUhzy9JNoaVnwTKlopr2Lp
AEdhf9CIp3TRrzHaN5zMVhGiRgr2XTo5InUEK62OyVpoc+qmWj8nUUmN3zEoqOGk
QXCWfpd4Rh7fvu8hRiwEZol6BcduCMgtX1i1yxOqR1JcKF+ozuUTLnDlfskvUa/Z
8mCb7PMNZ5QLHVDsyRlgxUJ9CAGNw378QzBFWtxCwHVeS+TactE6VZHIxVeUjIAk
ADHUn/vq+LicG2OazcTZx+w0+zGTmJbaFmECQx767alXFg+ZXewKDGKUoO3y0yOc
nj4D0bmC7kL31T2RR1uSxVqOFtU4sQKAhRDWwXKj8UF2jTb6otLdvDzymEFfpOhw
L6WacqMUN0pZx8gDipdYN4nFvAwGYWL6QpTBezqxneSEFXdTHl6r9xlZ+7XZVw3A
jXJ7nWPRYlE9OHTmuRc4VPXZCvCAyp5cqWDxJ5VYpd98bebDVBcs3RnDW8piJOBc
nxEIax9+kgGy1+w/voW8jU1yrlu2iRdcpxqY0CvUt/7Y3348gfPbBvzaNJ9ZlqiU
V4M7RJTKvlSCWSTrbxcfImClIx6zJ2JRWYtMBvIrdPXXvOXCrGBROCKXUVPQXR1+
y8L8Jy2O9+wsipo0zKSCLZivLTn94Em15s4kzCSjLdMaDoas8N2hQJKhaNTPsvP4
yyhJIj/L7mwchKonQHGNfKYFBeDPXVfnGxybjOvPR/QyGSq/I3/8VTscTwOZt0ER
mk3eFXPqbDI8gdGF9AeAqbWHc93fAnkEWuPDloM9pY4A8+GdrfaYuHsv3lcEU20O
1F70CEz8+GRC/CpLZkR5lt11G1NjkibUwsftklmZ0sRECQI2k4xdr5Xwldhqitpz
qs6nGXMD3aXmD+z0zWAHW3msdqDuZw2i5hyN5TwYYPvb1qWWg8yMAmlgHGdxqprX
as7joxQ3FE6g0y2no9dPd4r2oS0Yn/L54E12xpzMv1/V6/gpZjqR/kGnxnJyL68F
UWf0SdJT8ifaz6LChF20bLQHdUQTR1HQv88RLGquyPGl+AP9KP7m7I4nniJeDR+P
Pa/S3lRYRzelu7HctLzlv6CBSYQ5f7ac8jJKtdI1GaXzbBhZy4jWGhLSPdC+RQB8
6qorePekyov0FeLtzdyK/5Tegf8BGijv4fRQCRkExMWyLDCgIXyL1o9b+Ds1gwcA
8kmXfzUHSxt0nkrukA64mezqjMCUCaGA2PnVY+6Qd5KiIVTopdSf11dV0ISdRDOL
qHnQNbWODeTG91DrOddUP6eg1wT0YLx5bYq4XmttkmRaoHRfciYtivapRDKE99xT
UyfEiuJY9zaAB64EJrIrGIh0v7AshQTMhmrwGiO6SqgssZBJv6wHa0BTgi2TmRxe
Bkp7ZQgoXA19QOkakb4O2J4p9aS38092FjHArJ+yGpWUxsX4wtsKoLBC/kIK9Itw
YYIUbkcWej7Cb3y8l5GxVkJ1ldlSBs01G+kQXiy+Yib1P3E+59aRNVY0Ldgn1hV8
f2FgBOGwM1KlWqguBhxKGToPlP0RcbfBOizy7MEBPKvpOyqV4e+EHoBixqqAmR5F
BCvFDDsQIIYioMUWWXbJ/XU4aLfzfKmQa8vo8KSQZ/OzboIbwyLMHPSDZJpMOh2f
xm6r+3FcK+C9TUIf3IObq5AU3chHNCM14OfYL6NsDhHJXFtHa0BH8Hv45WG67QFO
Gi15E2iLWlIXIRCuNuZfW2pbQ0E1nX+ptjtk7+GN9XzAdRjMS3AnM+kR3LS6g9NH
YfpcLoi54IfonRw9BHVLLhNJoFAVONIoctAyP7waD3twvM849sBDe7IUxkB5pWUL
LQ7Pf1S6SgaRJAPIprCqwKPsn4y2jBoWX9mULnCwW8Dr/wBjnOipojeBtKg8aO+J
3hzD9sWE2vNS5C52yezO+0R5dqL5AChA367P2J/BkQ3UwjDuuxe04k+DmbZtGfT+
ZLZjdbTbHomSoYVSwllg1+KbmpIgFTMM+sq5mooBRH/0WJEKVwfMVtka9oGDn+h8
g5o3D5UHj70Xq1jDkW8aQtRMGdrtN/nQ034eSUkVDly1oRdchhqUIL7EdOk5WQLY
aNfptXO4VLF8axrog3j7qqNyjhtT/wi4OSCD+dyVJnSXhnawaMvDmiGbTyLcOWS4
w1nRx2ZoAUikr9esKtmjqY6ZRZvlfDKMWqBKMmOStLaMLPRIyAnZIijocJS59IsB
tjNZylqfClXGRy7Ziyy68fgl4gl91fU93N5csxlUICuFSnUYc4+WEn1g/l37k8JZ
XbQYu0owtIfkOav1f/KmiyYM5SP0a1/YNJnDw55pxLAdpbYg2pcRfmb5R2EApd7+
vYKvz1SAvJ0i5WXQPJYBGhQ061s5p7sEK0IKpJDu6MjK+SJB22KtypZbSSNzDN0w
pWUCIcTLyk43lqtmbY9LqKzR1Kz9zBod52LoqdhMHjGS/4cliNgCpcZ/UuDlLP2b
DbcByZiG78mpBBeU86oFPEeuZBvORXWvYlxPijTb89i+EGCQvLSH2gO6v8bBuI9T
sd2JFhTNK2rFGXSjqGYFACdpnoPPjkhJh3gF4c/zRe/ochRPPySX4c0mfijsxuKp
BmrO8zVptfeW+vpH5QRcYVhQOdfhIAYNowiEATmA1ZpdlDpPq2oS4bxDnQM5Gpjr
lUiIySTJ+JLAbC5chUQknrPvys3hstL+lftUmMf16bvvDzKh5lODxykXMRlYGT9i
Q3BlozU3nj47cPSNpWSotu9lFBXGXVmDioBT6dGUfMYYWxfV8W/QCHKRRjYGP2mW
t7c6TEMJ6e8hkZhghDBlQTxGxkJy4FQd6HtDkPbRfvxt/Oly8VNiw74/75SMqo7F
o/koiNpvXARIL9tzOnU75vhGa+ySRM8qHI+rK4kBC9V3mt8FfjLnTeoXKRff5GAF
xz/61WkRfUNWNQWt4AiNYyChIVPYcVAlKmPpgi3qymF71r6Cl6PEOJimHNdq7S02
7ywk+fHQ/UuexaLD0vHiJ8m69Enlbj2bZZJ5vTyHz307LNm2n8hZIAWAPt0419dW
Fby48EDHOhBuRWrX/I1B1W4i7o6EmpHzDTECxHQDj1Imr4s9hXEszkTFr2q66ocd
JgArdoaoFR3b2WUuvn+MPdxfxyFR2PWiLznKYDcQxymdHvS6kDdG1kj7ZkQAHzuo
eIrteo5MJcnJbJIUdb07ue/GmkUTVK71Qt6VBYVv93w5+L143ng/RlqQAKXWjwvY
PGDAKlhqzOX9R8pNYJ5kiv6bH1Tb01Qs1trw5Qh3f0qrpRhHFQHyaQmnMpvM6omZ
Qrp93/Twto/KWv2kG/qmhIyXgfQrXTUQZ0v9lEGD0LpErYIkNtAQQcAg7VHU+roC
mlV//SKYhnQBE2ORE1U8MYWg6Gl7F2uze0juWbz2QUloBesmpSeLqEH51PeVqPwC
yGnIAPiYspEm9bSC9jSVkuoMqYgUpQqtvNEIg1G1FOp6HWhFwkxbhec5Bj+xkZQm
p1UHpT8OolGAAr4zKjP6MJ3jSh6uqeMpdn65x+Wv6eS1TVKoa1/Ee4DQfd6agjMZ
Vol26hwfH+/mB2Aktde6QhUXiqWNgm9rlycXas6JDQLLDQI4omrk2BLht6FJ2UkY
rjkXAnouVlUojzuoj4zHcAe2L3JBwgw/LWsbISEsbXsN/Ls/sUmY6S+OYYPftK2G
K2fw878MSGpQD7cvoeIA+WwnpEjbYWO9dg6Md0ooMTaQbzdFJ1Qgw7Dy4qH7qqqA
M2FPB4fLHeh+F+GfTQKcG2V22LM0gHcHtFf3Z/nd16nDUVHcSyFtYkrLkUWUINJN
fhKT/UMSsNM8jhocLB2WBs8GZG2NWBqjBFqee3h13r0iBiTcGX5hZ8bwYX9uKPOX
HoV3+ik0OAb5d9tKHiU58k5iBu3ftqbuGI61F9ievdke+s7RA6e7Hs01X9KFnqko
HD++7igvIn/gKwQkCpWLE8W14Ubi0p2v7jH0EyzgRQZSSVfcj1le+57+sSHcAY3Z
6MmR2FDwk/AiRN14XR4JNq8oO85Rqq2yKnkYm+mziH3uurOw0Qbxke2zWZPSyzg+
einvkpgrggHrSt4Cd9ai5fnq3dL42tS8ZQ7EunOWHcWLbm1hcWnHhO1q2rJCHvw6
fKqeNlAuC/74p+hcProj298JQt1ovc3IdzklHWzXWz17pkIPKasa0mAc5KTPH479
d3xUjO/lVMkK1YT0SSY/ZXJmE1RoDVvu3g40FLm3cV3ZfJc3LoG7i7QuROtZOXJB
qQiLe0MPEBMyK/2FYehBOhI8u0PPoK7ObOM7uTVOmgaJKhgHkATHW1gRvTsA7QaG
0WOU67QCBp2RIobX8fgkKS8Hg6Y8F0EvF3RWslHG0oRtAgDtvWTzA3Q01y3rQgVQ
GLFEmzZNx5VrMdubNOm72RnenZBd+qbN2XAOt5J8LqdA7Isuwyc/gp7RafIt/YFK
7I6aaXDM7WPEsxIyggiL/nj78g41/+FGBiFGKcFFvLBduObdHr0WERG7u6AHOeM/
5eAHu6gIlp29S2r2TF9x9LaPqHdW7qc9sLfkufcgZLNSOo0f9tOZ4axlj8RslwWt
+vwfAo+W6jmxVHWDjj/ovnU6hf3P0T5Bq9Rmarq3L9qlBwYTnjz5YXpWsYujI8ZA
z5+Ks+6QzZ9pl4Bx8vvRBaAi106MIyZ+aCaAfRpmqskuKkDmP0ZSG2N6B8ZMfft0
N+192bzCMOGGYSyHaRDRawoQC6UK0I25Svj1oTFcqWDpL5oBhLkuYQfwUrtVK5AA
fPGE5rLYa3MoRyne95Z4cqn3hbqxlVjiYylkbjDwuAio6vwDzToKaxV/+d+yC3o1
VrWUu30yhl74J1N5VUsCSifBrLe4uk5DHGNUK4llMwhdodX22U1Q4HIDQfFGJRMH
JGElgs8RyFNEf2q2K39HNMYLgFkQvks6dDTs4xCoy7c3ELbMmXBTNngJR8/lWX2R
Oj52qyOxcZgknP7VtIBzgv+Hh0Vn6Ztswxu1yDTPp5LE0l8g7C1Bvsf23+Scx4Y6
5oPdXekzsgi8U7MB4HYK5jXt0zavGXaTsaGcPPWBm4qkM7y/HP1RAC+cVD3iSkOr
NFoAi54dZEfPRYtI8JZ/tP76WtQPifA8EjyXiUYXf5NEO0SGUxVAKdebSgByQRu8
Ta8Rxp1RnYdxyzRezUJ7wqE/iCo+4OVFEdVsVPUzDNRR+2fPWzRVnlLwbNcdzwNm
RrANK50MOb0Uih1cc3IArGzQl/QvDRhlyoJeFVUQLdSQUISGkqo4q3Li9oBNjVj6
izvD9WaS0GckaxdDJquHiiiuHBqnC87Nvl2W5f3TD7U0zlaImDZp0/0eU4PtrWPN
JOVjrR3uAEmm9lLQqrPZlVoeP4Uabu1DpNJU/26XuNqXffGCcEMdsSIeCl/qu25g
MqRrwnaVR7gXSA0hZCxPAPxc9wNvJfAuCqY2mwj7RtrTUJmQiYjY6rJ7r6M1jAeh
QPFrwmPPq47R9AOjFHcTfKE6Sjtp3G4R7mbpzFjky/q3V/o3i0JLYhwx4JX5Jlhk
sevIomA9xst1mVbmeIeSM+45jzx70KWoTtlXjmpZqdEuwoUFUtBOU26onRXX8w5T
Ygl5LR6d3Uf4XlRVUFwui5aUr1weyjulZe7iALCterRZ0qXUnvH3nJ2He99Ca9IB
gLn36e0VIRJCMCtTO60kRrGKP58M8dSjA6NVT7lblbr1480RNDfNiFdki4h5Pnya
vGGUo3vmzAc0iHKVTBsV6n452dJtsxFXaSA+vW7v+sgjPc7y2XWfdWl3e47eiBhb
R3cN/pUagVbLlxevcthF4dVHIiAuIOByBiWbxYFJ7H8HC+BUrR1ZwCbsfaUNNtu3
kAdDkw4MnRdtl0qYZrZZzfWs78wORN68D6G2XM9Zcc77Xk5guJcaSCyW9XJtHaFm
BsGl0ZLOQuGsWO/Xy1eUnVhiFd5fJ5mB204O5hvmoDU1qI6JtxiO5sXwU8Atzx2q
n6A1qGZMchACHOzGO9kY1ZAaFdQeyTrBA98z/FRECDQ+FZ74WSciq3SWfqZGvdbm
0enPHhCQzfI8iYldC2QS0b/okVlzXfTlleHGVWw9q3ERHcWTINH1rXXseBjt5lZC
2JOL35GQfCsf9ojGEfAxkfHVom7Z2xHZzZ0+23uLJNrzZMFCnb7JmmDjVj0TU4j7
wErCE3y5RVeB0A7yqQGYgQWHrXYBh4hO9IvRr94doHeCtPm5IjnuXoWuSATooh76
+pEvNRSPc+MHvsv+Lh4ta8MwK7V5VKSErVLPmWCJv4KDJECRvFYq51cvQQF/E+k7
Dfg6IbOuEvAlFNgQZyS5IHxb80oHSS+elU4KL8ObNCZAm0WxZmymNT+Pn/oypxUI
TR8s7WzM9pVSmS65zt9oMTRe/sTQ1WxYa39AXaBPzN/9tojF+kdHls4Lv1CRsWf5
Oo6KIcSWK44OaZQWNv8FOh4KtIaJr6RA0MHpNjvKATwIdGJohQlrQ/+fsbcsRXY2
MvVkq/IyrLdk/XHwpHdn5ega+WG7/2jws84btzy3GWesFiTKF0Isd+2c0XH2Hh/s
Tmr6FQ48BRKP3boleNVWwrwCFcYAXF1/OmBSqe5EQ2T/2KO0RDvp3nh355p7sFEv
R2ZOd6S8mPVeYrb9fie2tSIATiMIpMKl/OnT1w319eZNmG4FBZyey7Ie7khTOpfY
krb9YxyvYEekP1ro78wfYZk+7lOETRzseSjOh7oltB4lJBuUMPl1fTycHjSGoQnu
30cCB6PtZerOMJjQaI12hmRFlPgbB7EvGO0dQivc5jkd0FxrI0W1TdGu8Cu1vQcN
PjazEBQ6tjZnDoH7eGmKCx5YczJOXt1MfnHHZX5gj94U5JilgEDE3W+coJDFXQTj
CcL51q7tesH+qvUrByyJk7JvWAbikZstiP8n2gP1v4BwYqBrjURdVHe7jtIKFbbF
jeev5hEOJumQkeUuSm9E0D7A7FXahYOGt8idcJoZc4dGeoxgZ8XldlNDC2HWTmXB
Spu0I5ngaItsO9PW9Kc5TIMecyK8BN4gdhT06MWHkCV65dnQCuIclNCHiU+2X3Wu
TFeMvhBoYZb/uV7JDVL4j4oG9I6v3qGNNYeSToiC2nQdnMDDI5VBZIMqT9C+A3dA
U2lxHP3uk62L/qR/RbU5vdurfjxUNdnfMNhmZsmCpJQCWx6zOlxJxEEOGmpKWc4O
nofvndgsU9j1uGug+qo7pAwZXLHy+lQjjNQYgt9mUWG8xTvBaNAO7FPLGJv4A0bh
VQ2sOnlI788CF26pk0LgSpxJ/fK6xucLM9TpIX31pe3atYGIoQQbJqoAnfaqi1eJ
vJJVc7O2KLBWGglMbhzjB5OuM8Xb/6xolCz7eyGQAx7snfWHGYlVO8qFA5Z+sPvl
oOVBDPqD4ohWevtHaMESG2YsEseOveKer4yv7KmSh0gzigtC6uYCUrRma53Eef/F
1iqR3ZY/6ZbwXl7tW9sydSCsYSzasrNJCCPiNLsp7ImOzvCXRCACCXgMLNAA6fFM
FaxRDBiexT0NxhE8JQolgzOMNnv2HFQ/pTaoS4KdFj3D47F1wuYRgo24vOetSRqc
OwaeQzvPRrvgIOoKzxZb7Z7p04sYNR5Iiz2Q6P4W3dJ621lpBFx6LOycNAmo5RCB
Ko2fPFqi2UTBOwrrCr6iEt6eshfNHLwAOhcOcM8UXbzDh6ODNPAj5BnBE+ObhPEw
vZru0j8HvKDqfDd6x9jbviEHpHSX4kxq42m88LCuA6mvN1ICutKlQ29R6WCjuNnw
zOzCpkgt1RNw7KvWARGxVfXULvRxRVRQvJq1rOS7fd5osxmVyUZBFoCxMdchpsdN
oo06ryrqcAw2Em3mnAm7wgifXT+cW7hYi4Gqvq8qI759STN0o+ri3DA2/UYdNfU4
UkI7YOA1TmsymKV2BF/mrLYMz5HOiBfCh388tDwDlj1vSUBuHFz+h8zYLLGo/jGh
NAzWPa8elu8EuredPe6IDELUMZrg7Yb7rSfGIhx6wK81u0if5jn4AOHpVM2XKWIP
BEkBq7pYAFyR/Cbnyngz0Uzo8dh3Ud7N2Tce++1vMYn8P2xzkUoJOOluAlMnh+/z
nyhTIxUVxn7zU8Mql4wKk/3OUlLFjPBg/N1PWRxlRjn+rNSBbiRrC3AANgfdbNfT
Oj1cKYgBtDjl4HXmJGzU8lgJ3GvctZ3EWUbCQy+kA71zv9QrIVKBH4MUBwFQjWsx
IdcobW2KdIxwXzto4K1NFq7hecxIqAMq/b/e58NEp3K3eJd8y9mCtByK+J2M9rbz
E9dUKrN8lfPo7NFWbz26oQ7u3l5iJ/VYW3gN32pY0alSP4XSxBN9mdxoJ2jBZQZR
FjBsTUXehi+ggB+w4z6lDF7GMgL+V2//yykoWoRg1+P5L16hJ/is+CG5BbgIkLH3
fIbmzAXLqv8SaxlBbQ6qGrEKFg8ugVI6hmXXzHqTX4tC4WUOBMjf9V/4m6PTC+0R
yj6Ft0/7mSLykYxBzi2UppDadcIY5PXkbaYaPnZtsJuT9f7QPxureQt1NZYy5LJy
bnweVP0UYzqkoRXiovWE2RIkjF+o8TLk3q/Pgr4kHQbIVG0SosBN5P6yTQ9k/nrq
lAJjbwFlTgZlhe5fe3I+wb2HY/WsaVJW2sG/hOp2tQyhgWPagLjhqhUWQVW4GNX5
bb1SyA9lNjycNfkOG86LZCFX30v/psAfmdMjp8PONs40IXYTpuSW4E4Ev/T3J5Oq
N7Z67TQeDxW/uW7ukrgLxOSZwkkzH5uEyYlbk12vfs4=
`protect END_PROTECTED
