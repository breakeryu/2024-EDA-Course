`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSSc1lcMSgeBsA2ARPq8wEQfePCiKrb+/QCF+/U2HVQVBKOgKmgfBIBJlclxZH0G
8Rco3KlIsvLHKuNQFUpj6UUVkQ/N/FkMrQIOFqaLGy6zVDVWQBg/jYHSFQWMXUMX
LEcdA1CX3wwSWzXEKNf3KytlDGlWlTJFX/advVTvT0pW6v1nSU7/1aZphOdSFIix
YTfZnSxjyS6K4bfhUcb4Ky1/J4Ca1qQzeqXaXqF63JG55PFHrUw9fB7EW6i04Ag3
wsiP3cww8zoIl5+9uSi8uwOSIbVyv/nDiPnkwMlVjcscmIS7PDFUgcre0da2PeZe
DbLL/h4grZbrzbEB2uBnryZDwoydYlxGBxpZdyyB0Wc9gnKgVmsfj+Aef7/f87g8
AJUBw1/YozHlYCSM+3O5InecoZZDgAkuOqux5WB7qCvr5fIkHiZ9gZv54oA7nAT/
rMpShvKJ+4QLQpZH3p+wbdVWSYZS0nbsp/kf1SILzrECGafupLSs4UgQqrRGMwpH
jIgJfMTXhJWqCTEcjMCd42C3NXAHEFXqGWSllrW8USC6yUM6Uu/jL4KOBqdcRYG0
KUxKkeVT0KR9PMCrzQXI07SJpTvWWqon/M3fJNPfnGerd/FvirkK9S98mJgKeEOc
gMG3Tsrc6w24OTrtuTggfKf8zX+zP5PY6rLIwcEZwpup5T6QeCAYye1LSYgJ7Bnb
Rf7r7za4ulqgnYYRxBDgG02GEfV/m43PO1o48GhZqMSKEl6wXYyjaP8q7ll90S7S
1WxpQMs4hItwUKgGIzuCUsJkVTdUVt4W/QKf+b4MogHBum8DPLlwwveECojmDdN9
zbQvIQ2yyNwXdOm7IgrBqLPz0gj7Am55htXiiqTI//Rjb2Z1epyQvdH4lmEehD0r
DU1g3gtpt34jYN1tJVhUZ1P6ncPDcO7K1g25lvF6COKvwXZu1eOdsSoGW+nPXeLA
6Q/l2WFA91LprIrat1oAVyllIqC0igWxW8/WkqbnBeMz34wHpl4YkqBXu4IPW2Ew
pWKeG1F+VcXo75XodU/CL7vEBwAhRdxyTkLY8PkI7a20EyzEo6XYcYCiPvcgesK0
ah/Xqg6e3UVCqxOHMbgNVr7q9NQPQq8b8VpOc29kefqIQeNXQaEjvSj6djzi7lbn
Pi5Wwosozw95ZWE9MEc2gnlUWOMZ21nTCU9A0YtLI2Qw9FWOA71ZG640KIghvVEU
z9Jz2laGx0d62F98SwFnKynbDyOYblWG7oQs/x/czDCPl+F+6mIcSbu+42cHytMl
fcOmevQh+gjz4rPCHkHwWavNqxJxKEzocBwkdgk1DkmOtE9O8q3xER7tThCmllLD
mpOoUnMcES/VDi71ilXezsjq1Y6mC0QF17Ns6u/ZdKuzPuK6yjpxh1R4SW9g7TlR
uFysBCvSIF/Kt6fiZAG15p3Cr9x9lVBxGOPAAtMegjQZL6hez6OhEpTZlb6C5kIB
B5Izwz3o32Qe2HsBREvUCCitmyemk8i/xLT5T2XesK+1ioacI8zAI1LDaxNEGRSp
xTkBbpefwBNTvq5yzcWxY2frz9Gyl1fu2njSteoUV/znnfo2QfwgAE5A5fD0+6yD
Bx4Kivyrm20H3/XCi13EtTNilwYGAXM6HWn52EXphfusMf+Pp8FPmSPmI5OUirro
3xJ5hdRrCH2F2o/vWV9ixkYOmRsdijkDmkp+94mUYhM/6ZcXqgoEr/LyYAIx3fZJ
vt+Hb6qxV+doDKekOjL9+1tzDzaDYUkrAsxh2jujbGUe6Zkref83hlAhK3O9pOgF
IYDbFRZEpeVn1JJRi+Uqb/7gbLFb6bYCHhwr9Co2eJTHIz6aqhoqGcrwlpHRhwmR
mHmoZBaN1dvDP/YUm2Tkv/CdFI4uNJwr/nUfKsH0+sonB9nu88CSFeqdocJkiPM5
RUNHD61RZCjcwo4vMUvloJf8zR/3KeQ6NCASxG8sJ0PZXWyr47+YhmVqH9tq7vtN
zR5vbUkX9337SZ2wAM4rTTvmsgobLD7qswv+A9+WTH0pm6JqyVzEw4IsgSHMznTj
L/AmjM+iiSmLmL1FsRuN4+CNIhqHT1JBYV801pymNOnu/ybTW6be6pf3idyQsbrc
14tMIvh2UG9l0yybyLBWE6w42Ml2LmEZZK4GgwxlLRoBtzHSUx+JqrHd7q+KInie
91iLJhfaZeThAAkH/LCkF7WuvNRljDGhbxjm294lJq2GQKGIfpZPRZa4MOqDBVJ3
wFhIkvobfXxIkBBphMhd2kwPppn79OlVruwe+alF0UaDbLnyvdJ8DNJwk8+GIPyY
txbuBUMUJPHt6wzUeBM7oZ5DOphDLGo/MoXx/8rcpX3JNkXrKMnXUQGyrIl/F8Up
rWU2GZUdT2DcIzr1ttfho70q7/oPlcJw2SWd0+rRkWE3Wg5LEl272itnGzYliEhy
kwZhxpXWaiZnFyslQLLmhG5TJ6AeBLA2tTXQevneqekwGX+huJNLqnQWlnOSmbdP
MdrawkP1oAqVPcQ0289zuhTXxUismiLZBnhBT7+tQkSCXVKBpQX9ouEBTRGizdyx
YphJlwn944g2fe5bfv+U2Vyzt/ySJjihv9lcQZMwWgvRA0vdqZQxQQvyHbnigoRo
TZUZkvQmkd/iiOZ7xSwTqn7RX29di20+3qy5CkI+cR1xWl1IyjHSRg5c8Kl30ceh
+rJiyiJ4ddC4MNVM48ryEleyAIAARiLSNQjYjl2mUvRdwVIh8cu7aMja0CzEQmdT
4vGHxOUoNzO9zPpIuU62nw7N+zpsZ9iZoXNMB8NrMbi/v/8FhnVxJcizQ2NaOMfI
NxXCEkvQrtE0xF7f4en9G1fTmBEat0vLxuc4hiiiEBZ1VMfk0fZa2d7gaOucCfrZ
ruUsmPTg8atVO329nBynmaS7EPPclD/iTBpPvMedNA4D5SYEH5PMEyS1vUIS0AmD
BQflCNTsljgPwyDL1/ZyvT2fDQwOO5ua05s7hDy35OV2K3D7v6KtOp9vvSGVY6iN
DHIKQRJ+cZwHg3jzvaJFezaXeHR4jt6BHrS+KPqXfVuQ6xht8ZlnFlrQKct055oX
UU8UmlATpS+0acYuPSSCIYOsVUo6eb2BD0dmIuxS+thF/Lv+1o9z3/7A/SN+F7EI
uT67NUpfXT89zbwqisMoJ+elFO/X/Kz+jJGxnIJc9NbRZH8HUtNrdpEty9bk69cC
i+l9DUFXj7qwuaFcSXJVUacr2sVycB8tFwiQh4LUaSyvNtFoX5s0v0RMBbc69imc
fa4N2N06L/4RhoQHZZk/situI3uV+EBUtNJGhy12wqEJpOmIR8iyd9hrBE4ORvGG
VxpWL0zm1nNhkhsAXptkBinI5cu49Pd646XrQhY3MlDOHhewe2iHicDlPSbERRxX
wJoFB3L2UA8xIGN2rEixJZyeUH+19/G2QE5v8slA/jZJo4NGea1Re4t8wyAKdQqy
9GUQJoPzPj0JjNvBFWiqP4yxLGVj0ESXcSl1pZdVcvrDNPeE8/AjzAKWtRbmzmzu
b+5FAYn0nHJfLMS0GAZpyYSTSbJwTAU7gFg6RtK05Pq7mEww/PWiFloqguWd5tZ1
8LX1QGfqMjXqpknkmBmCXbugKZG0/uhE5KhEVNE1qhhXsk+TxuJdSIJxgV6es/WA
7utZoZcK0wg9I1ckxx11Eyr9fp8l2sbRKIo/mhy0maQ03Jz8/wkeBOQOtY2qKkKK
sS1epDGRhxf+6frVUUc8l+OPMzsiv49nvamW1oCZNkkU5wssU12r/duJF1zQJKEF
bhNI3oMTAjCqE4L796A4vNb//pRq85ATnQ4WltH+GhZMxCQJGCiRZQPZd661vYHU
FUXCwTunpLqQFV1v3UiWtp+a6b5oaUQHXE0HH8JKiQFUvRw1yvphIk7J3+ybDAkC
4CiRjZjuwHtoRpdQTKk1cqt2OyzPybODe4t7HXOQjlUPpi7SfzObEqpwKaclFQMK
rh/TCyaYv2xVeUAyNws3KymDwR40wpuFkESXR7lwE1MI3UoaA886H0tsCr3dI1fL
lX0JThP7VU7ZpQ3k3bMTJ7V6q4ahtRyyW4PDaMvCF9FC46amAWjD9drFWLu4pnnH
XwX8IKUUR6oFdK/7s0P2elTMdf+o+WLZxZpLEAGZxF2STDlqMcR3e3vAIGwlmE0O
XIM/PZu4dQblOUSL6wbSCu77AgU3aBdT1ASsukB4E1HL7W2XS8pKmJpN30aiYXH9
bCYZhuBORhTxkQIvoHgdQKMyjwcyHrYtVXkDDWWiIjG6najA7XUr9Jwf4ZOGZ0bE
VtifvM1ENXJmGwr5H4bQg1iaeJ5LCZMnOrZ62Iss/kCOy8/HsYVvlmXcHFvOhYLr
c5JRJ29dZKkR6WpilAM3dVf065IW0LwOJxKEF+AxuaFL5miEESb7Haq7Zxu5vvi6
2q+nc+lLVdS8P4f8VnzCPmEFveS2BoVr93CP/M/VF6hY3Mo6k3sXm3p1GUspII8O
ZdWaGO4xxsNDGoKCxzn8kApJ3pNE+UCYiuEfAMmd7G8LI34dK+jWR0L442fPOvSW
87y1xSoVGsrvQpwkz9BB/w2cfB9hk/oRWKY+TeFcI9U9CPjejwEn+SggIYVSyLsp
2BqW8bFU7kMIgJAJJi6mUx1cZtxGnhRyapsgPsPjHQsF/arztC83UvnIBZuCpCba
vjHkHp9OdSP7i43dhvYX0wjNFFa5E6GcPf7FghYiXmpujKUUMRd16WyigY9TJhbp
yFsElTIcQdogtnUmWhgm+TAG/Zj3NDdD4ELeu8c1ouwfVlJdryqSjFSgnwyiI/9y
Wsw3uvzpvSPxcvWKjWRxOus3t22oRjFlT2sFP4Z/jNcyS7NcCoarjXSDqmxx/IA6
LetPI5tG+BF/0h33Clb71hHG/0/blHBQCkTdc8jz3o4UOBHRir3goyVXIywAGTrE
rd1GUCUBmKY6kt4kIitQT1eRFUQ2jEqAoZR7iB3NFDFDfQpLR++DyDRku+6PgTZ1
F5+FHl2+OhQ/bCe7gXGYHAbnvW76PUzj4b4neXnB28IvIja7JpF0B5SyUUeTPM/r
OczLfKsTDAQUSZrNddeef0N+7fOw4JgjLndm2RKMz4GrPR1Q4WMshkPASKaQV1by
Yf99DROvEGbCO8ilwXN7d0l/1izHM3o8y9zmJ/5IYtXk5JlfXX/6RlTvzGJkcZx1
lB9V701JE8pqwR2YF5TvBx1LKQ5Z8rN2RlgRvfL+nzVKR/lHLQW9B3YYx7uq2uuw
eXq8mx8Y+2TmOTiSkcL12lP+GGL4Xc8OczrTEuLLtPA78JVZzzJFUZXEsYj0y86a
ifBv/t3N7FQ88NyL3P2gUeRetU/CdHvPcPC4uM0h62Xq3Zkes0GDzud0hmb0zdli
flPb0hqWezfz8FxblSaUt04gNegtcj2/zMinM2Sw/1L12m/HORQlNkMu4amob/TV
jYWBCwONIdvpa9cCGTAizboqWU24RrvupFslpxFh/OWHpTCOuDzIQE6mQaArpZwz
1E/zB0gi5he1DQkg4S96ai8Ed+uNNT1Wsjg4KCGhUhrCg3TGRuJkJwt4CTzsuWV5
mMn70Fw/A8KK6P0RXm2Nl8PGRkCpKSXsBUtVmW9vGmPP/hPuSOv/tytoEINec8TX
z1nP6pPUHBg14UKEVLEJ/qKWZBLg9Crwy07xaN+Mey+R95Wzm3w4TK6JH9bRluCK
7nbG2ALfi3pVbsFGeZQMjWBqi5oKQHRQ3i6knvQCCHGxf+KKD3nGQN4XWfnZr1PO
IYZVEX4mX03FicdJnUEABYpARxdKbkyzQPrsSlV+t4CbL/zpB6Er5EpzXuL+i/o7
zP0pXFpy0TGPum7kMozsfME/149dk/O8Z3Tdg0YRfYjJR04V9xgM59Wgye6HtIjx
NovUoKh7rulffg/SjRDsZU2tJKCLBiFpouSo+5l0Ju3QCf9vTWbZu1i7EeIl+Wk7
IrICB6cE1bcu53S17MfRrsiqBzXRp4C1CkaWr47gk0cXOsE7kylKXXvVZw/mCYQE
+rba6UccWDIL2SlEe2dVei2lBTqhFKH+Sqp104SVo/QSGd9xSCfXBEZzZISWsofU
+Xqmr3F8RXKyYiAm/YCEwdk5y2FtVZMu1Dr/hd35UKFTcWRO1Sl71PKVGAa3Iu91
grJ1rrsFiQOnGj0L8IvgP4vNjsdAIBAZiywWyx2e7dXBvxU8P1aln1lPTivcaJPN
W8vMkvxrNAT4R6y1UVLpvUx7OOAb4KVV9wMW1El7NcG5noW5XVCP/Q0AzUhfhlIX
zuZXia+diDTdmpPKjKGMT1I8k3S6Po1asnFSUpyM7D/4t/Hc5eSv1dzm9i/8l19t
78oKJUt9iQRgzqCFZfTHLje/qtpLSqjsJYg8Rx1SESkUzAuUxRUwrsNIrFSHPXzj
UK54K0FTLfM+RAXUuakKYwvg82SeWjRts90bH6l53K+bXqDSvfGJ1V4sZ9yURyW4
od2gSyq+sP0/aDJhJ5bg68klNTZjgRpoIF+p0cyoy3pyQPjBvBJaMFTxQ8fBXqOv
HDytyFsBTSAJBT1GE44Aok9LYdaxv72d77IbCtI6XbZu9Zz7QAzUR+qn+fMI+o7P
8iIcS1VbMPJdAR8CBPkxe+NuC4GIZEJcJoWD513xziTV1FwJ3LZx2ZDPlENv51Nn
ueRe0ZK4rVmzwInohao39fj8b4RuS5DKQk21zqBXM8eFpsJSTAuvaBRJfa7BsYP0
SdDSZz+xhKeJmJuhKSw1+/s9d3rwQg9Q672qM7gYcOn48KMNsnTcFV5egU2tQDCp
6wyF1t+uHCG/RxpepRKQcLvoBpJ2iA2fUvbZ3bUsoAaQkrsjGy3TEfNOfQIPAUDG
SwghNCzkS8fcVW/jGBUH9DuVGn2D1aqLVefNZw6hCJ/bxSL5goVaq5V/J1drZWc8
CUybVnj5s8DHZ1e9y7n8wom3iL5AdfwQmcmpIdXewanoW1FW/JeA6vX5M7/LREjs
YIO6rf9UEWVMWR/PY8dySA577Lkybv0Elg9rRZ9mjaqPmc4O+80ErICaqV5bIS9T
Yc8l+dVcdr8tDZK4sjjAAROSeBLtcyV5Kvrr1Tikx18S8wcDPLy6dYc0yYjyJp93
O/lgp8P0hVCJooSn5PbWKXnZZF9RZrq5uITYba0cgJJLP04G6/lg9Pv0RQw2gsU3
iINCKlczPCzAHN7YbnYfkF3nMsiXla9KiZ4U09ZgEmepoBkg2Lnw7OqauUGoTvmV
1nUbv8tORXkdTlnKGnH82I0WJbsHbj9HP+HR3vYzscUwMkHPY2VNJ0PC7+azw3ho
e8QKuxDuOAEtJBWhv1XzH2T2zB9bn/YpM596Dj92EHlzA+gjmymtFEK8djLHNvl5
m2p3ist7lW4RWSxNZPAO8OM+5Puac/tbo1vS/MIJh4QbysmiHwcvvLd7gJrLyROQ
t3+nn8XnmnN6mf7ugftvvDc4IGLGbwr6pJXTlb4xkYUO/xcfu/leGh9ztQb8IOWS
mFB/YdfOsNWFztfsxUnrewqnzY8SUFbeAKrsQcxFOrlDsxHrfXeUfegZlwOdnzZP
67dFTL0GO5eeAuWMlE0MeIODAFXc7A9I2BnhErqUeK/B15cXwodi0HTd0b35EVf1
DEIiq4nDLlKL/HrgvZY81Xa8CWU92eGPERdBTfqrRlntQA9s8BOOali8+B98baT4
Hgq09FC5bad3TKtfc5fmHpjpA5aE2Q1+l0wnDlCWx6Svl+LvPmU/nzoFIvFDijyg
eFHj9CBeQR0lvv3HSTRZsoQnV4bUM/587zo16rGcdTYTuEUL4lzz8AhU9iNXmpT8
l3pQHTk0XbncsLRrC2l7CNowfV+LEx8zmnsmuANY1SzUpIk069C0C7uS9X64uve4
zwxQ0ytM6d013qDOjC02w80CPjLpgQNvlDyDWMIFaaNrMqvDiAUdNA/RHye+Fx7B
VS3aKtaGHUPnQPf+FK3L+ysFBiIAi5d6NOTaGWL0485TMacjhOhpw08pHKF5vV8E
ccbrcgAabogW/wpQz6xAuKYiNbuXU49crwcGmhCrMGUgSx2FClNE9Pq3jTKSqgVx
yItS5jbmTTWQu1CHjV8gAbKsOT9pnTC7W8klPwuWogG/Uf5fseNEMbCoGed6P537
ZsWR5zhaFe/aDkkbMS9wCME1JU53/iGm5CoHpdrZeS7Q00ZPHnTQpwPKxaFWDekh
L4eNDK5n49iPESibVBM4s8FQgJ7BdkfPVMGEAyGpIVWVHumQpVZ7hKKMwsiGBqdO
EpnRz6w8ckH3/CUoOZOQ9PIPROg2eORAGWwSCmlgJdekX+ZCRWZcFPyk2cGnjXWn
n8QeVDWtZKWwItp991Js8akYmqMGTmJd7AGSnvTpiySWn5DvRyH2ZZcB72e9r9P2
OXwBYyFLhNqWHZqOzQ044sPWBG5duI3XB2m/ItO+XwE7w8pEEKsIW8UFe81QsP/a
XSrz2Zn1NjTWDAqSuOanzL6BGwp+xypDE2miB7ZXn9XjFuoQ0ltnbdbbtSROgZlO
6Sq4LZVav83owFi5OMs09YAvHRznRRdf8KX142X1dANQdWchFA+et+GHAn0dqx88
zxMmn12UGA8hlddkmjsyTneJlSZyIu5g+B6tGwbFsAthKjB9kkilJfJAml4Q1OSN
e5S6xAtBJdmQOscfaJ1khWOGlEpD8ooOXVDFLsBtI3vKPdcYoY5u4GytkTJ1ixDs
OXcYfQ+vqKjGc7asa+6IA+wpB2ANfiB8Ss65ZrI39mu6UFWWOkdrHvMNidsEhLRU
anr7Xaj+hNnwyVsbB9s7rn0Ui1r83wc0HXBUXsRp1PudWevM28XhvHHGmSgVuqlU
LXrc7ebC+O6PHWnqOY2MHf1rDv7+vcHYv6WDp/cgOp954M7jwmE4Xgd1CicbHZUq
zgIUsEx0zhI6WxTCNFKBvU1aEa9jVoPmvup4o3XC0FUngb8eMx+WMuwG4J0BK3XF
f8As/UrFJhbEvRz9evrpB6wFVCVCRBh8T2A4H0Uwog9ZqT8iSnKUUVW+QeqPrxiH
yfop7arHbk55+elWAWS1PJZnJlORBEoFS+gAVzLDNGnW8w5qv40Y9U7HQwTm3QTb
Q5Nt9RhY7JRDpbaGtQswsFSoiEstINK7iSRYkhPS3Yw8g8YjV3SOdBuWYcxyCbUX
hoKHSp+uiH4puFbpkFD+Af1b1J36GMzRpOHpnkFTXwArQ3uxQ1sM02voSOrqLmIM
mj83Gi/sN+r3N5hi2XEjMydeChworxpUAOv0KU9IQMIgdEST7WdrhuCZaWzkHh3s
l2Ov9MiTDpUjI9H+MGKltKqAHThyeXRBEhbHk0DWfp8+fE65pyjE5dX+1Pef9/mx
bbjP8IXyYxBi//ACTYX/r7iUconaM5c23vpXeqOZRcLlXRZoBJEzBL3lk+xLkXzg
/CQxMTwxBDGjvVlTdj0187RTJl6b7q5FoubaQWt8C+KpvGqzL5KJBYxj1ggNkC0E
SCdigD4NtZ0r1h49DxirZv3uboR8kuSj1uZisCsFinD5mSlcQ6kSVJZjSCpqoJfT
DgocutxZjHYOmM/sr+8Q8IH+m7RcvE492c9ebo8sTU4O1TJTak4wbNA4pk6obZ9l
5449GS3E9+bWh802I9Lg4mKwlbkbQ5ZaCHqVeNJY69IuG6nCdeOAEGDlruakdaWV
lo94kJa2PKOzYw2qsnjaQCv1DTKNl6a47egMGSV+V3fb1/863cPS3iF3nOtYNT2k
zZSoq15f4l+fiUnj9W5WlVZm/mstlbgpwyv9a0X7gg+b6UT6yQ8uCXlu0LDgEq31
c16KFYLGClrczw3zJocywW3KiyLnO7gSNop1g9tq06dR5Qf8Yma3fVVsSC7GSuFS
jQNDA/FNiNPFPfuIgBsUA3SiLQI1bY6aXxIZSBAjNZrB6m8uTq6k3OZcvMAIErwW
IKh24zDKCeDwaOYf+gXCn6y8+1PVhXdx/R22ZQzQQrFjSdhYMZuk+Wd1nyQiunlf
rnIVrAE06/o1WtiVfwDnDPCxX/8pKEVAQHfAY1a90sjxsJ6u9NaLgmQmuWNgBiC+
RfJ2CvSq4hUQf3sP+4jL6N9u5qdRn8gdoLPKfl5YtewfXMmhzddu4a/VmPL3VOrI
/dys6QMqbscT0K/OFet4MTuLvQNa23BkKw6vv4x3QXOVDsv7kTQLv2TUnIzNJAbv
Wl6pvNOOWctXZeJY2HPLZ5A84p649sqWUjb8e/GJLKEcMR7RmElV1ub2G3w5N41E
V/HMn6/2AzpLmxVuTWt9yO+WaqwpeWlk85WeLXKQhcBnMU2YK3KKuFyb7lQKGg4G
bCQrsycsDEQffAEyvxcN7zIZ9ot+cZkUMkKK0k7HaCE1YiYqrTK2+71HxHeYKcNg
kMsL+kJ1rawZKYELMgDFlE9ttnMVviFmc+wu7pQL2n+PRLb6FSgRwaKmKnRJs3Dm
DelBfhdQjRMLlDjY2cYP/1/Pxa16/MEJYGwtEKl5FBDxkaFuq3YYq/fnW42mziFH
zU9LSmSOXvwgoxhwLkrOwt6mZgU0Se9BGgQ6x5jgGts13QGFJCsnR3xo22shfo/1
aKH3SGvDmGocQsLMikxQZkhfE8d8+oqHehhuiJqxn9/8CN6lH2I91J5AfB3bviwo
oTnKqgp1QN7dVAFqPCWpnoOl9rOoNzQfE0nyF49zb6edW9Tdm2IUJ/+poSeZ3T09
jNN97tNzjnGwgDOQW5Ubj+U5fwR1WDTKxilxTdeuTEQCKZQ/+AhS1A+3f7FZ8WJX
naTFBWYNn28YlPWectHDbgtAsBwDe48qLT1fy/UB5xB72y8vbdYAtrmFrGZSkwEH
Xtt8mP892A/rYrPuksSF/IuDGUtDtBLnoyTV1Di4Bu1AVaSCwI4GmihQ+CH53m20
saNB/Ots89QIO5sOBN08r1uvlpKvCXic20nMqr3b/iYanVNaDNBnyTrAoAyZjiDu
j6uJJ+eybsKOV+4tz/nWbX+qrarwOkkW8qdJcaQzmwiOWl8lBgbBjF5vOyWuCU8x
ITw90i1IQIvoXieu5SBg4EvqV8l5tAhZDqkjtd5n5cvzYDuuALY2daMfNBEgqrXt
fjlb3NYsbg5XI8aOTq3hr/R8J37/pCSm06ETyMF9oqbaTJeMLBkmWCZ+4RPEp9dC
i9iKgfFUl00f91n5U9MGz+EjseJ0uwLfLR1sLCEKrVXGBt2OnZUFMC3rAkpSAinH
UZoANG5xDUx9ixrpzm82BFQ9kPXr9aWGgCG++WqZNkppMI9nNw5pKoxpCmOr1GAJ
NI80m4/XRqax/BfBPh4I5/qALA7G3lWEQbNYPBkzWdIHzKcCrOUAXwbKQ3WWmvjN
UqofTH3PSQC+11hpIBvuPU7BjFb5sN+/gpW6VDm9KdYt7L/7PMWar9M7yCuZe4y4
XBIULDpqWPH3BChCQYQzBoZrGOPnIi8m390JVCG/NKeQ+ZCDCC3IgKv7ZBo4aQ9Z
o2BwWSEOAu0xNkWON29GLfEZJvpBK6WRdVp3NUf9CEzCVDCoHGq1/0CsD0/Gl1bk
qD/gwFKchSZ43z5xRrajb3hITHOvE65s5j8UrYbv87qE3vE3sIKcQw7Qgk93zbsR
Li7r8UQF+VRCkUWRlSDGnU8LPMFgxzDoaY0EtnFzhd0IxG+DE6sOf+wNupeAjRuW
3fww5bUWycrpuAK3HfEdu1iVNnU+aU0EQHvMLK/gsgacnlzyag5EQCm3wWdwgP21
YJNdSYt3cUF3abqI9PbtiJlF9O57y3emeMZonkxIAfkPR8aT2Nv3dVvJpBNtaYkw
fIZRHlknj8oaOCBhCbIcLF3BvQO3vNwED7a7uMxaZ2hS+zY1tvkvXMF1+veGNd2C
JGi2Iip735WrB9UUhV7cnU5rRfHcYcJtiRtB6UTRPR/AI+UwA+k6Kqi+t0qwnz2+
VNhBsocLeUDBwZkHoWJjJjXGDWfZLwFIYpdRbuvWHbZOlqpYyaXFRLmWCIOWOCzw
N8WopWnmneDS+SfI+tOTwIHQjF59Ic1hhzmfZ/m+Iq0XLyTEITOHVn/7h0J/Z1ij
Xo2W0RBDoRbOEfgxYL/XpUf7hpmcK+W3Rn6W2EPpeaOX4QHOq/OdK3WSj8KL+BdD
Cd3/HU6MQe3Xk/XiX1g0o6Fj4b5wkCaKPdSLo2Rzud45dCpSWHfOMrVL3sup5z8Y
7KtxXfLHYkNuo34IhR0vKWs3TB+AQZ1arYP7cHFxCVgNmFfgliLdbYSZHvnAtEsx
8giDF2U7tr6hCsr3WT1XNZ+Rm2/hawvvZMcgRV11vNBMTGkCeNHNigOOh202QapR
6KCv1MgwTu83rJccjhoyoA1pmUr10MctmDXY6WBkkKp9BhJ1ztUF+rcRjC8CTZKQ
XAWix3kE49O83KD1qvRqegl3qyFgEmfTStXoYM//N9FbtnftleASl2ewELBKOPo8
Ivy8KPTNmG0iVYBOGfhkzTB/sC2RLi21x/2dhROujAQ+xGyYvxkM/BMKeACIwZ7J
s4HCNQj3TXSL9+TV4c6Ze5Qaj9nHXIhCT/aL8aFYIIGt3V7e5Wb/PsO55JRXbEOS
adMXkMW+cbbiuzJ4MTHOXjPrFK31wUgxVFYMDWdBqKqRbOImRKjLh65bsVm8sImt
jp5JKvfbB+VOAqqMKtQ8fFdKZtZyLt3aQvvAWR3gxdL72clexU4cNezDMOsNxAfg
+HAmhgCRFrrugGDLAXD9R6HdeVpq5sd8nFb/Pbe3QZoGbi+XnNqsykzHp7RQ75uy
0vBxfsuW+2dZeMteunEfEdmi1L7N9o6pQ8eq+l9RmLYcGJXEzeBbfVxHojxsXw8N
a2ouHdvwOFcG0wA7PfZvTsUvay2uFIBADzy0Neb4/dUyDYSPRIu33nMUdBuggEPG
OanuCmZtaJ/voWqh/bMwHomIwYvurg1UQsqmU0Kc+zXOSL8pC8ad6bCQILBDt39o
LfYQF3iqJ6rEqqfj8bvGthF+bjamshmWYbxMo/71rfg5VWuHmxRv8kC6ZHk6t36o
lwD2lzkDRcUlaZ6oFvoNssfQ4Ohu6Au/oCg6ur1elWZ8Kowy3JFqFJgSxSf/X9DB
29lKNNGSivAv2LTo/IZQDNTwXq8lu/zf0T4ZyuvoP4NrcGEFtYrY80GQpuVxiYub
8gEf0ov4qBEXkCbDGV8zrayq8L1AA8D3FFnpCQfkc3sVjxppw/vtVhZf8dSR0GXj
V6XXZaPURVNTXldA91xlVqxfCvhKc5UNBN6zPeIgvMA1PBG2KRQST4sH9EKkm2MZ
u/D34X+5RObbKylsHJ5JkT8TYAmuPGIJkC6l3o8FzKUqgcIEJJiprVTPV6cbW694
c1YDLWnV/G/X72Pv/F2Kc3N8GaF9CgXqO2ZDjY6MdQ/gfxIJnSEJWhQZcwy44AA7
k9rs0tvRlWq58XWG3aWLtPF2n+Z77Ovs1CYvli4LqurKFAkPnGkuGPw8ak8EKRdb
Ipl1AaPWnDokdRvGupNM7BqcbZivGXi0EfkYS5ZqeUoYD/lsGb8g0+giV38VGKC0
i/iJp/Yhy4UvOzPeL/Ymly4BEIba8GPKvep+4ppKLnBhIUZAOerGWiG+w5sZ5v/q
qMJD7/roFTPZx7BoHYNCe90WDqm+y1dgoGQIoso/BgiRcYzvV6KbOqWu/ztRPq+5
0JNzfN7dAZsk/Ca4meSuMpZvsUCM1nTQeT1bP62f1eDU4qyCh1xTXEpsJnqhXlhz
/N6b2Pmv9Vopi51UzN+Jm20b3SbFsNysVtmVpEpf/87CkbzQ7+ADe6/e8uEl+88R
no0pyDxGFWsGf1xHnap2SBqEBawrWZAdDufkbUerwHxOm8+ErQgwtRSOpoc1LDT5
flVyv3pUIBX2IrGyt48mqY+rrjOncnuTBt8r8vkwB76iTUlMS2XefGRnCTKfHTPs
n8i8ZaoTuKgfuZvzjLdofOGsqXGc018s52E6p/TvJD//qDTGyQmOMBSGB3Smg6jl
riMtdFDXFUsIEuEQVgup+zbHxsal6NVu2Tod3+1Wkf5TQ/gAH1y9L6EsnqfidB/O
EBSoLG5fR6F3m+gsy1wdIVWjepyOT352q7xyqTOehktIatDyXzbM6k/87JamLpzy
3yF9yuaJk4ow0r49A+OEVGzEmnyg1LCaSjbsqsbYk4jp3qInbHRgFYZ26r6PTJnl
tyISVwRA8QdATZnLWAKvoMtmK1P+oNW8tkZnjk3H0JR39b/cWi4r385wLsYzaZgt
odlytdud/oa5Ln0YTdqCgzKSd5dcAcX82yiJUdC+MRj+UW5vgnI9/cLtabp0lVvx
U0TWpi3llWZcUTtDozrRS4UH/5PKT80Ye5nY/G5C975QyHz692FlUnvE/0dm5V2s
nlNJ4cYpeXjDruMkPf3hOV019uJv6QHgShKHGV2aF/38Cu3txjEiPT5zbLJ3kko3
Rztv4g6YznwSyaxrsZOMp6Px1X1ZpVI/GXJcOHIwpxP86Deo2F6L4zc9NOG25Y7c
FbSxwTkiLtZ/Y1shmn3Wli2B3Q0mmsdS+okoR1KVLi5d9Gm/BsNehd2zdPQ60BAe
2D1D0Ah4V57Eyralbze3VNShp239KyuL/QBXgVp3v+COPl2j1FeKq2nd8nuQHabm
7nD7E/0duMCxO4CCMoEEM25V0DwnbbVQqA6RfVUoNLoxc4f2XGBsKYV0CwUrvNpU
LWHwQV3IWONygdX5xdAsVKYXldgpOHFCBx1/VH2YkUIK4fpF25NsLY4Bcy+F4exH
X/7nc3ABYpRH42ncj67LVb+859oHzsb19ywpQYxmMRBxeT801m0xo/z4xWf4h+S8
dNK8X9Az5QaIP+ona+2bnHqeuivW7a5285lNEvXWtNDc/d342rjmIGZiS7obwds+
p9/IgwdBgFf1siarg2pJ5aD90VmBeWUQUglTHW0U4JM61XbJLodw0c2GmszZzcsj
kqlrMot3OWMEciIBh3/+EBaxzSCAD5GdoDKTWzEQMmdThvR4SD1ZbX2bc73c3hGA
qFkJdfRo0dfLhYyYochsCC8FwbTDvbyjUR9SsHew3Sh22Ns5v6JZKT4TnPBLrZQm
mFU6ruQGF5CCM2sev1rwENqC0Yt6TerZnxU5bl9ZmR5bT5tVUNkX//vACfr+YATx
j9NRZKz59lPycEtYHF/5L97K2W0oINZOBcAw/6M2JHYeiyK6/Sbh+hXM9MPykein
l3jEXxaCTF+/8boXF1B8gKcTdn//Qd+sDkzU3JaZwSp7J7ep0LNz5TxrM9UaJrPh
juTOxFJCOBkodddUbvkI6r20y2XWMJNvPSVOZsOhwsXAFlekN/vsE6pvUeHp9tZk
8W19BSN8Dc4l6Uww2pVQBRID+IsHpv6Cxyuvld0Z4bSplh76GInUQcgihRQ3+0b2
VxraoYE+E/9OJtWGg4HCiVaqU3L1AgYg9GcVJh/4k+SgBoDIX0vmxdVK4WedHkTQ
Y2C5ixjpMAnkvpHeB44vnOAQfJY6cWXhxhQmelLYAAH+epIEjpI+l5eqwpsobwCU
SV6rp0Chkl0qpPawO6twep00Q8seFkm+fUIeesZLzLHB99e4Poe5E9gz7gKLt2jx
MISuaI+qnfZXTNcDk/Pjt/8KNKAyHegUFmXuVWRIp0t8ShKsDuRCrq9vucRD1vbT
NKFXcuyzmw5Oyh8bL6n1wpoKlghafjEmsj6Jg/51pk0MnADRTvLD0mpL04IEO5+r
Udcm2NrqSK18uuJt0ug1ZUb3jvqLfSfcTuS+8YfzpitqiqW3yM9Yh1fhdgbRAMmR
Z+OIJoqrPJ93zYtvvjeKl5cirNiIMshBjzc2+LbXdxFKQ1kddyLhioIGH5hR9xhW
i6fLZoKpKv2XSaKd0Bjd1BqoPQ+ewMFGLSC2wNBVA8RF7WtAnW6bM1wE0Hk57Ijr
q3GzCiJ/r5ovcvO5Qe7Rp4s31/1h1coe5sPNbhpStczJlgKSAEerc9hA8oCJG1wR
DxJuJdwwJOcFbILoQJRFOxpEHXFQiQSUG8nLnqJtL4IdS5pTdWV93CHI2TmeYsHy
anZASTxCfx2XhJT+6TgiORTR8Zf+9iISDCAzPqVXOsz8TsfPMAco+Pow9ltNeaaU
4/LYjFyZ4j3scxeh0AviCA9Fae/Tjli8JB2gOw5EpKBL55SDb0lvDD+fBKDtj2zQ
xBYNGQuPuV0yS7xdTu1d0b8yCjueSj6u1U7usFn+Xk4B55O5uwugXF1V6o9T4LA/
APITPheogIvkYnDXBmdIyrXKCyGBLfI/8spRHWch58em+4U4CyK7MXmLtzf9vYsk
sZCMH3MROBCotH4utONIKAiwU7VGb9SND/XQ+lkgEVR+/vF3ivHKg2YO2SlPEnoz
eObvBE7RqUwFeI1QeJqflN6HM0v0SF4BXUeE5qfgzn1iZzv205qc6ziBOEQik4FC
gnOhhW2SoFfG+HQo8PrKTTsaYKZ9GTdbPZGm34j33zRHjapa1uYVKw6QloJ94bwU
hcX+dRF6X82yC5r3QMOqhOfCCa6ftezR+tzouoJNWFPV+CtjYxWlDWeZmL1ktP+I
pAQv7y2sv2cAYWpWfJlqNRBrrOL9u5vk3F0uU5Zs9Xrxl6JFTl6nI0XqbQF3J81w
+Qh6sU6vTbq52v7SCtRBHQoyxFladYh/an1EcExqzz0NxOrfBRgI2RX+qUTwIQko
DRQvPQPg8CGZMA+Ch6K9oxq0VTSkYZPAzRgZGK6I8eOZr1/jaXZ4xoy2Y0ZX2CQn
f/AI3tJqyUNja1TNDxWVOlocb18GooSwq8pwFNZFPMU6qwX1oAVFpe51aZFvBeep
6TTlV1rASM8dfbXWfC49zocx3dtBlulDHiwzFnRvExNdz96uQfUCM5Ryrsbt56DT
EAmhUlin/VJV1PVvQT3DWzHjp/9A+y1PdmT28wuOtoUFNcP9Frvt48Ylga+bd32n
QMQwzJPkE2+KM38+T9x70MpYPlLyQ6VcG5bT0eVHQhbSCnKeTGTjRwrHLYFDJmhC
KKvGt5sofnJ4BRlsb17Pljl0Zgks8gTbXKB/Amt40F1Eb1xpbFr+NcMMVxyd51LI
EG/9mG2WfHL/sKPDLGDHuH8INeisvXctplemmNeG37T4jEGZlgmaSBHKzK/bPLbY
d2zCFr92n3DFlht4BWKeLvf2u7SYwLPEEBUJAj4XOhPy4BqUEW0Vb+yqh8VmzeN9
FXlgjh7fEDgxUwvjlgkLLlTqpuh+qAy0zjrOslEKcc0wrbnctwBuVaELunCnrX/v
NyqxRCbbZl+ab/TUj+KGg2vyX0Gg6ysT93LfvsRTgmkERMfPFSU/vEhavk0ELSmE
bo8PwEKSsOh0agN34LGVURNyKWpAEZ67uAqwP/uCdIfjPsZR2+CFDihtnwjD+hvJ
f0+0lHm6Er5VTgFUQfvREzs+Gmn5Zmxh2t7dvqTwiUR0suO56cjcTdgB6P6TRHr+
Qix9f69RVu4VKQ6jrX060VM9ErRAhrMg2lJ6REsfQ6yJDdlrGgcPCNSmS9/NwLaF
/5W20T9OoCnHA3y4EEZR/b7GPb3kqp1JzBfDE9s8a7eFZnOM15NypbjUZv7zNkTx
jei6dVLOkxu1mLdHHIx85hsCa7x+MaCYy8IevtpVltt10/hAuD+ZbHSA6J6p72VG
0Ott4+0HIdEAjEWMKf/45gnVMaRKM0YU5yy3JdQv6hmZ0a2BthteWnRBl8CZ9nHi
o6saI3O3mJafMPrsZ0QOzjt4JCqWOc2ILevEn+rch9brlAvDMOV5QIxxnBPVpjw4
vWn95DCRYwGC7VUYUd93gWswAZqjA3orvez6/KpS8u/Ois5PVu8oIceXWE1pGT6X
TB0N2HmTda/qmYUJ7qKaZ4YNS898O+s1Azv3bexSYFlIc3QPBEIpfzRgkhKOv+1f
QjqJjZLroudNYY9LX81b0ah4bqcnX3dDHtUAj9M8gVJNMZbX65g9JwiWs+/2+hNY
lqkviuVMKgI51xZeV+/bx6XC3KpRFQ3kwWPz2VwHzIp43QQG4L6j+UamLWaItRbM
DBrnqCWzB/Ao5GZn+QH4onvH42VQNIOCgAMY1Bi5xXtssvHALmJEDJWMKagksv6E
H5REN/X5DApsgj3+5OGIWBgb17wVDg3FCKyWaNKV/IT+KKgdJeCHvD1YURq6cAsU
1Rw79NbDm04f6otqhwPgFeN9qKBVxohcuA3bRB5Uybt6KBddzJxp8sQsPKho83Co
cUDrXuQr+iglnE/ea0Tp7Ljmgkg0fiMzZ0KFbV3SduAhbd5aPvCtXnc9+pDZgtYf
/HVFuhO4jVhH86Au2zl9obK4a3zkxmwrGL+uZ/KTPR/rc/8w6cOCEFlxveD7hUK8
3ij3eRwEWEZBMo7n9egREGZ2MS4+8+tj15vSqza0Rtg4IAc8TF7LsBb6Cofjo2in
gmXlkDlZ1C+vqF6e59O+YmbwkV8gezqbsA9BcQ8iwYuZNUsT509RvBXWk/wVDcmx
vx+3WrhL1WLXyWVdFo6ni/HxYgniYi6SymT0sYEAyToOd7CSvfFBvVzNtBupOSoa
1Y1cr6R1lBf3ZaO49u647sNhhakcoKOBP4DCeTkFL6ahB6TUd/20IgX5/0DYHt6l
iMqHPvA3Ueb4v0C5k7IJfE48KuRQEXhrvbergjo6pdB8+/KLeMeoRhfQ4pBIMK7i
n5K1X7rEdW1G0xC9RMBi0Y6CZsCwTkp5zEXGEQUuVUz6AEuoNTy6cxULn4ud27pP
gFEw6J8rfYbs+XyKaZB5gVJer8t96Um7V2lljILnYvgZBwsaj5DwugT8sqriISDw
VoX1FQuxuZ2IKGU5FB/0ombUNfLpqGgNfaUUwd5gBul5OmChTLCcHuJi760JfYov
myaQN4ztLGRyNrfXKT7gWW75mCZpuZf7+Rm8BI4lItWLwdvvd6m6m2kC4j1+TYpK
U2e1wyR+RBxkq31+hc1+PI++tP38TfAq9CXz4vi0XOzNmxY4JSqeO8DBzDL4ZoHl
caZM8fGtU6xHpjACGqTOVVHgzx38J2RVf2tWIxGEAV/r8hTDf0xA3d15elDun9qV
DONAYsUo6ivgyMmI4+aMrZxgPzB9oGZ8aILshfoSzqZKSLV9jmqjyOlqY6RdsIUY
YvNfeVZPtVD3sB0tQclRwL2d+slJbzkY5As174dQaBRLDhCMSw5IXOz8Iklho0Le
RGbgvAUdWSBZB2T+Ap4009Hi5h06ODA6fnm0EttTQAtWv9gWBDvNo/1ob5YYS2rY
KeHHZRa8B02wsgKdz/2zwO4POM8mTxIjClnq7MmBxtucXdR3dcqZ6YyjFJ5O7Azn
XvTcrf6u0dQay3aFd+dq58RJCaQQ/v3SvOYGB3WhB+K2yaESvr7ROo7iDNcFx+gz
eamew08j5hCVEerVHeYMicC6YCLWD4Qtby2zUnBb7J2LAQBV3BXQBvCJ/zvkCyW+
Lfu9ao31D4aHrN/wo3JA67B0cXR5sHDNt/kw89akXVg+NrDUz3gB019zoQgHlPq9
g7vezb2oDTtDgPGUXUIps+6Xqu7/nnv8N2wNp+Eweyp14HxoPP6VCDQrq3c0WKYw
Kf4ULMMu//Voaa+IjcYTXXLkQDa9pgFHhrdJKeZgWPYuXGP6AxhC9QeO41276Q3W
Hh/0/4AeCAnxQcnde24bqNjsjzrUyGwPUB66TXwhX97WkE23/Bkp8NXues82/6zh
Lt/zPgzwlXVKNlfKzcEv0c5wxi3htHPUQ5901fRDMckvcUD0FVlp+okoOvpJmxc6
y3n9IFauJtOkzRU+ssyWiCsZiwy4SxKQTc161kIuIeqzHGYcOwEYoWKn9IIf/m8k
ehtfR8Bv9ZmGRnDNx9AgwfQLIvi6nE/GCSOZJrscmTbKcKGxYsFlgOGU63wHqvZ/
K2/3nYjNJdcsvGJW3R0pa8ke9o44lOK3yZnwxWYhrynbc3Zez0YBYZWR0DaXRySL
Ywjm1atReJbdqZSDe+kiVfkaf5lJS5gaAWBQUsx5aTPsioUoFmt596oZlDxcCL/t
cz5NoqvIuScpaFClm8muUnBdNUfb4fsOAqIsdXim8nOOPljN0K2Uqb5U0rHCnv86
TlUDcHV694RqjNCxjmXfv8SfK2IxknSy8ZCEbdGPT2Uzu6dMO6guCiKJoGHZMsNF
CPXZ33R07NKPQghTQO1brrYgwfLoBsuL/1RBbJ8+pPVKezMw41Yf8BsT5fzVWwBX
n7UcjxJauNy2TMxhI5YDFk0+YZOZeucMweSlQ5HA7dH7wk+e2XStT7FoFWK+A6hO
wJnG5ZZuznrG+yVv+CaDma+4GdHwSE2D6v3cEiQREkX69DfhR0d3+fAKgjdVhz+0
CXiEq7lwoRDzzVwwU1gmTW/kUndKe6/nkgW9pu08PaFDBIjsx7VYRwqiMKcGK+mJ
WRYpSEPIQc1XyWRlzLthOq27mlR+6NJXVXcpqR/oJRQpWVXokqWB6XYHpG27Px7v
1+530bxRm+plktVn319WAKjUQYKFx8j1hwfBxytTdZqlp2A6s0ofMnKtIk8S5Mvw
ujjEW/Naql7K1/eIIsag5CSdKzO3Xce09Q8MFFe85JZQ4htDbxMJLFIQgDUGqc5H
yuN4isqm2l7U/pi4uRuCMCHKTAX1MuzD+C1dOkMWEoHMuc7KqGpFN4DrPO/C6Pd0
xp9FLZ+Qs6Izt7aCx03osb7vldMr/oN7NkG3E0UebYjbLavhn1FQkN5VB58ON109
VYZWFfoRvaVhhhRbBboSs0GfqbV1sXHleVnRPCC0KS5YxVsMfTRPDtBZLf3Ch5te
cK77lgtSX350tU8Pfe95y3DGB9w0AduWeB7UpP7D15DEF6Fx2Gf37TD4E9NbhSPn
g7KuGetKMNtA7G1qHoTRALD1jx29TlXZwx8CJvvjb+I4sZwrlwQCCtSUGfRK4Qis
6VEHFCYwiUISQyhAR0buux3MNP/oSFRrxoVe9x3/fQCzSGMBjOAsvy8mLfhhsDul
aE2JHbgJDxEy1dyN3adScMyhPHuvi+osepDEXB+hj3Tpdxw/Lj5VKnnTSvw+LYpp
4KdOTGFo9ZNgcN1eoi66sCmKjC9gCOouIAZxndQ+K/SbFwnFZj3C/tRg31EEvAH2
7Q1+xkwBCxzWcEuFmtvia1TvjP97g4PTSAqZIak8KW4E7l6V2FxHmnp1BjO8/pcN
8TprUhQx6ZRNctJhWbTzZqU+FSFewG+I17nCBKem5Z0XiSj2C1yjE+hiNoD1G36i
cyrFQbs2kVA5B8cB4PFSYVebz86otYcfG+o8k7zmHjABFYl3l/tDXBMbNuKRkqSF
fGSB77uDfQ7BNWMy0N299Xl/pN7WGhIcnOxly+R0FPTxGGfA8/YBkcd+G0BSPXUW
93GsQoWBokhefETqZcY7fc5MXD5cUX7djzW7DWoXCnvVwlvSLKWSvXAQV9cj9PvN
c/n5tnDsyJAOCCjQAosZTAEpJ8uM3M2xoUxLdKmmhrvl0oMlyWmoZ7scQFGfO8dg
2c0+e/C/4sXnaN/DAh3nj24L9nELfP/4pDObHWsXVIMn47Y/aOSGB6Je6YS0zj2S
Q2ELBfS2bBrSxIAx12dvqwi1CT9NJKUqYuP1Feqhi8ke4cgPuFPbgsIJAvO9gZPp
5j30uRwpafd3Saj/AJd8PyJrKXvn3zOl2Enx0oARKodUijnf9Xkywb3UEnaAN9Uh
lQEPyjScdCnPl7aT2kiesYauNYW8qGdyg/15yu3FF8uUjdD5yzKPP4Mc1HwQy47w
ei7WmbzWh0DbGytUcF6nRV5EItjB7pop9q5Xzt9CvpHeAfDh7oR+53C28YtfgAT9
6BvoohS0Amw9WUgt6eEmlkRioWLwfH1p3+SqAhFx5FgBVu94YnGkf6b6VUHDGxtD
6eQ3IHTM0y5oyRMoU04vFp1EvLtkgoyF6Snz+TPWQOd4G0xYzQPmLrXr2OUdgU8p
J2Cs8khCCWW9GCey7GKVxEyByIlvj+xavs4i/f4U11M8c8xW92QeHtQkX0zgdxZd
WiQtq/Kdb7gpajg4pMg+u1tqjUQAsjphtxwDvI+l7y25OoRgu7TT+XydRxqDS4g4
UZL3ORsdHaeASmJmrhppethv4CEj9oebjdQeGboZYZjhPI0R2pW0BItL0qLz4jas
1fwh80dRzpDjF2lrzGQiWbhXnVIjKwnmWGyiuiqo2wRkEgy2Lw1nZnS6XCxHnMnH
X+L8UefQTvZtk9VKsaH6hhFf2nBTzoGSNcoBx5dtP4O4rgLoA515C5c7joj2FV9K
ODp0AheSjQJRWs8mAeynzl3ssOdPgoypIX22e4dJO8dLXkk5YRn/wF2iKXwtofo/
Pc4WCbwGrZoYM5laq9Kl9ke5w+OIHTTvjAkjogb45RmBmfmrzpPyNQmv5mUbSbeH
w96cqE4ow3lhNBRd6RnbKyfSKU6OvuPlGcCmYhizttCHknd45K9huT076HiQZcQb
mddz651kqWMj8OWMncTHFmnBtV0I6lELwRomgtusk+i+ozTyCvN/tTP3/Q6b9cAf
TV/+8JqiIiCncFuNMsv1DRimP/TvkiknzGjliCEyYh7tvcG1KNiBXCyvVKjA65Lr
WJsGOY48f9Z+zS4mDmO2IVh1lXAawM6q9NjHi9VbYQHvwDm8miQOcifFkdFCL9Qw
SlcNOIzB6uTNF7YlOkUOB4vj33su83MBSCRCUgmg69gUERhA30ZlQpAh9yTi9InZ
De4S5bcZH0dUaMN4HDys30TWRd+BTTh4/qnpPSz8ulC+7PfnB3VoDCHzNp5kRelr
eQ3g7NoKWTLfbjiHnETq951T0R3P0AtMv0jhAHVpQ/WnCVD9sq6y1OiuhMWhviVD
QOaEmneNotwsjhhrI0K0RtpaPb318b4wsLhNYDnfsHHDrGrh3JjYe+k/ECHRweO5
/BDdljslTsklNhKTsvO7ZRqG6hSKW3ZixhuzoOzIrH720cRzdqVwNfEv/yihi7ZS
Z3PlAjSn2EETHknNcwjLGMxqY+b1ikRfarYbDzmK068k+PWUiFjPWf+AY18FWoqG
wSJgiseba8IEoArnDYDUEZ6i35RQzkgwT4oXlm+5hScCKke+c/8r+y0OKsp4b88F
FUf4Tph9xc+6/Vp6TZuO4/TOZPfw9zIXfj1J/1TsI60zEP6XnHp/1V5AzmYTLdir
JYDLB24+AkXbNqPenhMJQHRCWCiGWe7+KQ07jAneToiY0W9Rfy1m7SjH4pc2mvh4
hgkDYO4XgBGNuxJ6IbxBGgKNo79AuhPhTrfhDIk3aWl9SO04VoP3OLLRpr1/GyKd
9yuxT8SPofyzHLVdH91R7/v3WxbQOQ5anAmHPqtNLJaS537SJtUAKIO+k2bbQGd4
rn6ir62+dg6z+VWh4L7GjrvrUZ8ZjyRq0cjiff38nhvtNyZKQ5PlNPJAVZU3f7OC
/CrB/DCuRl7jU5qBiMJ2nn802KMUrTc4NScpTC/sviWspW5WseIGYl27BwXpfo0c
/xvoUUvRVatq8jD0wbvkLHQtj8AYG9+rPnElMD7+EwYSbzdZoMBs7JssDsighMrv
QX+2NdLEd/E3I0eJK8Z6vUdEzGD4P5wJZiPwuKkbnDwt0TmpmVR8aNn/BzycDoBB
UHpB3k91mBxGjGqmDprdAsXLbep4b/9Xua5DAQMXKQOEUTetJYMXBGPD0ff5fGcC
eDX3c8RWI79jIVmJ3Qk93L1PRkZbnS5DbM/sR41vptz03iAIWiEX8hw/1Cj1wCD7
S2Lwn5IujvdnalalJ11xoneBYxf4gixtLBLLbSvtEWAb+Q5HXGTxCif3MOKy4IsA
zzIH9EZmSenjM8+F8pPGrLjfXVPgaA1JpDuxQBgR8WUrYtGtqcNA8Tfcoia6lzYY
3fCvBKIY1yDXh/DcrA5/5zbrEYb90MDS/NofqnlqHCs+BetiR5s7Y0YbVRl7+zIT
fwunbLWw6AJv4gTh+g52KyfLAdePqgu3NZtScPkIzGPPfVzwXU6EJf/bdn1yVqVK
WYPnMANK9gdecifMEBCFMlYLp9iHanQoRkkbcgCqv+vxsqDurlpDs5sJrszC2RIE
T5EPpTUYG09upN5yWptAk+9lwao5MzSV3kQuqkHSWf6m0E07KJHgOWY5ZNjikOQz
9URxYDoGPWlhVh9TYMajKz88tF0wiEyOvPSAHOn8GOjy4LHfOQzaRhFvO/AfzD0T
hVifB5x5cilTNFvcD//CrfUnYs1Nqc0pzFQcb7YURQZ9fPSDTRRnHoPedptUi8qe
FkkADJ1vg3CfwUVF3UsU8ocYUw3H55GqQ43YafM4vPV8Wx+T+fEqwyRlBwKh9Dd4
qEv5HzUHdWCj+M140uWw52pTypeHQfHfpkB/d9agnerBoflhU4OVCX/LR5Wng4kd
vyb77J3xS4UJ5aDHA8No4sJihS5tTcm2oh0CPG9SSpHMwLs4t1ekUbKv6Rsg26Q0
nOp3iwc4eBrFFVdgWJgR0p0W1G+xbNwdZI8o6QRC3TStPX2HcKMXeEfMlG5l7Ly1
CZgKZQvGuuDOMYkA+yhvqAnBW/tAitftjHHmMWO3RMmSH0yvJZEBXEI+uIb6brvJ
iZBuJFWxp3a78KvcH+1wWDHkSc+FFiTUj7GUsiwvSznNqVAr8xpM5dWeLV5zcgYQ
qXBynjspLQ0ZPus8xzkOUQkVDGH1s77PRDoe6paNSEyozf71KN5v2DEDt5O/Rs6e
mOqj14UVFc/X24vEZM9IqGqzMa0f/Ci28A8Ch/ubdoknV63FHGxhvTdyjz7qXLgx
B3cIBo20OaDJ2EkQHbqWh8m8QJ6nkVEiv5MWi4YhNTzYDtnwNCgRWiU7PWFbeUgM
r9YVVtySmFTMtGIP/9fyRFIqWAt4HaQc4y5cF57T1uCnuf281kyjTk8GE8ixWzKJ
wKzMlD8EB1pe306mdAJ6+SBKMf/RoqSj9MCiqT2NXdSD4pewM+DbOIvkbvxfxSCD
O0a8IfGse8w8Otho6JijRjrIc5LoV5l/8Jd1L62r5abSIK14UmVoOaKSk6xov2N/
ps61j8gtzg2fkFqtoXAsLsERCB6XU3JMY2c1wULIzAGqwRYS0l6QxhCd1UA3Y0IA
btOaKZckz2h5qMxsaA3OSvhXwewkZ0JYKpfHF15fcPcFWcO2JA0dwYek2XmiQHtJ
Dd0VJSHN9tqHuHmVnXOji4NCOROqnqlKmFsRMjAPwFO8UmgOyGy1Os1Qsyv9gwN/
rme1f3gzFvAV/G/iFNR1bXn50ASfmouO8EaMj2862GPB6eRqZxr+Eo3oyeYZ0H5t
MtjDXfwLQHafQFySx8Msh/frm9/koybN6uzlv/bqzwO8ZDHdYai5W/Vs9DXkzjaI
l1ZtnEodXtSPscuAo0e7qck28hVdDIAyDtTJ9JZ1NVUmlsu0AN/snEDo177i1lG8
aaBJtaByK9f+UpOF3gJfMHxWmGIqIPVqpdmoRpxh/Jtpq7Jx6HkfNE41Ee81Yw6E
wYbgQH1njpTkxRa2fqeQZ77AJrcjRUjIGMO30QgsEwqbo4VKyG57NDinBsJ2d3ql
CPe4ZQqWDXyLmR4RiEM9b9vK5zZFIAtOAUv99SscT6DEXdcpM5voJhS2hY6Kc5Nu
cd677L7QVFicXUvNp5QAGlw2n0IuoJDgL505+x9f0FMkJfW1k7vMlwz8wWcPLjVZ
u42PqX2bYHlrsCbmN6G7BDU6vQVrOmlvBcxk09IJt0+gSKCE9Mjy93Gd6NyT+mVm
ZCyJWcgVNlC9hXCjxGNx6MKZYU5f3dGiH9naznACDCpdke8lr7smvjQbvbc5X0qo
VJU3cQm55U3JaOCqTazXwFquwG8pYsVnVQXDb6UaXhx2yR8u1tsi69hLr5K4jB6L
jaY2Do1lA//6Dis7kVwV7r2COdURla0bD+1cjx9rE7XmBfwqcG5wWzTDpG9QVZ03
MRZpZoZjyo/sVqRnTqhKUHchYLEbsmXCJWPvV89jQkENousOpwqOc3PHkqrRX1uW
4fVe4tEjn2ynPQx3VdML7xGXzsZgMCsizH2K8PrEZEp4HVQgVMfgUnOAs8AKI8/i
yZ+hGdx071zUl8J8jMZ7UIdGEk72ZD4L3e+ENyqGDUQO28HQ42KRzsEhYPt15wbD
wLdNuRvtd4FRZZCJKw129Nz5bm/CHMRMCIw1n9RhgFt+MbLlbsEsbwy/W5KweLeV
m/hstKVJ5C7tuNLJ+XhC6goPY7jaXSnqEvMN1UE5LEmzCgG9SoiL7njzJol4RNl9
863ckIEJqZ8Ziefaxw/3LryT2sUVn3aaMQqKZCzTmQgtfPbHXRQHYqdMTmLgb1sQ
h1orTaWTBSZBif3eo/cjIbEp/VduomAy5VnfLMXJNO/wIYPaI3O9/etln8+6x9Iz
6FeS7oLG0jpgbboVxB2i0WWmodb0qReWAsQpFdQkcC58DGdYw/kXkKHpOy+Po6tJ
093cFhfWCc33M6cn2vlX3sMt1LDxL7Ipt5W9Kjb4U1+quRFv9f7Y86SP4F/Swfom
rBAMiCnzpxicU6rAAjFocbS0WYIqhe95FfYIKbVjL5Y8MluDeL/4WYhp+lZGzKRY
FdE5G5zjYrG9ivztqPin9IEaoFWasBoC8ZuHqVxNvGOdfYBdhmK35zFcWpaV25Pd
2K+JwOnoQy0FWj8X9dIj06BstNVYOTI9W55dCXwEzlkjVA+5KBw4HFfxB87reKpv
/0bf2pLuarjYBrpMcArZfg6wf3vxzUsnaIkqCAlZqA1n/L+0enn9N9yvkuAQNtrD
c7fgXJZSCSrsHjAhBpOd2TrbwMobeaek0OCnWOmEwVuE0dRM1qQ+onUpUjbp2REh
SR613opLMr7nDGe+gSTK1goTKHHITfgsZ3RACYDfPhzcR/QPKL6CarO4HG2HLf+T
ZjPfUim+785wy2EdGMzXv3fCcLwS78t07hWREU5AhKC2hJzFqQbi2TS7+IHi6Hri
BdtmkCMJ+4ybIfBt22RHsA653I/f8atwUntZLOBfL9BPbxs9Y21l08rxdzEnQZ3d
fy/fHnBE+1+97fevrliYkzR50dSPULSHSWXb+UsX/9Jfsbo8BS+iSrodj6dtGYnn
ZZ4i4Gyoxuhb4f6lFID5k2pBj6gKNuD3OB+wmaSjAQer8JIHjj9rbQ+YY0U24keI
DkC6WsWBFB/7UaEAS1Zc+6nA2OwdVpZqdS0cHOCc2ipr4qUedqniYchvgckJTK7L
CEQDvRHX4o87pzSJaNJNrpVrxySYJSMqXhPiQuPZFEuqHxZG/NATZ713PHE7czUf
lGkTR/Sjze5lYORagNvX8VMgiNNqpMean3oRm8bK/hc0+T/rZMxP7b1Gb82+ddEq
AgUtkUaltlAOqiKTB3i2Iwcb615JL8HPDyrcxuVpQHcfF7cBgGqfhP+KCD1AnKgB
AOT1DX2SwkFMOUH9eRg3PIl95xMBFl43dLrwwu7RitO2MUJpDLt1PES9HJSIWUbE
2tn6s3U/Ge2L/b/1B/U/1VMn4ms9e4A7PmimlZEeZZWsWHovN8cWCJkUT1ArP7Io
CNr9hN0CzLDo5PqpldmzvB8J39g6ud1l6JWWdYXcFMK4EObheX3ygLzYVFzgId+a
e9whk0YQEKR3JQw6mkIvi/c/QOFOvgKTK1jRksn6IIYiS+fIMf+Sao7ClwmfE6vC
f5Elr+C+/gQOf6JeJ5o6CpIhT83X3IbCtppKN79s1HKNcQ57B1Uve0xqgSA+TaFl
Y31AhJBsDLLsfBwU3tGaRsO3QGNGjF/f+M2mLHG/xufqUOmkClOr/AFHGZ1k6vF0
qQ/3TLBC0feOauSpJlPkaBffLvkrUtpkCQFGpwAIkMqyw+55qQTBwiYYN9QKUA/A
SV3x71V1AUFiPZTFP0AaGo0LeP8kKVoJyNNspogT2bf4IZOXSwTlQuBTl1PwDDrt
wIgQyQRu3H0GzCCeaBaUVn7AKk54LmgaW+m3vmc34JeGzeAzB5SdGxb3FmhlVtl3
9DEfv7SJ8kIlKV+wlaAPeyrcLjsA0xd+xsQnIN3CgQ79pCc9bLzk9y42dC8vwMTn
8S0uUdon5AVMy0gq0zSD+5yfv64t2ZNO1nqP/BDy57MtUUKOXEX17LLQR+AIS2qW
Uho/N79npKLERmXPfmtANl6fk4K8RqJxyv+t5DDtDm3xYntu+IRfHcN3iVYEJMNa
gShKi9asrKHVzBdQeUo6xGXBV7pwlxAEMwolfdmQOrvOy8T0jdxJFnZBRsdtk9wt
UlepkZuJ/EoTT5/2MuO7Ou3jAwJV3aFxxDgAGzKnqeuX4afJRXQfRAQIRxDV4e1m
MQ64a+HdUrbwePU8pZQvCQ1d6pbMa+U6XJgBODmVaS6uAg/66TjfazjtzwSfVfM9
O9eOWQIbfKpW6ijx5CQvQfzsawEMaL+NTMTdOgummqcj+uOwoyEAlDbcFhO7HxAK
E5o6gfz2E9riKdBfMC/inQ4IVnBXQsor/EJR3UTuHzUKag1W5A6Yd81RNKru8VZ5
vot8gX0H3O0zPRY7/XS+W/uxUonPUEL8rPfdEolLKwsn1uUbOQEyU9SgcG0dYvgv
NXd7sSVRVp8QyRnkRgWsZ/qCMJNmofDanneZejN7gVFRk250zX+v19Z+xTjWXzcj
qXv8m/E5Fayta1cCyxATrThjhDurMUzMds4I/CaT6ts28uRcjiBevGzfSNHoxoj2
9Vp+GLHlo0SHOjR1+cZpgyTQVl9baei/MEhUZ/am5Tmnj/+mAf6y1NfQBOCMvYnD
TE/jWz0uZV6xpoLW4pvrmC/6RriqlMh7b2nRE4kgqMcngFONisrWTh2wcZQoA76n
cjF+mvRJ3KU0Ks+Nl+blrLKpessSGO24h5rhDNqAtGrZBjFS16viGIF2GJHmtuRk
WYA03KPDBtT867nr8OgIiBOtzlhMQWQjAbyiPdp62R5tUo7kKLJXyeV8QA23d4B2
2k7P9jmUzj9xxScVFRu11AXIFPum4abjUNhWpvtyEUWrOnK/6WvN5EmfwwLboi/Z
lnm5itU10m6AaZsZkZXtG/GroZF0wEROtD+zVYp6avUP+eJjtzakKIs1plshWOkB
2lEGzkdyiazCAVDa9uuolq+b6KSMRzuqMbiFM06stMNgUKWhLjP7OkbRazy8XgrP
PP+ptGBcSySXqM7pvr2GuqfLe/hDBU8xQ6umpTIrGsk0HtyFjRomZuiZNumroSr9
7NLC/O/7ULYgAOhFpi3TH8kEgieEgi/FvSFzBqpncHebqkRUIAUqTB4qjlyflp8V
w9hxzzN4RUQEe8E76+vE0vxNFvYG72xS3Ixr52vjZfbL+RdnXzPQ9Iz3yWdqNF9d
lf3G0NBMa+Gd9ilo3h+eNY/lnI6d7NGARWsQqtde4rYzckmjw5E7yl1zqAhC8eG6
IXM0Qv2QcyK9vDETe6b1yGoOMthawhkCUi9aZZhL74XaJer0RkUwKjJWNz2scPtv
Wy3YLH//vMDtqnWAVYCPCc/Vquvi8kq7By/u3YguMrI4y4oLZ2mw/tB/bBeI2qe/
TehUe57wZu2QiaPlFQWtFPq325MOd5tGn3Slf8c1XtDC78YhcE56HJCGTE9SnnJK
uOOy4Pmgdh+qzHDiHA5WXiq/sAk7R3VySxS2KyFSfpu4FubUdUbQETlfdFEpbT6O
L3bxzQr81CTc1Qo48opPXqAmAAhkbt1l25Y0EAaKi9Ix506S3UsWbBNHtRIR63L/
dYDDwNiKUZ6MmhgbcjmMiOXNB+iCqBqlb2wuirsOYTK70st/u/EurXxZWBDr441L
BxrnLLjnOaLbQknhBO0mCD0Y7AcATvl1RIhhylc+oQN6QMKYHrtuxPJc6diLMDFZ
+EB4eeFojpSlwL5+Dttf1H1HBaWkODqBrr45w52du4jKs2ydGKMGe4Nblgf8jnNt
U2jtPj/ugIA+WjFYay9q3kpqZD+FuL8ZQ1hNTgNnFzk9ukhrriVH40OXDhhZhyUR
yRcvWh4Kt7X4DyCXX5DsMrh00g537ITvA0Z7b/vMv7woLpLFsX+mFQPSCohCMFJB
fVMyG4kwZRd+ZXLTDFuWhXkGEzvpKec73qfDmZCHIyg4yrufE/uupOlrHRX6530V
pBYetvoMAFdrheTEZMK88cXbgdXWyzOd9lVEZKy2Of2q604DRqy3Ki3tIcMi+JQV
edESmId+hlQYkbgZ4zUZmMoJZYjEXcInIV93METVt1O+Jh3BeObUcz6I1BveYwpw
3SIoop6iGhNcbu8fTDZ5OyOXSfrWPUjPKFIZ0Shbnam++Rd1300cv3+aWMeAIpHZ
+SsxTYhYbBv/QTUTfk7sb8CaO9fMWF+ploAK+Misuw6+abqsW6r6AV7OBDNrvWjx
pNrJyBRAkwFV6W9594+9xvlqOQWkc6KFdiHBJ1kvMNXKGIMSTfSBs8xh1/zpZ1fJ
scwvb2nfTMxLwZCWbtZdkIJCpOOXVphSdRRNnEvylTuWy30x6YnDlUp78E6Qsqav
c4rmZ9XWNnscm/QiU/bC2/5lyozmao4tDWybYzKaVUrmLEt+KDT54XxNbJ+M1NE4
Ne/v5e2eksLtORIilUGUCWFqC86tab08hVnYkpp+EO+4Y4TSXg14EAiD8wiPcInr
+c/cZOQnMpjbIBZYY0aGkLAcH0IW4AFGOxH5mbJ/RRd3pOr8SLF3PcbLMUM4k0G8
YrnAfnlptRu8JqF5SJgbSnD6W9Fx70GCUnCzGoS/rzVHsZYTpdVe2YhdAJPUvrzL
D8ta50yMFtxppwIH64C9of6KDIW7qtHQPzBW+Ai5+kkXzDBxhRfksU1Ce1apYTAv
hTTBQK4joM/P/0qsDE1Iqy58EZMzy7UpLlepbzH3qNqs/NVyyVjHVqy+1p1cIMYN
klP7JU54Q/hXqs8H4XsMIHo/CZ3QGDZoL7bRTONR3dB0oRQASk1MNswvx3K1FHMH
CnO2As7G7wEM5WBtS9xN6EoESVSF4dkDkzlp88e7mkXYFLbz9raOZKQI4w1mzPMd
T3p/mUFweTrrL0LVgJAunMkIo4zrNC+C707xX4vUZK4ikXxbsSXMZMCPj20UQp/+
JJFqWr+MUyqAKLGH6nUlAb+mkKgNJ+zO7egRnz99a4mrLfrnMhWWlK5Lej21fjRu
zmDAfl2etIPdB9NEEHj007lG+jzfrlX6KuKY1dvCgsr7sFtLmTPnV22WqTA3GRDj
2ue5dlMStV8F92GojAr6YGync4klbbmX/XqmNCppulPcjSzwVXBxi9JpJ4NYnLE+
ZxaW7OudOl/LePJ7KYLksUibnvwGEOSAFfwiYQJT8QF5AsL3ySajVOeLHRRd96xO
dlaeeHaylNzWTkUXsLKjlkU8v8pWprWnfqO7yi4s6NBriYP0quEF+zHpDdsS2tQd
T7QHCTxN97BERgWg2+r5o5eAJOvZaiFmJ4BgoTnQ/oi7LkSL5kmNhEZSyWumnAS5
rbSvPvEVvgI2/6OkrWjH1jx+NwbGCPQJmaGEBsfMJ/3fPORiEVRHWvajgXdSQfa1
idHbxKzQDAc9SFJRkw38oh6x+UKR/zkdsJMePvLewC3iwgQHQWi3mpQkGsrW/2c0
LUW57Mnm+zugJRhSCti17g+yVXwbT/KSSmRQLTWUisHCDSvdkxJbFGsER7s4y3ib
8JtZvzw9aMM2yYAEk/8Tp2TKqDqrKj2DeNHyV3zS+X95hM8Gk0mLt5Dk0bC9pXm7
LBPQEWo1axJIiHlWIAcrOIuHzgX0UxUYkjICSm8fjet+Vl2H9Ec/QBp04XwQE3BT
qIDd7U1sOFxr172gRNeveHDFX1lwMSmmSaEHWjS2diapSfW6UolbT11DADWQ3zAZ
PlEt4epA5yXyr2S3Z+YXSDsng/WPAM7cjiaMi33nSZF+hk9dBQpRag90dta80756
R3L01zFBE/NyiSqgua3s0/Dsh/cFHm3R5JoLK28QUlAcLRra/lC2FZCSiXbY44d3
tu1LXWHuH/8jYPzW4aDs3vecOCxebCAYC6nrTArR+G7K6uXyP8Ec4I31nX5MiXo9
LK8Xp92zdekYJJM7JZgUuTu5p9LW/4vpB65aveVSrA3w72ZWHl/h2RpTQktLINvR
02obz8JFLLqDYzWF3GA1IQLleEqTn3CpQvNa1SIycrCgb/2Xz1rHLEIFs0cyESo4
zUcSfWfygsTY8rzI+XPRViJq4C4Mjaz/Gb1HE0L3SoarnAoBO6JcE0Vmi2QtW8Xi
eV0EI+W7/nVdNJLu73QBD8Rhf4gOYPjFE8P6sZ2onLDOKAZJ1mS7vp6GoBkuGpjy
HLpilLOWwM6SXHSZvQkJf4WEX4Uk84tk3/V9pMxtc8sGxnhihGsHtTys7z9o10sD
LSRKHAYEgzrcPMEHl2R7LVeKLhNidKHXw6YdnznROrovX+IPaaRulhSmiELRFubY
08Cd+vZc2i32NT+pd5m/R0eKn9YQWzE41GGaYZm38O1jPi+A49HGnvu5PWU9F/Dr
dlzgJ8y6D1r+QgtwRq3C1XI6kxJxKfxZn7I5Kcra/CNsxNFuxas8971svkIpkjBP
TF2x7xuvtnp9kcP0IdeDdSQ40etkPam0lQAgkh3eez+pX2fj0Lhin5dn6eOqwHe6
aJMwuIsF1bBjAeb56Yo1Q5HHFTkmc45fc9upNQ169rZSZfsBXk2FzZxU9HvhaOZ4
+vq7ELhFs1L3Yay2uoyHeqB/Z3BG4u68x2UExYl4J5y+b6+2lCBC1bCHxQ3cIFqJ
2IzPtyCFpKtrJipxKzrzJDPnsnUrTbP2n7iM9eNpg8FgjU22+t5svxYlWbG9JXIm
6uBh0E6gN1B8G4LQ9o4WZdRN1h7vCgfsGF+Jh1A8deHIQyXj4y/4clf5VXQqLpn3
2ghaGUGTCXNttEO4ffJHJopivFIzLXpBcCAYgwhEYaQH0cxNA4r35H93JhtxdCe6
GaC9sie51fZzznynFN10esXKNacfh/WS0PaTmLcY9fkyD9WYAO054ovkXEJUu8QQ
gZhNeBLVMPb+AC+3WeJ4oyABNTQtZ043PK6WDfw0tUSP78N0pkNz5lyu9skUbM4c
hxYNZqLSGJwcOzFbN64Fstv6Jqc4+cX/YJJJBEnuXt/4ktyMQvH4UEwf6FH2wNRz
G6At0V74Y9lvZtq/QVLmMljifj6Bc3WLTXf1lycP3sRxEly8D9/OH74giVxtGVEJ
XVAMbuLgORS7saddKtBetAgfiB9kxByvkbTch40LejgrLtr8M5aGcnpbpVo+YoE2
jfG2PLjfkJJDrBdKIRbEQ4uqPkxhRzf7ob+41FP16JxWXAA21Vzp2BTl45LbspdN
LwjuzArL2gODSY3J2VtnRHQXD4mVJANsJNaGb/9szmpPnZJd0Eh1w1HK28d2cABK
+veh70A9Y0oV/5HdCsKn8IXYmufy1GFJuvc0Z8gHI2psHufE3oNjG4WjWAr956KS
cO2w4KwOd950iU1PmeMBOUrSTKE4SKD7KMbl7XInx1imULWas5Al9/SqlXkrRKf9
hOb8o/OA4pQOEMA6iIj9kpCMhNlWoA0lQWQJ76M9kvJCjJ6P96oQklSzFuQGIsej
mdVSLXRJEdTKI7xIbZldxcuPv+bKz7/HmliJ2+nBpOHGIGLrkyWXmL5kBDnO0pe9
UGep2k93WRA6Xv4MKFXXOMUjuGBg4tT8f8PjfLDydSNfZfNeXKg36jLwRTn3CBTq
zx22xdCjVX1UUAOZ9Bu272RQ9bQYltMWuM+Zivdp3TZQD+NIPThSEXyQAEfhYavp
Z3WGrFyCPLJG+TY2W3U9M8GC2dJAGRzcbQVsHk7pTstv1JpPiuVHI8p+WrumCt1h
FX3xJLeeKSBicZnS3ApcIPa/Ir/MdWBzWxHV+/9claW3/aDVKQnYTCxcCCL5AYn5
MQ74xP3TGw5Ow8lJIYTSPSHJkPsUpS6UYZaIdUJ6t+6P4ZJeTBRd1Z2OxmbxISw8
3g+BW6JcERoAAhsuB6UhKRAgE+2IFbQnCZcZf/l82tAiuEl6V/eXDdrqIZ1gc4ao
wF+bbfOMn1xb4AVLilgQxehmd6/pAVx3c0PFU4ugKKUvz51nGL7CHDOevt+aIF/P
B4t2PcTRu36l434nb2aSLbfHfcstrqhFws8+gURpl+yn3ryZrszsVJWiS/NaTjfA
+wKj8nY0fA/4tvJznsMaVcK1l/vy8clnvd1PWJOJEgCLLu5FJKwVRT4oJE2c8PNF
3UnDBCGvHYtFs+S8ujn4B4kUk6GZoqJCou68yImrqAx5w73vBRBsstOgNDguk7gv
DMhote8JYcAixdk2lwOIP6UvTI5X4J8o/qG1BuXkH0QBaa/jubN8WRWlxdkvphqA
/MiXqvSHBHRuzl0iEuLSGHGUf8WvRBT9I09bPMqmloNvjVnLo+KLuuoceN0+7vVF
f0wGfjfMQy4U61SaIBCsLCd1KQDsEKy+eAge8amF45apsKEjwAsAq/4oWoYQVrRn
mlNDAH1vIhiiNK5XfTUmpx+NsFvLQXnKQiDgFKNnnj4c7VXPjJFO80IW2cwJ/sYD
QXROJ7wgVNH4oqQ3SvJUAWm35Y/EN8mYaSklPJSeWbaEA2h7qW1JUpGGv3XqVuE9
eBBujC8zT0brDM0aQ+XW0RDuaS8QjqAUWM3uPucSJptfd+iKGZjQ9BTl6a9Y+S3l
u75WJIwcN5zl132pD+KeX5xe4lJhPufFhByDktqndvzzlRtg5+kKi7b6SEsfGRR5
u6DHZN1NgNt6TALxgFc8ZVPSasspiKqfWFjnkHTTmTI7Ch39elGCXZDmbkB4qWzX
+d8R+jUQfEcPgYz4OB/XsZSX3kreRk0TxSOl9gqw3nKfDtaZdnKKpAgQIeOouYzC
q+7gwpypomfreuKnxHIV1n4mAJUsKHIZjoJRLd3sezfzGML/KVavciDxDpR58f8G
B7SmRbBD+fYrxFE79FeP17bCW8gsu8smNK4gploN0HqLia1irddkHhCXu9wdgV8L
aHkGlF32GSiigCvIYW6X+J62Mv0J3mK4dr2j22VenazRfRBSCuJUUK2tXIpzQhW0
Od3H3xWkFUc/OM8cLXGm3JfHJoBkjiz1ayBsMgegDDGMh/FFpYc9tsEDWZIewzex
V2reBFWSxspwBHxppbB/8q5xLdgRKXHuSdhBQZt1Cu4hsdmupF70YdRjyFH5Uy4r
smiI4Fnd7sW8M0caKpnpT5J9ygP+hTFKPYD38rm6nj0hsxtdqu89wom2PtZ1S3o8
MO7DaH8G+06145iWsmxfWcibCEMgNTKvyIQ3VMC0/9/EpTMsVkBJwp+8Ovtf5QNy
OgN9iGn02Jqr8Ish7KHTLAZNc7i9wmNUuAjdYt8KaVlAw25RsOcbqT++I4z4h/Us
iMNcmt4aDwxWQgKbZQvMGQuMatft8h/EX8vxHAjCFiksj6hugHpnmYMGKQp8UCc2
hQKA4nwh1dqcdVNF0R+Qu8tsQaYq2LEIU10a/hAW9wIueuCZdXUcdhdKYMIFkw7N
yWoMGyAAiPSzVdcQmziufBlanmK1KqS7Wyf6hgFdRA5vJ+gY2jfuq4/8wcrqtgsa
rIMDcdZRbdYC1vxt88/3uCrTrt+NOHuVcyjLNfzIJuULMBPoxGVdP2w8diuyTX3k
qgWdSIjQEHBCzG95CwgG9yRmOVyaXZEAJKIQDWeiHSpwAkLWsaQpjaxGvpXfgdS4
+HnozQ3DlPFbSCJYEYq9GLmS04dn5L1BZGGXCOn6E+NlMajTdvtYlz3BRtuH4YWG
MNRJWyXHGq7P71njNa3Gmmzn/kOCYjo8Ia2T0qCdxhnIy6B4oazAgzd72JcQcUR3
lFR3UUwhdASK7MiOoZf0kyLOWPZfjUtYPC3rShzySNMMGgWA0EeNF5YlTMwzoMn/
PXp3WK+kRgCO3BH/8FeFqJSxBvu/DLTxJvjLUuAiD9jFEXwr2zY5Twpgtc8bEzeF
XTYm6k6+qHCNW3k3XWunHEDWGgs/phCiZuJlgRt6rKUlXpDLeUygtR7IOO1uYdKn
yYl7mqQfQz9p3fOvzlKrNRtwcgtajiQRieg3OCTghyTxEg2lhIsPnRitcuYe4ZzW
QwMAxAIcutofwWbucvl02hNpq4YJptu10l38W2/KkNgjVVAJCHZmY63NTQaiBnzk
H30DEvGUhNwmnbdN31R1v1BYvnuZompryLxp9MT7sEW72NbgSPO3J2IXZ+QLzqwP
55mmw7mUGQSMhc2Wc/Er6LM4fYHLjvW3FygIijEK3WObpTekb1tU9XPJph/qcL06
acZmkba+54uqOEXLMFItIbsdKszOVpZLJVZ1Si5r9O70DFtkb8w5NYoeI7nj9VHN
YMW0aB8wekSnK7rvKD0IOA6mvQaIKZyNWOYVZt4GI63aZiLgy4ZM/1HSeGLWuBcs
GkrPrTattxriaspZH/r1IyO+jx1x3kShaQxH7bTCv/iVstIF4VDrcS2ithFwGolw
O+VWBDHR36YjA35Bg1ZrU/W+kt1PjQd52AQ/Ngk52fYohEjuFsagrdtvP7a6pR6a
cObrRZL26lnkPBuEx7sYu6B63DIMmIpjn0MLXWbSyelzXA5GbotoSLvy84baLAHP
+taT6RTx+evUQBPNK7X+T1PKdTo95QbkQauuLd6V9hT7AIZoTTBaOw4Timp2+D0Z
Y04UpWpuaf0xreLBh1A6O5bqgrVeK7+Z1iIaFUFjJ/iT1DJXuLxzraa5K5p4EzsU
SNCYRlMYGAj15hJx2jenJXODtOTcFRB4UAN0p4l2njymq8Y3rkeWFZAENXA7jvs3
DTh4mQQk1HZC0f4oH3zVhOGCLecZffisg/SaRngKxhrBJCPJD9yN1rHnXup2SA7l
TGxa/8Zd//MfLuqPsXohylURoAJdv4tKsZu2+llPPzCCmySyasrFuRyK88wokOhB
liCXl87nvGpa5zK4slkbH8TJiPFVzmYHq+OHPZDE20P6pwkV7H6eUZAlEgJU3gWW
5Kz4vkQpWWPepGbbCzwfoC7DFbnfYKrcPGJ9Bf4TEqlmP9IIledYgfR2om9vXB1n
snzI+P697IAqjF0Z4seVEjm/cENTYNBPZGvqBDCUu3SskBIVaWfm2E4Lmjt5qGFO
7YmTdIxIXQA/frqLUXbCa2dsuB+0kkrqeTYGmR+LiUKLD8X7PRZN5KYasCiF5Nc4
JCLhydkLel5VU6Il5LYbEkCPLAAcOo5lpfESZaaIVXLhU8QNMhcKNOGQhQJ4c8RC
I52BmoY7s8q8A/ZA/a+LwyYd3qGFLqwpdW3qJWzuf8X4iJUjemC+P1Xd585oWPCq
o1YwSORqQiQPCh2zoTwo1JvAFwH7hR35sm6j/K7oQspnlUpu62hExwjktoA4DaPK
Zbvt/2+6cpsrGNZ/dQVKm5HnS95/c8PC3AWz5bneJaSkSk735uwVp6IGYVwgi+6V
n+mz67ruUfI5/mInBiJU4C6+eqBXuhFNz92G910i+OPZqHBHHq183l2nzWnpDrYu
0qCwo8ZaBM3daN0XBuZgGN/AnKl1tSOlriguvFilvPg+jf+tdCTXh14OyFxnCSp1
3S1lDz5stq1dvekM6IOM4oxkSmIeuC4EJ6jbFEY8d9N/bNEYDG7nDyM0ZZ3Qbh4c
xmLRwKD9LkW3NlaIkN5kwAadqejv6A/60FeUYAbHOBgIFd7f6DSKZ/e9BaSVGr3T
I001X4QJ1RQJ29paN3/RScgowo6au2UmffQ5LTC875fatcCJkzcCUYA9W1us3Fg/
BTdL+eyk4xMFv9cvYdKf/kWRlkuVT3z/pbAagfSlllFVu+eXr6Yg7MACEgjaXvPm
RG1Nfp4H2GFPu0FU04TvXycW4Ls2VJetE4fZ3CJZED3hQLJe/L/74E5P7foat+kc
Rme7acpn8KfhvJrF4ZgI3txTY+fe160/g6lo6AoUKohC6kqisi4etazp3Emebc8n
zEuMK9JUEjdN7lq1WMBqQZZ8TFB439ZAbpgfQJeoS0lElR91kkjgHB33MJqLI7fq
Cmnp0yTwXVOjo62Vzxlay425iTsGxLYDwAHBNRwBIzC/MKMbqnl71eo8Sj6wZS5G
FXu36UyDPgmGfT0ccSI67MnIKM0CVi2fMmRYSLypZUtavjJ1213NI3SgjYllu5JF
rqScS401YZwFoef8A54wGzNyXQvvxFP8vkIN6X7Y/Lw9RF8Z1EanJi555V3CU00q
kRgbHmF4AfVV7lyYb/A/WNGHWi2N/NXAkWXrW7rA1kDv2SrV+WvpxSGq/WUN9+m7
ilw2E5/56JtjzxU7n6BEETfiQbqKony5f5TjfDLKcv3qbqTBu5cmFEhIYyGqF2C/
ZGGgSXZdTyFdvEibRu26Wkt1dVf33nYBFH073+Wo9aep4Vk3CBauTblLylN+Tiih
6IlIuBuvyi5z7nVFNB1le+ioLF3VkgLPTlOKSBHFfU0P+k3PFjXjDUpL6dR7oYCp
8QmdcbnrCcGbXrO9KntJG+PAt80jG0kv4YwyJm+ly5Dbr5Ju8KCOuuS/lOybdqZr
PA3AV6a53be0scrTW49Kbpy5kjz6cfEsbgGE1NuiQXIHyh5nV74bQqjZXgSFES/n
2TPzc847hNe558m22TIpv7q3dhEUz66A71EXZ7W6csRFEYQp1bHPMDasUAQcCghI
Ct15/0VhMtqBhe7quFKgjEXNvQLz1JCFu82SX9q46a+XGAocVwPn5HkL++bNJ027
390AxXJY1k5tTk1fvYNwK/0OXCC2y6EKEcB+OrQW/h5fMFnyTWltNzKsWdpbcpKl
QBBJJFdopJNW+d4p8lRXAml9HhwxAiKHRxukG/dn7SVjrATeqkBvnTzPrZfJcAGE
N4V6nQLz7eP0F/015EoH5LMaKz+Cb6kT97gG6akaaexkL6ABpDGHGP2IDET1dBUq
iUJxWooS/tIINud5Ramahk55cJi7gMi3b2I1YjSldRfTswydMItePjvCFq61UiDf
1mixN3s9EpI5Mm7qQEk/n317lGFdp8igYPVzG2LxzQT9YETzWmjYs5nC4a5Sw3Nc
+CkbooHiaSAn2JUq1DIsvJokWgtvaZ/TwiAxoEIFQn8K/EFt32R2p8UATJ0ja0Gz
C+JJonNWLJ6l1MWiogGsOFY8FFoDTp2w+2PuJibOfNe+cK+RhuMPo0O60/0sPMfk
WMCu7MSjzYge7fviEO3MHCkRkYUdDtaqpnnEEQDZiJFVl05rDW6L5ARE3zkHFltc
ex0W9sdy/q9tudX0vBDSB1I6piKEUzLkz5xdiMHpJDHXScor4RVOJYic2LvnPX6Q
bZrP3Iq91ju7zUBosZRdn+M1i6Xs9DTjgA98pqemVgm85uxejkTuL0SD7cZWU6Gc
aIS/UL+JUBqpwCkpAqU01oZRAgw/81+aXP+NmWGv5YTqBuP9ZIWlNH69l1OnDUPz
xXBwajaFOPMxRVMjRIT1KP4eUNFWlqfajINOzIAABJtXib6uQUeRaeVUGRRayU2K
jZsMGo5CLzXfe3OVSWElY8IVGgWLVsyQbfDbtEZPfMKog3sjgzGloG1vZLNdpwKL
QhVTEwEy9hJ3Hn2aulwqrnbiprhEiqh5W9D2JcU8yXWt1Syu1aonhOAp05O0u6CX
`protect END_PROTECTED
