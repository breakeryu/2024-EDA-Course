`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HktzYUQuoxUiGLvXI5cVR0hFvgzbr4uuJWY9Pov0mv2LbFxspvbMbGnRg5bYvdba
NStF4RjXTKbT6hO/uI0o+/ImBUx9/BTPMdwhpHW8nwUpdAZR3Dt3KR8BQQXbDgpz
0iERLS6L880jyoB/abRUos6XlKmb7xBMebNrKCrUI2buatXI3Mz/f+Ep+h+tVyvi
+T6k+iregUTP/LdRRJe7lPAWSDDFAe+9C+Be38aWxAJceTpWyYGCtl3NyOJJdhv6
I8eqIfde0nZJ5p7CpJipZiB3LxN5vvI5XtuE3Ad8SUC+9hCtRGCYQncz9NKPkmc5
PeUvQChBI+CH5ZbTdE5fvuwAdGu544GY3DNGZrIrZ4De/65IZZH1m4blTbsuxOY4
4Om+M3Vb+vX0UtSQAxFhgq/oAQrTJdLLNsA9LB7pZ8cF7NL+AuLhOk9R6CpmQsf3
W8TiNpg8KVvx5U3UP/81ua+3o0zH6wMkJAJcje5aww2cfcAyuib567Nsp/Qsv+Zc
F68MMlgQRDPJWMc5Dq1lUpS+f1MjssXR9OzxsDRip78D4OT5gyF+rfTsXcE38skJ
lkYdYynLqbh0tktjxUlx3EKRX5D97MpGi2JBIDZbsHyateBnFFhE/J7r84DArHWs
r9qVghtEmg+qPhfopNwrz1FXwn2AxmsVuzDoe5V3sUbyUvsCrkDJOzrshviRKKuc
WP7+ZMQdC6BjZi9iYpPS3iQItcrfDHj5acQBX0CAXuHxjmpjHQPgcWNElhYBTa1H
6JKHM1jjJESREvLSsVaOHjbDuKSNAUb5jMBUJS5A2bTB2sQ0ivfr1l8j4gvdpst5
GXkn9UjK8MMC+iRHZgtRW9zPV8bIYdPseXgzJ64mQH2IXOipmdTUCdj7HF2s2eV7
SyfnmWGs4c/0RTAzP7pOM4PlOccN93FCE4SR4Geho+Zas+ktB4RitmimqNMTAb0N
qDAgwk6EL2RzJDZMtS3iCE7eoJ4Xdw03bORiZiGTTUVXrmdANCdEcoE8K94HoU5o
k7PTAHT160XONV5okuHmLzE/nbQdXPYRumrcfb4y2S+2GPDWjafOqn5h0Ixjum9d
/66Ku7u+LhUbdP7/UJHJ/PtMXVe2PZFBlnUc9y3scIc+RYaOis6U5HVm8w984r9b
5k5iZpGRMvIIcjxmj1nyHmlPYm5v51w9TIc0FtfVy7giOfJUmI19D2eXR+47yXTe
+TZfOd4il8Fm+FA3vZE1AeDpAKnagicX8a98J8nWmLf4J+N2+tVRmrjlOWRQcthW
o/UyjeijC7OzNG7PWB390MeEjYrA4iDRFynPEU6kSUm/dFhwCTnmssdyD9DXrcvZ
NU02CGr5msmmVPBQSW5e3RT8P1vGR6BVhxaxnp0efxeXMyJ+WcjUohEYxA24/JhJ
47mky4fTarhiswslsolQFChQZkPR3db616XUo+3bI8sLW741nhwkf/JGxaXcHog0
yU2Xs5aSNduuutUsiiwXDbndwpGkUzAO+TVvPxxtF9O8cDyUYPjXK77xLHygKNyC
yzjDwMgpo1gAcn5uMC6d1VT5et256h9udEe38TSJBF/fsy92nC/ngDB/gUTaNYVV
2iWTJtFEiA0hDlrLr8x4Bs/IqLW0GROmQEauNhyR+J4V8RERvF9Wile1EKP7ys81
QSpZVf6Uk2tkMyYyIoj+cAbpVR2VSBHNYHBEiR9hyetHOzl05nMp8ZgSHBH8eLvl
wuZXWyYrAoDd6Edx3AvJ/xTTFZOerJD+Nuq+6jwx2fLxSjfRSLmEBnB2S6iCfX+3
gtaHZEB7LQd/SUQ62g3z9B1hsbJRDGW5nRc9BLhT6SgaZUVH/o4KzI+8tkUt2p3r
EL/hEFde0UezjDhPXuJXURMrbiGzly/IdzTj843G4nIqyU0iO9ssYvcehvWGCP0L
8ViVhRChG/tOIfByG0LY7xbiatMO8u070975X7Pm6YHtl85p8n9QjfXPnEsRPTQ7
bW48DkiBNbC2OBlSFbWYElb5o8ubZVip0/t8o+6VyYCCa0xuvofPRK5TUY4ToldK
YVqvgfkCtoWctfr541Fv71auZobNeAa3k4iZ0qp/dAZQg04UrtAvua+k+xH7MlpN
Y7Wu4ck/If6JZOL8W7f6dwFyipj/RniOJ72ph2EhrLG9DmO3Mi4p5T5WBLiYp9pB
PKNVen/JJaAsyhDc+feGzIj1he0J9AC04Ke6oqHTnCmiaYOGK9baU1PLOYyHdVMy
jPHCEYF0UoojYGZEw5xeHzsJOoh8Qosbi97PkQSYbGdESRvSRLQ7dVGv0773OWiW
Nfc+kjludMqiNfbxwoGjfohufDKZ4HUI9dEsMHkWTaTQUnZzwYkdl0XQfkVReBds
R9d3V4KNHw9SBXsyFeb/KxkpgjZ1a6iT+pinvlc+0carnIIARRPcABkHv6de+lm3
Az/1QklXf2YiR58Bqk33jnTRWArpfff9h+sLck/ZuKyGj3B4RIUWPCOWfZ5kKRTl
aye8ntm6mtpweobGkVaS9/7orqfR+u0dfoTsQ874Eb/r9t9XKiCp3Gyl7zags3g9
7qVndOLxOYQn4DDXmt82mVlaK95k/SwkYKERUoH1l0yL34KAc1x4T8wJCHrX+7jV
/9fPcMo1/jht3zs9TkPNa9QlsNP9SIqvMCHbV1UAHnqF3mO5flMf0idxq636/b0L
ULD/wyDFQqE88jB8rpHXWrfJE5nhg6h6oH3RadF9S+kSmIwa5nw46t2jyxnPNdI9
liTT+FSvl5ls8qTOGOfU91PC5ppGLYns3Vk1tZ3ZywqrJafxUn7wGzKmHLg6Y0Go
jOBbByaoF662esoGOIAmTMQvH+J+hf9q8wQw5CMtLYEHvw+joTdbwVRZmEX6w1Md
4q7/AtDCUN9XgrXBWz9xEMJ+TAVBqGxlBMRue0R86Q14gjwjcFqvdMhOYpdJ8eqT
yYXbWmnJqg6aDJHeldUrsXJVchL8l5g54VzQSM7aqFSW6wrNpvUZAMGik7F/DY39
RVYgaEtKlk3YKEPU5sdKulr1uklvmem3ZDAAig0RYF0JYcfwrcVMyKYMj6VMEgVP
U1JqCs8KN1Upz9vloSttDmTlgqbDu9fkAZgXXTJPW4KT0XZ0FWvzmvNuAfRvCt7I
2S5l3ZC00lOebXsVjTzQuhMPvDns+r7WdrrP96sivyBbL7FyQBIrAryR30uHOLPd
E793MtqXgfyOq1RWwlFlWBJQC0r/93yno09FBPpTK0iN6TB2xM9IE1TSSbs5BsEx
81eT9jpZvxDV8C/0hU/QWjq8qFusiq2s/ooACpUv3qKoVpxizy/Zip3AvkHxq74b
RmpcNX5jc97G3O8sJtjPjTNEtc98O7b9SwxSX1ICHq5fJ9NJ7UvhabEBkUnM2qXM
hg0zSBZsjJP8mbt4E4wtd4x4Rlihmlj/VI3xFua9PgpY5K4nb0CpON48uTZGXKfM
DmWIVmaxU7FSpkXQxT3EWhM1UYLcK8yitgUltv4YSB5qxdvjhdZcDFTCEe542zGx
qskjjkcfjgK4Alf2yZ974pXH2ITp2lpt4EivemTy4VcfRPfSa+ww5THWBDaPk508
HS4cOKcVXgfoPI1BsqELpZgGknJbsuH85M+70Rxz/1/yjtONEB/+t4WIyq2yko31
+9JNvA0/jOSe8DAFXtOeZvST6ybBM7jLjoyJJ3aAgFCNSDEBADcd0yqAlenEtWBD
8TNjXErnB+neyLWzHPC5MQch1BISYof0EYGpHNy6aQKpLkxRyrUXlK9//OJIrlqb
G19GkDJdfNpVm5itDNbVBRbZANHjacYrj2MHzUX6fD0Sdd7t9h8pEd0SmDOVNRoI
Qs2smAuHxDfNoSsLmksVN8RUoQ9/YEeTcj5ugCffg3gChxJL3D5kKx/587B8i+/0
I1avOOuTJpLugGdEPbj/j9W/tIAcaBkHbm2p6d4O8EaO59AoJmzrQkJhdKT3znpz
vjx2vp/ffJsSXn/pImA7u04Dt+UhomUY2KKmZJrL/BS/wdLDswNC9atm9JKkvH83
PEZKZw42FQDChnyMQIVXf1U+CWJzcMEJBiRQr/gGmS+pWqxdo0/7vim22Lx49i+c
xco0NytoOBNCs1zXTlGKovO+A2aEx8XY38iwn4rqeYgNX0gTm+vORuv1mPO0S1fA
lRHSf+5XNV0DZyjR5kHVKStQTolK402GGandounEBMWQPgqiKmQhgpJyYqaQXE6+
/8lrYLZbEIWdNVNp23RFf3U+4DX2ZWU2D9p/pRVt6+fXwJhORZ5DEN388PwPmJVE
sIUm6nDqEt95k+8Yfy/MLlZg91Xd1o1CD0KsPzdqP1SL+tHX4fxZZxl8NtEpsroX
8ZqppC1TOt6iwdpTz9F6cm3LDQHQOYlhYBHbyaRiSZogC2CWh7nGvEHTwm0rSw7f
qkt3cQuXztYNdtLLvhBOwJiPn5IRJPwJ8Np0zQ2kypSGnPjgMfEVn3rFLpXkxbWn
l3ZBCEymb3qE4iJYmyKeS1l8Mu2o6zOXMhjfo64Z65tNbmFlPlaijtDjPGdugie/
sZ/KgwibC8DR2McPfI6nG6yXecbH2JeN1pmG0XPQOjx94roszlxebMSIGe4sXkrt
4yByUz8BiW5Rok93XzDq0Mbiq7ES2c/5BmkAjawbxDM8jioD3SP91KwLwLklFXvt
m24e+IqBYVsJ6CQBM5kx4e+k9vp6T4wodEzMzTdkhjCpD4uvH+oz5stQgGoZ02jk
uaTx1PH+tCcXYsEmASJCdSkO49U7D1xqlNHElhL5I8RIz7gunbaqaK5NIXTH6mXb
QaRXyso3D7pMiKdGjMMQvxN3iaWxTeW6TjPHv9ALHK6B2AFsjM60xsnb+nUi3oSA
jr0GnrIHwAbMfXNXRErqFMjEE33+OwD7Xp3qZrH+4/07XYS4zTN2qNaYpqay5OZV
7WvGhtp2ziSEguisEJS3dn4O83EH/ZFrHddjq0N7PyrjSVUhkM8OBHMgtn7iR5m6
ghiJjCwCw7gSmRWvaTUwZ2a7cMPIw90soYeOLWoXIdlweXiMmqgFJ1hQ6UFhpGVe
HkyOrkDMBTpeIreozJ2uMCYZgQXUY0eH/DH4F8vInb9+4yq1vJbOy4UPrsc2w4Tp
uz3lE4mjlTUiSL8bnKR1dKQh67NbPO5qZPYbwYYUc23NAqFvka1FDLl5UihecVSF
SKIVIfRzu2eNorIbrYnjyR4SYhc7Ww4ykhY+DFi07oiRsEGLWGQH+5JrGjcTBzaN
CZqxhI+q/1EGk3y+UWT6F7jY+Q6gTpAFM5J9Le/PM5eBwCoqhnt4uM1SHeGIvhkU
ABg8aXobsiY7694y4wHevObYf/as61QFZyb50cVXdlbykP2ZMI+3g8QBA08TeMdN
2kwUNWYgWttTF0lfuKPrFyU7hvxh8A3YcCDxfyzmMhTSDjQy+X1vaOQZQYI92BrW
5ENZzRoeAUR9uBqA2DVdF0bmSF1IA1xW1oVQdZaAjsTJ5ZIRmgT9nT6scp7wsFRX
po4uZQ0MM+vqKmgD4okd3W4G3BxZqzsFDEjXDkkzok2cfdDcesI8I1mqZFrcPqFr
V/rq+j/VGB0XpT+FTTV13hcfPrPHzy1dW/duk2ScyR/7jC2CnsnMNUKZz5AQ9e9d
iFbJkRgxFkRJbyKhLmHyLCICTBX7di9Z9ecsN0A/voKmCTUlzZ/k0lc8NTUixLiV
zKjmFDtJ4LhCgNGBSa5vD6TGN7mio13HQ2lbjA9EojipqN38v5MpPFxekZEwL7KP
bS636RG6HYuA5QfeMKfYry4QhT1+7iqbu8XKn8MnDattQQAJzZWqrBAbJ2H1znOd
DuSUEntip6ILl70MG5/vGOzepth/mY8/jd3b8v7UsgtVE1aaJDIDH+aQkoXHlKSh
SUQcodacsDhJVC42UybosPdZWGVEuzWlmX6b5lTtXQFtIGiOUs5+fauIdVU6CvmJ
m3zURHzkxP68gMQ86esaEDrMty9zJQh298MndohjybnQ+Yuj1JxeL1Dr0OULP9VV
2ol+uzPz7b2LQgt5LPrzGTkEEF/X+KkucWzt2PpDZVGl4tzLiddu/TnOcwQn+kIO
23hy0HD3UDZ8cSeWsrJYAKot891q7mrfx9DB9DuFKf02ls2IrShL3DUW8woFxiLI
6v4mxPO16D7105gcuPo6Bqn+m1Zh6FnXDOIDY+5lOKuy15NhHc/hXf3J1ZXJ/GQ8
NLg2rvAvSSmUAojchZT1HTeQ62wK9TwURLnohZZMNd6fwzjAkaIlrO81Nb5B0+HH
S/8MhOVcmCfmCRP0ItPvgh3LHQ4nc7AtzOe3p0+EMdI4WWB47l5dtpNRL0mBm5tR
dcQZZeMA6sKT15mZqNieJfEKZu40j8SDDf5UAS88AG0UiiRxWYOxxgFUNObwYWH5
xWxeJ8GJWCoqCvq0RafKjoFNQ59mI+x1WVHXNcEP7AI2F3ZUhgp/xUNJ9z0zZrhg
GsYT+JKCQFq07kLZGAPoPdTYPjdGmg48XL7X+srY34FnpmoIBf0lCOrFcUfOtC1O
lIudX2BgFJiZ0EenOFfCkJm+rjJ5BZzTi5PzBrnd7giuHYnZZveg4Rt6RqWJb8M5
rMJBmOCgrSE2EPXK4uyqsA1/7+NvbBiuPSVAVSBv7HfGZbji15Rtf85UFlZHCnig
vya6K5p0Gs5mfkjd1flBd1jTkTTR6ilvItGl4/RnY2aT3h+K7TxUgM3bxXHJ6U5D
gFg7tzildOg1sVvgzX9qLlKUIgqWhes/oRnpzPbN2YDwoqlqkp/PKNjIQaWZA4fn
Qz1fcMKjqdw8uhp7h7fhbGssunLwK5onkwZ6aSCHkoVWZYZhTi/yxDa6knPJAbIm
Qm3uABCS4eZ7L/z0FYA8z1YGbBtFnufolnGVdTl3vszls0IqSAySmKp+AM+/ahY3
5JtyBwtmsH6DmfwtS5ip/O4a/bssT3Ze48WQTU6nCPPSfUlSDH+77JuSPi7auyxl
26/QDr8y0AFSbYRCLzPbyv8/GutAV8TbopTFcc5AVX9eAV6CaLeL7CHlp52dPuUJ
DGf+lBWxA5UtrxCoJdCqr9m//l8/SIs+eYlLmZ2AQDs+Ffu3zRFMYF+uFrjCRizr
Z775JFhkOfCkNR3hf3Gda/4mcNjBHLp0rrORQLGbgt4i4J1kVLWjaVjjN8PVDGhb
gD2nxlYzJ/A3IIVMmr0tzJpyeC6eqTrJ+AzSWCh7CbdMXdCcx4T2Ija+VlmfOev+
e4mGmMd1QQiHLYZaQMWd/xQ60sf8iKAX2ADPvOEF7IRqIsa0ZqxhqLO+eZPXvhcg
mQj9oF3IrAU1vX5jzHSDbbflCrBB5E7zINaPLC4Bz3tBb1ZzHzcri6qdFRxhpEYN
XChnCXsdQd+FGLPWAOFccqBv5r8+8IA6z4fSxbHUsM8IeDTxBlTwGRfSl49TQ3lS
MVipE+s85Fpv3MDpGvd64EDqN21XnEp3XCW291OM3mOAYltLChBXYmiFcW374RZv
FrblN00y8605pAmH2iVDCfoOMMq1GAisrSmmjK4VkTbhzfUD69hGORwzIDFGhUZm
dfoo5VRz3jE7EVkK1bdwf4pCf7Aq2Mlq9TEs7Lsx9O+N2Cwems1b8H6krRd1wXI4
e+7DDp9sHGlHfxLsJxqOkBRzJYARAxzuNZE+oZL7qBDToTHaDir46kl+faL8BkiO
nG+CJSVu46pzYdfXHIoCTTIX1nD8bBeSL+Q5AELEiD9OXgtG0DIsehRR3yFLttv3
14AWXzHWdiCVeS6YfM76Ovbw8ToLty0X+Y0SVtBDFa4Lj2Y1eqG2jheBNvuPNO4f
LtMtV6rv0xUxZ1KF9XNLH0ExeHYViaBVeORmcyqgjJynwroJ/MHh7TCcQh+1McAJ
bwk8Tun4QzDPsELYkPeSSaZCI/OxbMSlGNnbzb5R52Xx3iQAFzMGfaIa+xjpumVn
KSlPD6giR25pi0VqOligk7SnrJr4HrcQs42D4Zhp8maxEZS85C81cnD0ROipvo4w
gBBDH8Pd7t9G0alEhxSt1/pQ15lV+An6t4f/iWYdHhg6FgPoVd6Gpp7Aew1uPT31
vlilBoqcHqF/Yg8qPPQTvolEus/7EVUespTBTd5oBSOZglNZMexZx1esK0Sf/6cE
jxKw/FyCLWUNhih4lRxHWOi6jXeJVleUHDcXzUI1iSyl/32XhIuOUnimHQPCvfVt
NpQU0+2h8GA+Cixr0ZTpPwoIsdG2p+D8yESgTm4ljoZBM4Sz5BTEsgpPgRp1SiJT
NctHs9PCwdAv49+uqIJBCMEqPWN2mG9yjBhu0ct4BzcvfriLUJ42eLJvZ9M+2lXq
AQEezlhydebx9LHC0wZqJNMAphBUO7Wp/xoMIEsUVjLF0hmET9ZrOmG4A6fyiWsB
c5dU03hjCYAOV8E1jED0TZLCjFjkMHEc+dxHoI2nWipd0ksnjI2eLINMSC8twg2/
3O1ToVyalB9WUuOM2dK3GACTrvRWN/wXAS4qCU7Vro1zGBurv+0IPueUUOKXA1Io
ebjIh3eWYsnz8xX00TcbWVI8cmjlFGwIX7o1Cc67XsECIPdTsw+AjErxA++o1uPH
rg/UoR5CnpNfyS9c/akn60T0L1hxZrR96YTkMTZ4kswBpwVluLubkm+ESW/1AJyO
iJYd663bfYvvUeGSawEWkQ6xiv3XSD8S7e26fIYdBdSUQfXzMeLqSAKa5CwtBU0L
NA/XOo0WVN98daglIogak1piyfeIq44B7BydPXV/wa9qth3xrvicyHYpVoQPB6yF
OyQzCbHWa8fksn3Durss7fwRrWP3qf0+xSdwRcpUHES7/Hi8xVy/KN4ueptTd6cc
lbq/L7QesUej65d4aaKDuYk8ECggup1woL+P4Tdymxx7lQuvBn8u2RjmH6yBTS2v
wS6f/+2DQyTsagCo1wEIFQ1wNB8Ai0bxUO/zsbNegmnWO6pOLf7MVnvKBrSlZ+Cz
a7oOs3s209rJRh8HSQlNMW7gVtQNjMx4wdm1kEGuXIZnHTKXyrzIC+Ef4SKCdQ+b
b4l285mxa0ILYhbRz9FKzon4HvPIDzKMj6PWmYc6H1uOCXSS+nrels6SJKNwBnKh
8V3IVzp7r22FoBi5ufBK54BmuMRHxRIEoeE4VcOb4TPmNQFFo2ZdItISiKaH04IO
g4Q+7wQ6hJMbv5NVKzTncQcOmVFBQ2cMBkGj4zij0dBC6KHEkXwkMawoqxA9nVfI
eDcUgm7fMpUIMTOZh+yxhqOV5UZCJjSKgxPSKuMQSwP7J1MIbRk/t8e71wCyNLV9
KDmMdKY+Cl4i1h/bKpPr37NafO3zHGaeu0K/+2J47j2CR2sC7tgGF41/lmAGs5QO
e/yNOBRRXNBBdktD3/UEBIpqEJ8oBDUuLwLMxPxWoaTAWQ87Fnbv4C+wzvLKh4T7
5QFGjLBmb2RA0nKU0bHIymwvyjv/PJFR3pEhIRg5oAVZgBaukJk1I9fnOtl6lnxI
ZpnUgjqiMi+7cO0dt95oM12cyrofVaAdv0Oo9swyYBHLB0BEHGJia71YHb4hDDXK
Dxpe2dOmf3Q3oQZVihuxHSiylhx4brKOK7kT4ZD0YnkeROj29sXugZjNW8Oi81f9
bYqqljH7bWt4o/1uH/z038y1Ov0/vCpS8hJ1S6QKMjJRnfE6wlc7vIHJyugzjHzs
VyEL/6KuEUN85RVK/6Ck/3HBI5coafmDeDpsThh4voa3snaAduuEKcU646L8peL/
6JewagUpXE7XrL4emzBfHQpwfMUc7X0Ei6gpPe2f7C2QvLs/EQt/hQ+ROw8yJfqM
KzXYthDdvZcNrIzKhbqdsSzFDvZF2uxrbzyHd+flv49BX29xaOxOSPQ1NRWb+8z5
YK4or+d8/DaJfA3yaKB/8CMUVhC/8BdyNHpb/qxzpEHANrBHQUKC4RSX7XZURcIx
X2plP0QHSKPDGWY6lnduBuEVkqP76YbgFrTBE1YjYD0klQdEMuoa3NJqADz41NNU
oNknUkQ15hQcF0aPTOA2gAF+K7spwI0yMFWEDr0SF/Dfm9ub1/LjTcN2i0ZeayQN
oG4AYTrO7NlkvmlrMrl3GYY8TjzUEHB3HKU4n39EL4RYNVLunu/qN8reMX7q6YnE
ACW2nkEmh7dAGGJoWvm3w+LUbVeEpVxAnE+sNTAgWtNYVS2qznBof2uXPjTZr59R
SkjA8B9jtD0mtuTB8QjcaHCt5bFSWqM7wTf96EJZKbB/2PgJTfnSyk6caupzcJ+M
o2NROgdKObdQ0cxwzhuj6zQ+5NtnCNMQdckwzt+iRcdfWJWJ2mP8C3cCPh200KCQ
B22r0kFbOhQFR7NM/aQqnbXlYp2NjTWy4R10KWmXIHimWezwFkPfIRwhxgfFEeRq
8WKHJbTCcoBk6/V95lSDqaJhU1DYGB/646T7pMrrYr4zeR04nj3xcwWurElxvKh4
lWXbOgxkBrcnMkDXfYfm4ACkKgHBQZkHjHXMsIOqaVV/2vmeyKapY5G/93E8rKWA
GISZAsTXeUSpfKQ6t+JMcIwviYUoBvQYZ2lYEQyvO01M3iHeatLv1hHeRKuDACgH
rUmCN4UhQvFvv8YwD1NQCESOANL0xYehK73dcxmkY1Y6XzX/CxlNZYWU6ppg97Bw
UqNO1ID1O9zLYlZffeox8ZQz2LQsByr+OgACFH0adeAVnbZBwhJeQ0JPhoT3ZO+z
NtYVj5FFhwHMkU7x3Ni8GnGUELEQeYticoXBtEbB3PPn8p911Bzoo1CrO+13g8Dm
j9tahHxlX9GJA3b6uyDVIaVtSyzpzxwB3z050PLqUt3Z3j7zKbGkrFHSfzRHPjyZ
yFtktvMZaMT1bcXOEVkAPbO4JM1Stt3tu/6KHzegRrwVCGI0+/cVrKPqNxz3Pztv
4wJmeeOt4EsZOBnYqhyjcl3WZ0J3XvaZePo7ovsldR9NUmYU29NLm8QQdGthofpi
w6s6/GnFLW+kxtTf0tYXKQmO/2Ja63i2zqmynlSk3jzMnccRwANCg22AowwCzZ9r
2JXhqEm8Uwoxa/tbIPiwp6UjSdID9yTejW2/1ehK7Bz8U6//j6/Q2Gm7hT9ScuAi
dEM8BZfnzGkwHc0B5ifaP5XMi6VzHBRdMDvOQTIkuMurZw22qQDDSzQVunxSLgXe
be8KRpthpFz2pF6++oCBG6ESWd/EVUE8ck+1QVFwbf6yzGeo7tpXkyQEHQEl1nAS
vi9LleaxAcQQw9l0RE9I5h8kNB8vBuCL0Kv+aXdmiyipXQ7iLUlnx/7uOoYO/VXn
Mb7WLqF58gZtnTVbmzOJC7EaNolGIe7Wl3lFdMUYGqMW+pvSy+p/jOY6jENFjLTv
0Fyshhft14/DI5ZRii7PrlTO/vtar+b0XEGkfU63Kx8+B0KFuLMCAgk8++8JIoJJ
3xizqPArcIMTvSqzPLzCB15aXohjIxD28UpgveCKF/AdiodYJIC768tEpn4ANcjc
u/qP8oobz3DlYNkxVtZvZtMMLR8ro7YOETguwisE/sFK66rq6rNY3d3sGaci2OCj
RstCFCTYb++DsfB6YH/KjrJ2/9L/TYzyZ+W3fasM8nt2+4ZFihQNjTBRFH/zH9Oz
ptMXK0Yd3hqbGLXvz/IcWYMOT0ySV/WKS/Pnwvt20iLv7MfyW56ZBcpSNIUNAJo+
Gh6XsiStSLJ7kea5nA6BW7IN7YxeT/1/WbAkBRSuGV2Zp1WA7XQuvOZRlb4dZNh7
Kdc/569GMGEm2NLF5sc/ykJelj8Wo2oIPHAVAuxhVsL3eJz+klmAAZJCVkSfYXIm
1btSKmMNf3PlpIyE8CASz7zaObIr8vDVwHlmJhhQ7T+ubB6Car3A1Z47+8TC9Ac9
JEGyvNm634p6s4m7lLsmlL+xdB6MC32Xz+5ztWWZiPCEXerGp2ZBSOdQ2FxcfpxP
eClYxKWpTPhd2V+R5GCxl8ByOFwwIx6ubKMqAkbPrbmMrQX4bbuEK4dX82OJImSg
ESSjJuIPeZsKeOaDs86/FO/QNnRue501RjmvScHWNZF4y6mSu1nSA5z2QaiN2Xmj
i0QsDlgsOvRWqNJsuy1VzKfg+0ht7N/vZMx1gN5/uvU/WSZ/jcKUClHXfyAF5ugj
aV1TswxmqnsujIQUqXne+AhN8k6bKAxFpJBp/e+om2nF1jCiHgbtek3/bE+plnx1
/hx7NzAKo+WQuWlwKh53Qe+1suir0WkobUJRkbpGhuBavaASflkoN8RxxWhISiCq
+xNQsEJXcDMVwTYUyd4ulrf5e/ku/sSGXKtpTwa2UDNnNxwnnZKy7iUN6PG3pYkI
5i93lDyGCw8H+ZFn5B8JtoAXyI7M/FakmbgihIaEsYYaHWkG+g7OhtHTzJyznsdX
8y+5t1X5tiMTL1kHZ/jq8KJ0vY0Xx34S6V1tWpySzWGNnA4sjjUS2RqJrjItKTVT
rK4n6rsdo92ItJmk/Sv7vIRPyx7WQ23P3lYZDW0VTzuW8o2Q3MQXKkK+R3MNEMU3
o2UAgRmqaq2DYoOeyWwm9UxehvreVtbGMLyHBubyCgzIHK4/exNYiF9zDqhYT9HL
R0S3LxmPCU751yVv634Q0ItYPSMb5H+y6/++N1zzNALRXQ1j7xTmY00vEXOwbr6H
6S8U5qBIrgb5E/qSGfVFVug8ihZev4wdfltO1F8NaYb8yOwkw9G4X9UlpIO+/Vvd
yiSMl66qXVAIQedevr2Kafl1zC6PBQRVLsE2i04UfIhm8hOivXuhUb0IQZVturRl
mAtTIG1882SsdDJHclsJmxtSnEZwsYvEdBpvVFYQTGXTpSyJmGJaEM+BNyS+Rpco
RvPjhdm7taC4iLKKrfrxhuCZHTpCqlgTM8UaxQ/kQBw6pCwbcwIFPt5xge0aem8H
f1vOV+KalpP+2PNnkuBcqwEUiw4QY6QVoQGfGyuOAv4b1Q1khkgMiec2ESPWvhc8
wcJW+LOkqpNG7hWe2JT7UPa9WAtPKlGveKlLHDzuLuV+lNCTEljYlCKrv63i+l3/
ScFk1CXy7ZlGJLGBDUnQ6Jcte+EBwynlq1MslDhtb/rmlO3cbap+t5j0MpP45eTG
QtUN71i+rEyqWTqTcsMovwehZIFCGvjfc+xeEZ+5OW7v5MaX6Ppc49po6aW/wFet
lrngmQFi2EQK8sSWG29Zmp4jsnhAlqeFc1Mb36x8BCaMOMu1ZZOP09GhwRX+fIcR
OPALIgPVMTaI0mWramNlrz12Feq1BK5lyo0jnlVitneFbPV69dS6kzDlDNKZfI5N
q0gkyN/8DzSpk6m0Z6qAgC4ZOrT4j8D2B5s66QtZMt73fQAMiOldsBNxPoe0TO2r
7ezVTvvkOZn9YgTdodlwgFEXUk9ene6FBrykWwdC6zlhhwUJlltHKXbLCtHxE+pX
C2rid4aSQwwvi6OhATgVrtytVlWFSMxvJ9aL28wdalqftY5p0myHf4phNoInkJ/B
RFaizGo1DAKvAWG0iC+XE5LfwKRWGiVNzekx4RFQUr8TAG0Mwca3l+2Kic0eqhSh
+9X7QZG1PvPtQTyYtX2LsDjPm70TxXU+zpjguExbV7fEWG8V7LjR/SVfbcfBV4EV
gdQ92hVny5r2Dx/Q+UXaqd7ssDFN9pTNJfvRXntYpICWTinitVGBUzPVvAG3b4YG
wqCWVltHd1s/zEl1deKtYiL07z3PjhUds24NqCtDJztt4pjl9xkn0AEC9Tc39l82
CgwmkzppcXdvQaovEyD2Y66Wl4JKDTn+0nRsmKqs5cFUGumeY16oEBj0X7/93I61
8BVMTnbN5dupMYHh6IqdoJufx+e7kgZXDIr66UVsvtyULWB2sMurdYAdJaeWS0vJ
xs/1qjG9gie0zHiUpBseerfkQPbYsvYq1x+yPO+9LkJvAG7eCsHdX9AWdxIS4Kxy
4x9MlTwDGuz4gj+VnDVkBcbiJIsssIlrdtYyl8zwC5H3dRfBZbBPhv89QU+c0E83
fQzkkjHVXFG8IKqCx+KX0DXXoELvg/f2l6APsM5KoDD7/ov7DNpBOkcjOY1VRMcj
S9db4y7WJU9n5o56z5/mo/aKeCOOrBT9F79olslp0jmwDIlbvBe0z5QCmiBDzw/i
u0E2yNBHv1LOIhqbu5wzgIh7ajcJGE9FsZnmllinqAcIb0x68ELRmxrdSyoD3FNj
p8l6Z9Xa2JbwQqVXV3vw4wkee2TXyiPTD8L+9Sin/3nlaLudBB1FEwvePMe3U+tW
1hV2p+vt9o6btHsKFNCnrgSOPaZFvaYvBBUdBr2JCqjsMJu1zZZ+xxiDIDj0zun3
YEPT6jlsT5NnGavzWthNdSietA7Qj+sYOpTCj7K2MMIJ4v1OTmpyIsKfirLnkEIy
DO1lOqYfwPZ4tjXyKKUUutxqOdYDHTBiO4mP3TMHN2zMxHoskyTtgkma92Fbq7vl
OKgi1Vie8HKrlz1nTnbZrzdNzS9Ws1m57LlORgP6/KhrqDLLax/AYTnIag7f5nrL
VXRJZYccems/AheUA4CusI+9AP5FAYtiaFjEoxEulf4XZ7kmo6aAJe69Jsn78HOd
JXp1Jn2eJgqeB7B07Ij7KsLTmpXZyRHEewruSQuJ+6txUeR6+W+CJH3dUti+bL7E
3eTBB4iY2f76rW/ZgMgqckTMa9YlC6lgUsgcScmnycrNlAqu5g3HKiwgAWHOecNx
QbE5yeLFq0pyMj0A+dn14pagvvfOtcpz8Rm39FGwaN6/segJINVaw/t7buGpmCjv
0Dil/p7iPQq40SnVN4cryz/yoSk0KUbby8a8chHNJTScs5IG2TDod3pdrJWqazrb
Uo2pVPRtIo331ah++eJk5eI4HJwY+xcqEvz3ibK1XxztN+7ZbzQuLJsthWV54vU1
zpr8GGoWessoGxwX7kmNF67AiUxSjd6Ebwq2bkhluc2x+6zM3CzQSoA3eZ1ndrx2
0ZpZnbpwS23QRX/plEB5UhUSswyIPoTErJWnxAfYswNIKRsmGJsIWcrnZN+HS+9a
BvhYYcEc4dAEy9QXYiroKnAum/OfDPpqilcnzRhSw/jmevdPm2rUjy9phSnYp+WG
mGk4WUjk3g3RBDITuDrhqFFfIv5gq4Ji+1jVJw+MtCe1cDRYGV6q1FLDEWF25XbK
qzpKdLZ69OiJh7e174hZ47XI+kbKuqfxtwyZeKC4d+SWg5YkL2FOm4JCyO2mUyOm
Q7SkSRBeY1+MMhrEQCSncNcKZkQmdVfhN4DrzJHycqrx8hzEd1qMf1jBGWI9apZl
XuFTpRoIPtFEAmZzYUvLNemP0HmGeWHvzMY1SlaV3vKELVnFzpi35g5z5yoSCqC8
SWJ4+Z8Mgw8Te2FB6l/RaCzIisv1HjPUiu+4BAwD2smLRyReEtSE4nrix+0ua89X
8bo9Rklh71KPfVg4NbOLJ3TFB+YiHpleaCg9edhtT31dstEO+JSOzCdoXbsZ9NL6
i6Rh1/iItiCoCrtjdbOkBF/tIEnG6P03TQcuUGCnzs9w6QPTi6WqC++mxgTMu6y7
/8+i5scKgZ9T02cbNO+DLY5YpR6WiXo6Ih7xRUfstvvbfF5ld1sqVqEzOWPLqm/O
Y3cF2u1jI2nE0Jw3CQoE23H5I4pn9SNc0/kO+x7okb8Sz4QI7xSb9yH+GfUsfi1i
lRVy7nIUzXLbj1q0UmiWwdbhACRXT2t+zW74VDEmNSvvlsaojXDsi/vNbqbR+XVC
eD03KMk3qzOfU5XBltza+sU1U32Dx+p62hLa68x7xctBP0FMxu1U/RqcfBwlRWZh
q4hD5NR3ygZ7m8SijXtQ/425o0HhWqVdJEmrqI1OitinJBYLAz8u6XgbXbnlDDe0
5YUix79/yLtNVmERi4tNH5Xj5fve7cS2YmO/pieR04lTxHcNhZcPkvxfKZQc3kpJ
ubqJ6YSwkdC742jZwu2v7P3UGk9V1IYiT90TSp8lqcqbRy3WSxRXjj4nIv60wyHd
G3+jPwQipb29Si6XI46PbJTeh4GMcKCtN3tjhntb4G4Xg9zDObKFgbEwfYJae9rO
gDcn+05G1ck1ZZrCbJCcT4yWlfLBJKAOI2nO/dJDlt4u45FWdiqZXBznfSHGmsRt
/hfc6n2zI6YSSMn7FqqAOo2eLiDho3WL8xEJHcD+mBTLKZA1Fy7cxnXE0rRkZqDG
jp596JtNhxSZyxzeDsGrqI5CuGferTZ60dYyt3ihXLFLDNmI4SSTqhUOSaFS2rkA
JfPT9bCF0twA3g7KrgaVHbhET2sYtD0DctmfENJgjQ+6XvB4+UMxJCUaxzHa2KX0
Ly6xxVzprv4yhRMbL4dh3b7SjGdApjTDp7LN9Rqge8D1cPwQCMp5lMcDYTgYPPN2
Tm5prLBjKIv7qjzFWO4iiu6ot/IyuEs3QUcE60UpJqyxbMmh4q8BfuLxzPn9EHNR
JOFYOcRCDecJkSq7Z5UIdnkpbrkXTIJgrSU9BMf9JvBGQl5Gfw8mBX6ww0S6qiDS
UJJSu8YRLFnyYm6D413k2pXRof0vjXOPDzsQH2cFtW4UpE6dpBth3KyUvH4xYwqK
mrgL0CfwwlRGxP6VJ2dwXA0dZmiy0rN4FCPY8M7KzFQm51fw8O44y/SNOAhw63DF
ZzA3TmaoVTFflsRN3sMEE9MgAaidMlAEgo0UEj5SAcm5yoRMXtGo6c9qUpIQKDDW
NP5YRJKknV08NsE2kPloGklUmdfMx8kscdvohpJUghS6ehFrBXAeYoKtLf5QcZQi
hUClcgZHQoJDZqV3zdfapkqqfmsKnXtSJNvceZ4dTPsh7LiJdbLRQmOjS4iW2fy6
+ruFM+sBtiUu7LPIzYtoqTCgZJfbn8vV6GuKQM9Rs4yG7STrQPYeJnY2eo8xoUTn
KmXP4JHM3X9GumH4+mt0+dascFV6oHYjcP3oHns4B98c+F/b/YWjE3lxh9RsBdWQ
ynR42Rk+/RHwYULtXPJid61XpTyFUnN4LAq5oplgZJIG6AvegEJ0jAOZdHoN042b
JaT0K146g44EbmFPEr4tCHRtFrm7PTlFoRVNdXTse0xEsytJrPtNv5pRBsQ9sgRH
PAX+3Da83ET0NAKlJjX0cXh6C6Xsn1bNHZYu1xGFJYeFjladLJKhvVTGxlvjOuCN
4S33/i/CSh7ojIbbQKFdSXI3TroAc6F1IzapiPkZwRN5j9ZU2dtdWCfzDpEXkPpi
EcOxxQs4AMRy4G55O/w4S2ufxDQsHaAdEuVuuMewtgmkw05mbswF56h/ELG9l738
0G3hhAEfIZgTYOmDX8O6TiTlQHe6hx8m0/KxUouEIJZ8eYKKrlLTvnuyMdrNgRcl
3gAqILnHqEJtqGXC3lmkfRAxlMYl5F5RsBc7hSjR/2nRoS5jfO3ypHLg6Bkjnb3o
aRT90DSQrdRRvXAXNwQeJnBjx7Wa00ndfs9GBluil8w+k5faLI11niIJ6/rb1zee
xCUgUbzYJ13ZyRyHewqIUkx9al4T+VKxEXxnwz5Xno4TDFy5hXfeabrq3gmQJID1
Qj4FeejJuO8xMkWzaFxxNwjfJdJ9CM+6agKDw8HVtAXGM05bw4oZtDWTRMMdiC27
U8XGhvo65iAa/NCsrC/clxIbmtZFuShnmtk/wyMDxzYxwc1YiZCWCEFlT10poAOx
nIovnc8j1qGYVNyXEJ9v3jKIzNVBg2K+sKlY0DN6qEQcHqC44+eBp60HktEsAK/a
0bxaKq19M7D1uOBdkCUWv9BK/y52bl8tNG29iPHa9Vi3d5m+Z5DiNXvfbpyNa88k
vVe10Gvuxslm3JsD3DTbo6XIqHzfUGaI7aXVwyJF4K6HIBO7g2GTuHVu0yuBdvsz
rxj/IeJbtiskqjtR/xr0PZcff/0hzeVWAj6kF2XAH3gl5SlpsPMvss7chuAVq+Cr
3k4FsYJNDzzk5AH5oCLbCe9dp0UPEGd9DpDiM7hoD6k2QDkJfm+sZ5MK7WxQMxIj
PHVgaYF9qCA4JLGgjKDjm73Ps5VlNxNVy8ljtJu4feIPfGHnIz/rJ2Fzb3GrmRJG
SHItDPX/ce+eITCK78FU6O+0OYxwKZ0UcOAgrIhwRyMHNwASukbJWpuDwEJlxRTL
RWXwPkL+hqH0B6XccYe9MNNTZkUteffXRDJWAMsoiJV5Xm5cyagDshr4qvdg97oB
YutUsa/LZMqDfwLsP1BA7T2bZ7kp81dsXSNEEPnD8HOFUItdenei1yR35jbu5VyL
S09jJcv+bblG9ydiYNn0vR9F2a/5LcOP7s1yzSuo4J9eOiqm0OupKnLpkg5w8KFj
NoCHLkmF9ftBfk/rVi2xE321yD6xMCrdOXCGt6in/HP6r5S7Vq/sBxBsvhDE44l5
ecurPyEZB9+qsJxumxiKNB7O4xZp44WrexFnF0mxdO+WPa1W1xlhs+rHPQcmwDcs
DqpJQPpfK0tjYnwydztQPgfCjP98ba5iEpb8qVO2caHG+GwbM36TEQL/sm7TQ22l
n6yVrdD3LwlqtU6vhSTx2UJ42IT69PRWG9LxmDwkiJrWPnWBUuTTuPDSi5k9FAj3
8cj7DzqufhiCho7qtxoyAUD1+FjE2CCezYOZHrwK1ks4QFjLQUzTEAfwocg52UTR
Gcs4b/Y82T7fMniBfkytm+XRPsRIusqRcvUEii/6M/sbNuegGG1F2e06xXGESIpW
thqjeWtHyRqdGi4RUHT+UI7hf7Gw3MJ0GJEkoZ5S52hFtihXudxEkPQB7y7XXqM+
Keg6GHOn/s4fR5urotJJglNMyoJI6UTITkJWy4DmWKoen0Tq+PjRECUPsxoABIED
UtTbBZ0dDZaMdxB8RfYuVBUWkF5DeIUjC/CW7uvn1vUGTXMJ4URFMn2gyYsrG3PL
HtNoMlNylB3Kuq2GFN9/u+RFyV4At/T2jZsmnalX+KK5x+ZlJ9HckJQN8e6KwPaF
DdAO02wK/hGFDXBek2Vnl5cZxRium88R2tMu3DKHlcDAUIaPG/OHuT5O87sIY6m7
TP4nITobf7Pzk2yaJ4HVdFc5a4+ZCJyIB8tp8svJ6yXODBZL9tapiGhgOAtiT7Xo
ssXqn7OFawkgkTBGQUsPm57wig3TgYFLknmXfRvBzD3uRhd7trimYLCYkHTVLlY6
wk++qqEeuuXtcMVrJ3F8kT+XHI0vNJg1/48gr33EXeGkzCjdLcFFBNKA9ZqabzWq
EMz+ZNVKu8/g3io74sjoRqOcaR5mR/rpm3lujWuuGRNgTiqzD57gexodne1kkStE
NEYvN1r/M7p1tSG1O3t86OfV2nW6yvVU09jscEXNKE7w6ZRx0WADa1Fxw9Nl4RN5
AiIgpZk8fqQGuGeKUFa5X5u1pnmRJOGLivsLiz8tfMNVjbOJjynq85EGCTfD1qnZ
vt5xpQAac6lx1RMvooF8q3HsVwngenDQI3snM+NU/utyqETu8lu66w9hkfY1i2eT
JbytSTSFktw9xWSmouQckQmZsq9dl3Ar9YbDWWzv50dNf9PDMirjRVeEuGWZnCdQ
ZuEgce6E1v2BCFmRW4kIk3JBhw/sP/K7Cdmehlh142CUgnVZ9RU5JQbMADZcqdeT
3Ik3jknuQU0g0cFobSEpKNAoG9ZX/0Wi3uvpkyZvdrPvlMgJQSGBg7DATMR++cEC
4Emj5VR3RyWOwbaMS778BaD6PLoH/AQI9+7W1+bTIvh6asCo8hyTk39pbPxG0HmZ
WWsB7A701ldzLaup+chbUT7nVmVeiau322V1MoIHl1tIQm3RY5W91wbPvoi86Xvg
gJ4tyf67AJE13BesM6QE1LlG1H9jiNFq5tsLhvePRgzEhsx/I1Nxx8vhI9omQQPo
pp7AxnwYTDKkhQD9NhBwpugg9gyJP6StbJoxlut0YrwT9KhTHYTKyXOuE6aYEjwM
Mzg04vhwUcoXL936eFXv8Xhy0dvZIcOdQqmuEYSe28Q/Dt0mc0PAJQCYJr3Rr3RL
EktQY1g7dB+qeT415RqpEclO/Kf2cgyUAiQmopIcXJXEZz1HGUUFlwMwJN1TxW+8
pdPPf6rCtFwkqEfsij3N8UTRKPO96BibeareJZdovnc1ALszQNAh41v7aokzdBBu
R2mmDbmKNt1PVcNliMdzUXWNxD5MfM9AHBhBpKPfdFQ9+/6D63tsVk19fKXmXYiU
58/Y9O0iwL5/4bSgEyBPurpJSP4WVEG6oJ8akNWYH1PPTrSZ0mklVp6zATlzjgTU
Hc+oV4fJtF2oLP34rpvRbs5XSkYfoq3LZ9z2uRyXLcFzKh1rAUwK2R59VPHpyP1f
Hsgd+Z3yyPNjbXbZKvAHAdVJBqsMpfrDbyJJ1Rc71wJFy/rbvo+7jR8wUHmNA4G/
n15wAcWipKTRuS5/bJLTalzIu5VKAV/9y/20OhLn0wN++8OMX6YtfQwUz1JFSzu2
R+0k+gcqrm/M4wkXS7KkDjt0R3/SuzLxb+Kba9UMeUxXr3N/RMU7WYlxKdWMF367
LDO5DYA277RwVZIaIakN3IatEjgfHRwYclJNO56AGYba9VNBPh4ZDXe/Ot6VFv57
WW0ZgI8GuCfnVww/Qv4ZDTGliG7K/kKvLpbOGrZM4wQrGQkNwtAO6xZFdaBZxTQ8
6T7HQ6QaanFM0+vsACREXBQvAgPIKq5SVYgBbjRe7mCDARjEAn99SxbWFjFTLYT1
lKmhkxydHtYf3K/XEAgF6Qtr+xvwUu58CqK3fU4mc75qq76YHr3MQdkHk/q3YER7
ksMRbG3bydEsi9GxSXc3TMgjgBonypW84V3Vs0GgarjzlpmmSZ06znvVvOaFj+KV
5HJAdQU355JTFDX6L4aNT31Wt/J8Ol0Xgmv5OmFmmnGZoy8W1So2mq6zxWuIywwT
LWgBmArYdcLSCIJhoT0/YzrZpqt55Ofo96RbUE3cjht4JE5aMj+D/Jk3IwhVbBlq
TlCxzFsloM9Eax2Qiw7ZEI5MVAYxiApH4mNBN+Ba6VP59WmnWKzqbHxo+Vs01UkF
oWEv6hBHOIVMbdxEUPCyVg7DQuUvOC3oqQ7Q836LPF6HsmYBTLK1qQJAGjxXTyBv
+8Djp7+hqnzVWhtrIV0FVoBY/dph+Vccan43PwEcXLnEs5UZjr/UGJdsOZw7V6kN
NQN3yN720+60yMWCgUPJKIjKtkDBZk2aOsRhOEAIzNrv0Yk/CCO/adQo1yC1Zx/R
SHSykrw6GNdoHoMbojpdPMe65i7PaoM9VSbyRVTi2fFvMcUCcroD/uW2sF31UNON
4oq7Oz3m3/5LotjGgoTdgCBaxGOHV78NMijds35OztsIq5eMaBEdRvSdtPMZjFYP
mthq3xKJB0jCCz1D4yLO1J/5G8TzfeYl2KXkIhLSgxOKHV3yOi0KKkOaX0BU/ZFS
DOoqFnm5DvtRKuXBerRzop4bXMr5LQN9soQeMPNscgYzGlUS3ddoYQFvEY3/wl3f
8FMv8PE3FnV9sZ+V7zhtdPAQu+KS5zM9opQ2UFZvPykrdgPze9yzjP0CTCmsdZ5a
PppC0iyaSVD/T1YF2cH/sZDpYI6pnVlkhHX/CQguIq0BYSdU/XgUZUMaybdbLwPR
nQCAxsf1++f5YauiZJIOLWCkLeW8rSP40MRXTdfpv8aWsdxLRcUJTjgh1hi9umPr
5XcV9k+jAlYaWfKhRGdeO6Ssj4xgctERsFiqsac/+9DwSTHqSu9iZztmzu+ezG7g
5r4RS2agi3SYQ+VWbDDtY9zPRyD+FBD9jgYAsjzSWWVB/zz6jTnThNyv0tWNT+e9
w9CbvEi9V/1a8C9EN0HLcZVASFO/2CrEBMEM9+FZtDFCo+y+X2f2KY2xlveESXzE
K7LRDg/xDwl1qsluslYXIBSxE/tye9bUL24tNmd4TsQIWdvSlyA+8H/lUFWoC4te
fvzbw0wSg8z3ZuFX501xzu4+kHJy+iTdvrKd5f8h/PXUmNMxZ9DbT6LnIuZPuIFr
5+dGTeL9pvfen0i5G8GWFECnCcGPm6+Ltntr8e4+edGhQQZhULtZ/ocMptO0q1rq
wB26LHIafuRsVgjq2GVhgoCHdkAquJ5tfnB9KWiFPI9iBSp1NwhWWRI/1yC+955u
7yT+7O+RuEJENgUPjYZqbaH8Vg/Hcw2llJQema1lPFJOyrvFzdf0H2Dz+3g8aRkZ
rBcNvqKvzH9tDY4K6Z0uUnBm3dXK9AFGNPvmDFpM+m2FzdjnePzn6PS9AN67yM62
vUP0ddfU4Ufyf41b7lgy6d4LtySFy05T9qDYi7bxLbjdqu61iBvwECup61O2GA+i
Vl5oeBcKq5KrbokHIF7mMyCkEFBy98MRlfKN6IVigVcMs60OaFrYL5qeeTFxGw6z
BMsHJ0axade5tRskf5BdmyEqa739VE32A6BEvE6twLkI7kWI3CAEoJAQpyJz3Nsz
KM0q7RBtpt4zao//dEGsMoMEJ9yx5QMt6klwvRxRC4CI9re8Qfl1GtdDDCz03IIK
GcsoQ3T8ytpy+o+D8uJtLcxzhJFNcuLTS5/OTjhkKf7BoS39xP6jCjMTuCpXT3O5
5maLD+Qv35nHZ6b1+dPgEdFXjvV4+XIfZ44HEkYVPQxGv9oIFDOIJo8W3vDk4M8P
DMDGRzoxqonZUrXxjZc0o9p6+IQ57+6zQTv4rKa/vkaroaN5Eq8mm6ROl5hAXlOJ
bVGmjZr/soi49ejuEq2WukNuKauNxk3OAOyroJtBSMOAtn28nuu0wCpPHtkTrIW9
nN7Hn5dMyS7W7uPQ0XnT7pKs9VpOYyKYeaYoKVwy/8q+0C526ouA1zVa7DuGsood
yY/yLehtdcbH2TdY646OAoGejdlCjuYqxFh872tVk/FgPVHcmdhLSe4ossNdRsp2
oPPfaEA+ky34yS/qBvTIjw1fd7/6vB7oc21ul31qtlwAuTNSCR2ekxtMGuZSI36S
lTKlr27KWIPVsjLzE5dymrSuZkIEs03Zd0Uot25WmbgBztlB0nCnxlO7/SzYc/0m
+2WOzyHu5fUQgqX7/98Ht5NTnTrNSg4ogvce/Q5//trYTyHfzXdIUfpumL3BNTwx
cQMkhg7sPjPh+9B/B3DjG3uU+1+yCwIYP+9RRQMb/+VObrHlOGhXS3ieVVuGVZQ3
n6YHw/PJW7OQ0E0+XxQv3GEdtRJKVFDWUb6+dhAGiMJ8ezINreyi9XhXl4lLW48U
UxTw5fE+GOYGEzoxauG50F+h4Z5CTbY/LSXiQqyfsuKtqe7wGIQr0M8FnaX/os3o
EQenY1CdaxWEL2b9XyPxM00HyJE5jQyhrB85wwDD+haD3qJMB3U3wQ6gdrOKmGBj
a3to78VczWCo0EMJjrFxflO24NaWhYucw+A+Km++Kj+ZtMLchQ61pciZHQ/myCXr
3Q1HLjtrsWDfmvslak6aizCf4W6jlADdsZfLU5nARcO03zGaUahgIUkdwsgtWUK3
HDCkEml0QGw85BRZvt2qRXclggVq05LEIXBpYxP2C7pRQqe6JeZbHjFzXwxz4Z1E
+velBkw9xXU+jZhprVaMw3xNgfEHjjZqL9OAu70xskJ2uTNtnD4OX7ZY675X2nwn
o+FtG4k5lwj8YJnnU71ROe8KR418pkctleWEqxJThSZptBlAp2os8XBRoUUDhREB
LdxveGQwX/q4jTr2qJ2fyM1pXr6J7mbBOxdczXNw+klsYAEq2zO1lBMLwFm0deDm
xMwPvSOjf2vU13qqHjfE7koZWvoVx0RtGzZBZaAIft7BquKCEo9Bfr0y4BfYPbs2
pWXbB/z4Qz8lcjmvLJO6ZEVQeCeQaD0DgK5KU6qkFSA2H/kUhZOyS6ecajR+z28p
C6EQZU/j/rkfujp30JHSvsMB2LLjP8AXlOxF0oXCbkYZjSOsXWEf0uPs1OsEVgSW
feHpRh0PWYt51HI3IjNrYLUDQvsd23VdvwvSjcOiO634oT5Ng9rZNniwxb0JrYhE
QduccmkSycdbPFwIK5KrdfUuJfPCMNLZO+rLBEQQJX3bORSvYmoQj6raxmETHceZ
7+7BJutbWz7VskTYyHTDhjKt48qxDa4VKhQwUyWEZkNgLmmIYbm4BfhZSlbCdqq2
jDzUaVNLXrhQ0YqayY5uVp2zW1NKWfyGfvfKEKDkT64uSCSlNyhjt/ktbewPODS+
Wy8fLUsZ0fHV2M9LhUtOmVkd79nBr8KYctEA/6tOImYlsHYAtZuEyRrL0sFcisIw
lcyGld8g2XQf2o/z878YT+fGiCYqW94CxvX4cssf3MErVMeTC1JyMacd3wZoO01z
/iAspjUzllxqyJJKKIK23rZkya/jvSZf5DPnD4D1SsP59fda9IVpiULax/R8z97B
/hoFHyx0En8W1XJnTWtcxome/FPLZJ7LqzRi0xDstYkcpwf2SawXw/bf90KHnw/i
VXwL44A3N+860E07gVGC4kLHEG++amr8tMpo11UOYinyi8/RPKMZMBHUTp75ivdT
g59bkk7ncfheX/WAj4YeZwXIiYdcCEnNn51YgLoWRw/jVvjS5aO/5BIR2d4iAYkW
yILQpF9/qwl86XOs8reaPbDWTBTtmzmsASgBYJWxTPjAgoN7x7iQd5XPl6A/EOVP
ctyP7PvWnRo8GQvGZF2eJ4G7KcR7n2BKVcDCp1a1HrE=
`protect END_PROTECTED
