`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xAlnymx4HFWyqQqMSIPmjEl1H394hSvXSif2erOAf/zKucvWR7YndrRi5+QAOutP
11vpDhI6NJcKVFbgi6XEmniuFLikNkCn/sCLSsby6XyPY5wzib2xFTuyObXI9fFX
L99JTBCsVLrolzqLLpzzieuyj8ccrsqdMluqE34MLA5PQ26AJ+UVRgIXj0hDRm0h
fhwFEy1bgzRnTWnbhQsi/oKieJ+tBwpxQ2c5JQLBtERIExtesfQruccp7MJr45Bx
BQ19R6clQ+TAm9iGWj/5NGySQZb50VaOxdolff6DY7ahEQfnaITBIDgrOYeRGcli
DTU4olbaoKb9Y+fiD1KZAq5eGSSsskHNmwoG604Cw5flDTTQA8AeCalkOs+NH597
GdSJDrtmlgdA11pK6Y0GjQ==
`protect END_PROTECTED
