`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hc3DUeGZDaS0NBDs1gFj5XbfhjRVJWt+x++hpBQVel0DARJzhU/z4sNvPhyz472K
DeeRLPvbtzyZQj6GuAM2KVhfK87JvMGW7vN2KZ1RzEsJaTADkgbvlpXmE+jK4XM1
/dX29r+4DpawYqRzwVjSFqOyvnS1wuss6u8nuXXNKFPv9V0Dd4Qta4NfLx+x4NNG
3xMWiUOCmCPHBPSK2MFMen4vz+uheuN8AuRy2Jf48l5DkpsgtL6FsOLCib1qCC2Z
7j6NEJIAm+lIMeyanF1shPVLpdvS93Cc55gsapOfSsr40RptihPFMYCMwvWI1pQu
M9TFp+mmTDcaYkvvlAW4JxcHLL5NrUBL7SKDh4r+FqhfwOIBFpeCZN/73/gfR4w6
e6vMu4ufDzsbDZfECwZD6udGN7b5cpM1/h6eEoKF7AHCWlXTlqfiSZmI1TeV7YqZ
xYVZW2hLpPspkIq1gOi9L7W1eQ9NYECKAPnDfcqp9ALFPNyIJFlkLWKUo977WG01
mKLwzN5OqW5udWFATjbWBzxw95ksE2TiMrtLB20QdqfzIQdsU944+p+x/LEroCYy
bfOx6z+X7uuuwmNU29/0eFeanPJAlTtbQ6hd0OWMt7B5oXCjrg+Cj2GHnApAOSLX
Y3HJUQ3qYM0VYRaMKykAmFXjNKMcxRTme7rLWod/+lkG1e9B3wHXg3hjIkupnmd6
YvKdVFdhyytjSwTaMMcfIAPEbtZYexZ7EG8nmBnSBF4ZR7POd1eRLoLTVeAC401w
0/HaUJ2mGOvGuDqgesdem8vO7iTja4O6FAghYJhpcVScEtZjImnv3/ugWYe/VQ8P
RohH2m0rGP5DfxTUN2MZQfbj/cYDG1LZ9/agv9uueCUdI6IfSWv0lkqHRp/Pxh0z
ERc8jInr1a+5uASoEWsVQ6W1kozCZpWCQJDzMEjPgCmX7voWzse+m53DVHx7F/0t
OXAYSPpQA/s+x+cY/NnmSLIq63EeNvAPhFioyvs0MTeuzBoOnTCfrXjWhg5P0PvH
ioY/6ShNimej7aArIDpT4uEPUApyzOETLxiiVisEn9/doLLtJrGj+TPqEU8FTzT8
2HCeE8vQlBHcjca2+yTuVMz0BsBj46iV/7UjklddEpqB9pbNR5mNfukQJtBH2Yj/
IVAmbRtBJRUJFe7o9MtmZ/WdBorlWEYTRTDABO3ffkhObM7cY3VQZr+DK0OSc6X9
ek7b1nS8n2/n1QF7p12D+kRxjmmtAb01aZDro5DyOKciSj9ytbOG15ScTEhq3KXV
j4gqtQQiDT3Qioz9j/aTqCUir8MFORVcr/eAIe975PBpQgEGXpapWTvwtOMkMSCe
yThS3iaIYpji+ms8aiBUd8sKWBYP/DTLbpZT5cA3qdvftnhmrwo5zn79uJCXICWO
fCyO+f8cKG8wNZr1cqjMG+3H+1bNUYKqxJXbgZuBLxx/KMadiRolySd7qHZYZc7U
8WhCValqzSZpR+aiA04quUZsx7avHFYJ9XXfnjTY4hRPF9cY9YxEajv98e8F56z9
b9qSvYUFa3c0umcMkPTermNJ0Ipp/P8sDOMtVwrGlGdOrwnl75OAPKCKzRDyHWPB
zg4S48+TKv415rBlGFeQ24Bz3RE/exETbmCC5PMiOzgv7mlseBQ4jZedNDFbKMwe
oE6Aq2GLdVAKPOr51WHnJuBIBrYmtVVdCdfb0idvAHxfibQmevuoz6mGSfRj3fsJ
zxY1lbfGecvLquAc+Faj772YfndCSmV8MW7/twU8xhOMO6UfenN2uvJ7FdUKR+/0
VlosFhsLpGinVQAzABXF5oBvaqOYQvNIxv8f4GlhfGSKFUsHgNS9wQJCyaF2YJYH
cmYNeXLVCZonAxsa6eXumra54EzC+U5Cw+OSwLHA6aHZn+pLglOECg7UaiLWoaDN
toB91aXBaq0DIjvwyuESQpMbK/8/Z+7HDNbI4bfE2D3nO9lzlIUYmyKSFD3EPs3/
cAgVlzCvzQRtWn6vpV0zUd7fP+aREVEH7ZZMknX+jul0bIdGirDnz8EA843agP9y
UDmkwjINM+TQ9xCnQ4KnTdn//EzCz3l9czL4Y+LHODd3MuKwPD3CvxFx62SCbTCK
S471PqJC7qXzV2j/JtWOcPwkvLRfuZYU3QqhrGbrbWu9iuMHCQ101jl/jsT4sqzE
gxPKMgswMxYoSTWzmPRcbdCPe/SUbd6Lcu7wVhWn39oJhCLd0KhNA4EGBef40DNa
Qh0Q/nU+CUpfl61GunhI8ySR071DOMRn3vTNjzdFXVaQuw1eE7XCXExCGMC9IHDV
g0t2pnzfEmpP2nICPo5lE+oGEOddbQ7JJVasjnexwJYiWLjV8/7BnEij2TYtM18z
f4JaYToy37p3ShRQkVSiJ5JpVKsn3zYbzZ5Cmp2G455XPcEriaL+1E8zTjsD76ld
eQmueYuYNpVLS5j6CPdIxojIFCGx7bAgnklk0pezTOX4m4fULPZx2CzzKlbM+6ew
O1cw2q5RLnioJ5EGVM7I98EilEoWNxiZlQHJ1U6AN6w1vCmHtA30UgvaFOnafmH9
1K2xDizvLHCcu2H4NPEWGXsOfqFfyszQWdO7BrHiDuS4gKCp56yXbpVnlkTAwNkU
4g7g/gJisVloq4NE6SWzRnl79lrnhNk4BeGOC3jkIvaC4+7/xfun0y9uLzz6b/9K
wW9p3DC+AfPBCqClO01h3NDY0+nBWW145lQwdv041OwlHKEs5m9mIAmSWfVW5k+M
+B9Ia+NpKXvcVLSJ/0LWY+4VYWdf16E/9Gz/LEP1mn0tgT7KxZb56fu4HeyY1Fse
2P/t4+PE5iCYPhYPjM2T6nWdVeqNaywlpLunrCnLIIpypddzoRYfDWSZA+MjEtgz
ugYdZCJbOkngh3ePSS0+cYzsKj+J+uqtmJ0OEpEL3EYL5DMzmdd09Si8Xg5J1MlG
a+Z0CXGPcILLNDap7D18ll/9D0bWKPsjPLu/yOb/TCUikbQWpO5hdG7zJW5KdaL4
T7155/LqX1oECOQmeHrRoizTID5373lDE/qkqOrgVULSwsj+9UgfyJL0jYGA3BCT
B5LqEAWOLqjvFd9W0gGjQrp/bkhvGRRjcAe0HYiBZ0jluydVURhxITpsRToGAakY
q6x0M2qCS6rYv/aHHCO8nz6Lhao63VsCT+IkTLnxzhtAgNTDZlueA3nGJIJg0Q0P
ksBJlkQhRJ9N7XFPhBw6q5rBahJvWMxIY4HsgVYNW6Fyo4kz1S+WTTTaZepMdI9i
T5mwOvza2KC9cHHsDgeV7NSSeLwLhzZlxA2T+ECr150dZaz6UZ5mvddxFBrbxKyc
p3SR9DYYZpE+tkmXpmR4ONKmQtYifX1iClmTf0id5JHhEGjbpfS9QmkIkzlTjlfr
nJsbmcCkgDAsO76egP6Gv+QS2qUn3p1j7GQfwhbAs4dd52jREjUamfiJ84ShKJLc
mc2v4w55c43mXi/V/+l0JrDillf0eeKP6wHXfWrogJbQrbHyaImbF4uYCeMWKzJ8
sd4cy0fnGZzB38mlXZE/bnyaUhoU5nTL9uiL4z+VYvdViKVMZNVhm2EneuKEQCdp
E1QmxYFlZBzzCbZOiri5ABex7a4mepUJL5/rAm4A+jMWpubdZ1ooLu8zmyjB/6Z4
4w4bWQm6CwyaukCJPMRO6rGSa4yXyYE0EKV+lWYZVru50CZVJa6eJKJjtojlmaeg
swXx6h5oL+aldoRUFSochcvYBSo8U2tSahlN1XK2vaMTb0W5zJEIJEuIIQ1088sA
+X1kWDTQ48+dl2LlG1tIPlrWE02qraECVr+Y1SsMGcfUaFHouGU0T78F92GGfzYp
IGDNjxteahh4QOCppLRvaA7XLBWEc5u/caC3Vxzg7PYvpROVeOwhcoce+L0mzkF4
Esq07ehvOUlrmSK+KDJVObBFVPJT0lTGpKjtL+/sfHQ+1xcQTKNIzbGRFZH2aHb0
RKSkm8upEZJ37HhCAKEEBrDh8ka2Gx4jv4I19iRLWuuHmVNyjUV4fQdR+kWAEaX5
CzNjMovnIZCRSH/uiOsNfS43FLQEwGY4SYBqLMIt/vDg/AuCH1V6ij7PGEJeXrRQ
eVcgyhXYKQ3xGGCB9cgebA3Cvu0fTnXkwX08nxIwfFUom8TDdRSpTnPYJyd+IWEJ
NY5z31qwgmHu7kAuhBeyyAXyU084LyG57aqTJa7HfgEn50tFSdOYpTRvK9C4Knk7
/p+jQFfD6jHuIIhOdoALeAfpMQgVnb62U4NRevcLrKDTJepfd6KPzIoPdY50YpF5
g543/UPhatw8cRehc27vCFid5P/agZSne8gAkrkTZhcNViIYqa9qEnt5JHY7Q0Vj
WBf6877rqcmEWtjCovd79oLU3v9r7AKmIjZX1ICct9Tj1HUYZBccpsTniGgKUH5/
D3aMDsvUXL0RaPAplMjtcabpOj3fAqMfHAeT+03+WgeLV+04ko9O4VtLzlKKkCw7
DovGYhmz5bynmVmcarHaDKWcPjYfD/ncVrpPUT6P1uF0LykRYilICoInTnZ9BUBV
D2sKogI8u9CpRoaEYEKEkcLR6debgpehtdv4dxz6LduZgKB2LdOhNLueszKbQtSF
K7ETmYyjrw6M9nJ9xYD5Z8sD3mmDFthRhaRvlLs8wkOWEX0amW5IegDQO9tfsbHO
bjGneV82XAiGCL3zsgCW4+PI8/Pq5aHAayacj6SUkCfY92cfrYw1bnos5yVUyeFu
XdRP+KnMTKGuNo+MJxJNPbqkftU4ZrwH6QBRNOuxAzk8NW3h7q3vmbSv5+sDwMNb
Q0dyU/VsZZBdstK+h9x7aF2kPTKthFA47zr67eyL44b88gq/+bY0lwTSuAEjfcFo
Ywn23zjqyjihl51L7Ymjmocp0AeRqa+frl9/N5CxVEtr+3DGNl/aozpEZ31ultfV
YeQ6Z5zKxP1rsCfokG2ZzuAmO7/f1wunTMt1xJ+bshlf4ByW7F1oVWRTtZlZgD52
DbzVBsLrTA+/RHD9jBKqQONsRRUnFKuCWi+Qo06O2RJR+9MR15Fkv/NB97LzPSrZ
8z4bQkplh6Pw31ldcKXseHy2UTWp4eH8xluxp0qAQNdhMVDD2k9LF+svjTsNMYve
nRHnV/vgyuu0w6EEcn+3Qoh1/0hyyUIwX9XHc228I+YfQxFsG6r4UcGjPuLKXGbA
cg+THy3JTDyKcUHIfS90qLak0OAXiLR85YHqwfN/lt9p95tChlCTdsSSv8dCd3iZ
yBC6iYE3zMFgQgWC8QM/XLmj3lSmboK/6/02Kp2RLZ8ulqBYz3QeNPPgI2HPwRd9
TxaGUZwnRDo4W9iYA62K0J9irg6UH/4sqeLPgTHqMChS240zxfNey4UyfeSJXAxn
QNQcz3R2zIctg+eCe4YXW62Y71EzCegRAwmLLP9XcskI5ru7fohqg0i9edQTCl45
5zhfLYGaJM+kn8lm2Qgjf8oPBwNtFgdnPLXZn3EKzder/PeWPAr5ICj/bAUSzk0a
t+ZP4iPcjMVuqJL+GQ79aegpCT7eRxrX7S3jHbmDtvjb7FD8GS8k7YhaRVRqUz3d
DQOySutC2oZmb7bIGF2yuLW5l2BhTjC+QYy6lRCuTFMpu2h4oiLfUSSxRnl5yLO1
wmxbCZ7mqvp6fHrY/PjCwR59ktY/HFgIBIhYSGczfdzoZnevoptQYkVPb3nGPwTX
mtRdlnnRqLx4ESSCPoIgRcPWfqvPvqGXUJTZbikYa1X4teO4bWBMKl4oFxjOkZa1
qS387P7c0GHQ9fzjpO9CYIeqsNfFihRmurI5l1bJGepNq1vMHfQ2fbbzj8BpltZl
ATF+Y9PL3hwAPFFGf1C9GF0ISTMLa7lglI+r+dqrJtf/iMR3T6A3GaosZAZo82YO
WLmDoOkxc8atB7F6Kmx+VRRYZw+f4aZaulho63DJ2dg1M2bVmd5w+yrRy+91AHog
hzG0bMdpZ86WuPVE6btE6NtGdlURXGNj6AirgiKzh+rFCOSnCGg+D0/srdAg92aV
bdMIYcyW59iwkfBsQOFn0+SkeJyAhl7ZlCipbCaS9BnGtBNctbwWuY6AXin4JgEI
m1QK67uEyu+gTWRkc08EGuJ93vuG9X6bKd0ed2mcxGeXrNMO34bn78S5i72F9e5b
fB1fH3IP3zBpc1vwF1UZ5oQcFd1sBUXkTTdbOH2z1ctEA2fkpRF2/zeeEvitfDrz
yOMVE85LVeHmZ623BnONLGogGVaQR2UOUnZItcjFf/AQEc+aRNcKm8SJ5MWUsQlo
ewLED7spEe08wLutVBLRVhd+2Z4sPIyFCrOQr33V4ToY1VNfgJWTiE/207ezHuXw
GKnY/Fx3hQi/HWWItA40Os0IXRea6Q0YMZ0Vi8Sq7p+6awLPzB7KsiNkPRahF76w
ovF7xt5aIyIo8O3FWRAD9gnkWgssaXRe5RHmKqVHUIx4dVALLYlHX0vmcO0+lUZJ
h/E2VnKnNm+b6QN8zUVj0sa9Ezc5RDWdsLXgrGDPkWLA12RE0APT+XbezMuLsIvJ
2Oe0ebqFwubJZOPFrvLLLU9J4tlSQf8BMyQsv9Jpcpimy5uTPlxEqUAMy6t3cyO9
kvLrxZr1RR4vFF69BHoJ+txEQVqk5zmXcDaA/45VdzcNCzW3df54vXPCRYmVi7aT
m4C+fA0JLgeGKAkpBaNaiuoVXApfqOpv70w42Pq2Xh89f7HbVSTy+bsCLAIhlmZ4
zB/QobPVMH42LjddkieWNGx+uPqBjMTMrECTF+tswVLOl5cxC8RZJrm8eSDtxZfB
BhFab3e3fKbrsxGLQ4wZIFNPFi8+5XqS07r3xclAiaXqsjy0zE2YKdZeqZijdJkR
P947nLSEvkMXbCuRqJU8KXSjKEZ3FzzAOWkrhcaYMiyhTwvXsrG2FKUeTsPEecfD
CGCiPcMToNLL4S7tXmJKnMW302m+wsOdWHuFeJN0vy6i9MWwcPbdJ5XeWXtxxPlG
rUmCJqRB+7CdD/RjypRZkQyq62brt8um/oghln1TY1iHl81jmNLbmJSrTdWthg4m
otVAGi59M2dQy6ZxffHcjOKYMYuIcg2rT94y1wnCw+dLGY1mFC1wcIBO5bwaH8cy
OK/BXDWvdtSq0eMd17gf8BC7n/Zr+29ZLPKYbWdvwNw0gsaQpAPASbggi3tVHs9b
ayqNrZJEaXQU/NbGpKNb83svRqof4maST8eXH29KAfN2Gz3IVelIBw5V9JjfQVQO
icRevDV0TMXOGDrF8p4kCwSCSnubrsTl9zSZGgrFM05GWWPbeRZV3pvLRsu4hqod
i8bkB7yoQM0jEMk5jjVmgM02dwm7L4b5r6Cx3k3bD/AbgIf/QrN8gCsGXeKDme/B
3OKCfIjlJnPfFMmRqAfpz0L7x9a5EJvYUZFTELZ5JxOj1Eoo/f3etFod2zz0Wx0r
qXZ3Djuwk35705YnSFApvvgq2gbTcR3vSMNVmSBJ5ii2Ck0v5PvFva/afQdK/lkA
3P540hAiNChaApTqife3Xi2oaEU0aXc91MrY9ohG1ry7N3P3eaPQAzNhBKKCNg3I
99bV5GfwpgLMFutRKWJphIqITCrpZjuK/zggUi/vCUg45JHXC4Hc5h9Frw95riJD
YFr/qRgBamJDDxpko22u1SA6sr7W8woKMK546yhrxOfGlmlNelsEIMb5n+A617Yn
jODu6F4j5WT5p1Au91fh5OXY8xHAqUnqmqGXdtUXbeavvGcZ1XhoTsuwNciikHc/
VPD6lneSkSR1g4NWg6t+gncU5pEfq+Kz5sjzJJcw/f4WewPxlIRFVVWMlDpaH2pU
ofP1g31GY1CsLWfTKlzvibpVfDMzl68MzVRubGWDG95hDmq72NOCUtzn8N9GNwWU
tW0iXgtpOJ2y9o61FoqCrMnf/LtcaYDdYlA/DJZh+lFR4LYRB8rb3RWiqA8XQkQr
M2IvbshU/kYGsxU0FwbsXPyNT1bVxG8qQ5VdQMEa6vPnu3NEXQWb86zyvs3mOnTx
LxMmgVL/3KonkLHA2qLC4O9GB8MsjkocPcDbYY41ZlRmwoVWOSvPfAk3UMRDbXEo
c1BQSWJYNh1QbEBnz5kMA0mzxUCIhnOFoJmZgU1wEZpQPfgK4dcdtT5PimX84hR3
QCQTbX3O3eRwQ8/vdRODUglduv/hUf01lxZpJwZJZarxdMOoD6sWTk4DnxpvUpgr
64BVcLqkI3kJnunH/WAjXcZwXEdJBfmks0Vnkqt7j6XvxPCdSboAuBn6QWBIxuiS
Us+JPgRNEHeLxnjJowE4uG7whLJgVjp6T/w64wx7o2QCzFXsNI2tr+PgJQ7e6Hgb
/N+kdaRKlUYqhRGJhFE0PKuRg00eN3TYX6V3fiVQaJmE4EDQ9nVBLlI+LdWjUyCn
2LxFu/kqIcsvrTvFuVxwzeSD/A9oIPYOyuJfeiCP/FtMesbjrME4CN1NGs9ibKPf
wCwHUitCXrt+SXtxmryDfEp39Vwpv8eViOuzcvuxGKJfdP0rb6ZIOft2Svfjpl3e
HVQ0kZWHrC3Yoja5eRHae3PNYu+YhIisi08/ImbUJf87k/bh9fY2JArbd58y9LG9
NHYfiNFNfnTd2ah5l4RrTXtq4BtS0puMRGiDmKHHvslMRHTZ9r4qd85eVeuv77Dt
q4B7GSox5S/rvUQYMwg0ouDhthgnlT94PKplVSojTMzCZLCE2cx6Utf5J0PfNz0l
rADmXGIVBZK7Jk1q3ajGr7FCYlM68n4fI1pCPjOJi/cszgDlsXgSPJSTV58Y96W9
3B9yne3qdVq+mhty8PYFS60SwYPItJKukZYwvEoCEsJBW0swzrlZbDNuFH27ZeSa
JE9DcI4FzNH23KWDROKJsLZTCZAjphIHAWUTBFnFx95idgFwSR9Q+3CYOFs3d3Cu
VvVHC6S6K4fKoYqrjojI9Pwpwyhx064wfATflJKK6hwm5Xv4UTnDXgciOCKr8Q0L
NTML6dF3PqBBiQcXrLIEzSOAH43BYLsphMvNTq9rATEdKjwWvZ7Ez9nc+NfS9Tvg
aoheTcAypSZkSgsW1MVffP2F4DWsM65MZxGBvH4B/YmSYUkyNBBLXoLiU0MASAKh
IX6JQCuTXlPNC353VxWhsP0As8qYfq065CxeuwhcWldP86J6ANJXhXpuZ9wuBKov
pffsCdyMULWrsfKeAO7TOwY/H2K7X+priIixDwJtvyFX2uvAo0SX32B97oo/4VAT
FZ4D+HMBIyR6p/QeoQoK8AI1A50c6TCVC82a0yeDq/XffuyLipLqlfR8fzd4Et8X
NUZQ0uBA9tTk8gNg/sCXtKazhqKaAWpBBKe7qrFAXuYmiF1Uzk1QEocPSRoOuYxH
E60CUIkRiPlQE6bRYm4PzQJuiuV2VOqYFX1x0ZvAWdQaNQHXf7HvO05vGwrQ48fm
5VNwwqO9hfqfB9Wsp1cw1mNtSRLufGvH/HmcOn7Osrjd80TNDGi5rXdd+om39W8m
Xru2Ehffr9SUklVsxTR8F4wcQPKj9DDOHLB670TCbT9ACC5gRtHedPica+kPD0PO
xgcdVBzPeVxChBCL2l17M4XzFoErX6Nq1ckMPyjth4rhlrmTSbhoPFKj98EvpwzD
6ukYGiJVkCAP6GheDjubN6ph2JeA+R1IGWwcs3P4Pf/vGz/0FpscmZJNbEmtn/d0
BxCZYTxgqFr0CIh14nLvoGbD7kRsvoGw1uGPxPWCiZiBgMoB4wKWB3LXs4W4hgTV
jtcj3lIPTGtZNV4v9FnEO/Yz4eFBx7FGMgGCbkx6O8n5YQycIAhLEwUtRiX5qQlZ
hJVW77MBAQmiucActvg+sZUGEoOrmggklbk6wFjXT6D6fUFJL5FJJnbnedOY9QyT
2+LFuiWJ/CcgX8IS/f9Nhjt/T5D2CWJBAIfAg9jNEU903gWOarLhTQcVTxzbTv7c
CkjgpjutR+Q3ousZ4rPF1EK/L4ZnnogNIEyVSNp1SYn3+j5z37HeukxuhZecUK4L
EbZinLSAcbmivdMers1/gRZJAkFIgJo5/it7L0pUNUTbSIDcbscsQdz2ey/fIhXr
NDu1wqdUyEyzFCmeDNn9+eFrh8XII1Qq+7Ie+QVndCwbF6OlJSUo8g83ixrh1k2A
8pFmAxtJRDyVqyvAaEe89z7PCggTz/FaGUOkiKBDhB5wcxdQqo+sEZaAcHWd6k91
fOPd22RvEzQkKfCbWpPTXQGq2070bha1EK7fZfKpjaz5Xj/eeSy+CA97Ht6nt4I7
wJel6iClY5oOYRZGAgUSNBSwDKuxbLpA9R1CCNH5xXQongPtopj7Y625cPM9sIzo
tyNajd4qnnxFOy761RD3q5OUar5ijOYj8XWiTOZq+S6MU2PniGpnczoDdSdgiXNK
g/OZknqnL/6CNcCHo2x0houtu8vodII7qiCb8kRHjR0e27N4qEeEzrCgC9VqdeE6
GFEaA+TTSO9ZZDDHzhmRqkhYDEI6JAdvhXQUObHjbMkJdaNjPtbJLhgWdYiUxrnI
S3CPpqiI6a4GVmxMH8ZrprzkslzbjVAHTwBU5MKJiteohSXcs7trBs9iykx0DTlb
9kvd44wi1TDyWRT1flr8pX4R7sh9YOSmlAypEU4EjgEAhWXGwauqHpTBbj8UrSWX
ulLEQjBJbNkhUIvH45/49B3boGikXgC/96EE0FkwSz0BRvKALVYON8zbkYPBvXdn
L1XTh5Tl8rEs1iOOH7d7j5MnMDf4E6djNin2aZM1TVCiov+HuvhBoLkBF1iwMq6H
ykuXeeeKGbFE6vt8OpefD1wsqdXNQnaakucO7K75ZwgMMnH4erx7ooIUw83TQBnC
Ngp/PgfoodAR6/p1sMBpZWJ8EsTopceUCCrqBbcgev/bKeuCjvYirUlIjTjdlpme
0Jj+SIsp4uZrvwBs3m37gw5doOEl4pVfnXSSHzncZsMSSgqawNvx5nYxo68okwVe
1z6ZYRQG6bb61rT95D2qKrgXaSMbGLDJ3s8cN/7T4zP3eS/X6QR9+S5KRrqmF4D/
9AtMfJZejUsjhO+HK2z8JAV/O/woHkf+48XcUgKweTRbYJd1cAr61iyrCH6wwrpz
prP7SuWcedn2zBzNAeUURGRTRQklZjcQJm5tbOvjU4JzlUpNe8BTsk65HghQSdD3
6FW20sRH3wtOT0ag0Ww+lR2fDTQUDCuAwpn8mBLQPrZGsJ90OuKG7j1jv2AEPaMO
QwbrO5hS+rRlqQHp/VgVba2ba1541ARNYWqxxHP3N3kFaepvtwWW/qXR+oi8VX/v
WndrqTQrtPFFdpcIwVHV1ra2VfdGYcHBr9RiC8o90rEBPf48/BLgS0KE3LGGoeVG
jIus1UypdQDSgLHHkzrQCLwZWLDY4AwnPDgUfohVNdwzNj7zrE1vpy/mz5nMpai0
98E+1Ejd/E8MIx89R4U0dU2g76wgqsTcIvv/oIba16pGD27FSkEviUB+3vJmqBI3
MLhzI0ZvB1iHJrNR/2/uyCGJXV4EiW/6kH10omeV3w/DGpG/vknpSKXwfk+8m5zA
IsHWt6zME3u4DY7XVaKfLwwsVNY6WlNc3NgUP9EfwrC0t0OW71jk46pkKya8cjs+
sxbqQBw7zQ6+Mh9e0EJ++62u/8uXnJrPZe2epvCbU8dB6GGKidXjXCGGINM368ge
nBxL8OeZ20gL+79HNQJ75UjZIetb/jwcdA6ezGN7oyilWgAXlLH74gFHOyhGGKKC
YataXfMslYbU77pRP0aZkt//F3WyxMU7EYsCqFu0+oTke1AwfaDb1E2x87NN/EYx
j3+aXtPDYOKR/bPRLDVrdMRZ29LiPGAa7yd/xQop+/vvFCWce6+lsZEx2Dxmdqqz
RfNiv4mPSpA1+ow1lb7NKgUdapZjkjlnv/mdorWA4TDTBH7qy5JqCepXEQZq+KuY
nnev+J3XNFUkkKieilKoT3zGDWwdex3Y+YCk52bDVBLNOahecNI1GcfuAQj7qKdR
KCXDUuS7lk0we9NpYIuOuoRpjPua5oxzUAti5Dr1c3vOCTg4f3Qu3EyFImXO/u7c
cyGhcG50Sb9DxWNR+XUEv1owdHIQ4oIe+r26OV/LSnTa9j8IZvNnV5zQU5YWSGvg
6jW9OBfhKqG+7aSIVn2j1a58d+dmcC77FPcBCYOTBcExb7QoNXqIR9aOGtbsqiHL
gENlLKSC9TgxKL3Frl5s9iRE0rGSoNzUw+IbQNRN13C7T8VLFWZGiyXG4OI87CBa
4KfYZEP4JnHUU+/f0IA8znFWEukJSToNBX03dQlS78C3ML+IeE8d1PZz/BAF7mHH
v2xPoy7N4ny2+qkkZzQ95SUu8zZ8crFjn5Xj0PAOfT1Aruj4Xj0kDjPZ2rBf0qkn
2b2Js1RSm8sONV4Au873FYsT7hcRfhVsdNmO7PFnPHFCodZdk3uajC0M9+LelPhi
ytyEtzEP/GEaYY/z+qsAvxit+QUmPSy19x8oNWdriDWLJONh5uTvLYPOdq67Hzpy
vBMfpslM+hO5QykqVEjPBb+ryYRTqOvV0jISwMmzYpCk8VphnLPqztf1zWtpatlD
A77cV27IV3Njf07AndgAkw2mzikt9JAISMFn7gV7o1DtKWqZSuBYunCyFAyA1ynb
BZA9DPK3ZJUfx3tSHtuHHsa+wE97OD/yXYIHnJrfKHrhk9KgfuZ/8W5B4q+duQ/K
bBTsJJjT6jABHj/5MS6ckiVo/7fqCVA68ovRyCNzBogwaBsBcnEuvgEeISlxDWQV
jk80XNvoB2OdRr6LN/6J+A9qWN7aPCi9Jgb71ZsxXAjP8F7Ma+qAMphnSylvcQhK
+8JkpWkckXI2eSs0ALoMogoIMvN2iXtI+EzB40f7bA1M2vyqU0kZOMGPP0l9B8Zw
qiBEZpLgZoXJzRnKkPKkqQ/lgM5mmfu4HMhmZBWDq/golvrE0Bc/d+oWqsyxXYhe
+Zs4qdYwaVLV8FodLaD40NUUgJ9T/+PUU3q/9O0981NVxrbvAoxfq1cg7dWwDQLC
SDQJrKiZVW6tP8LhE4xT2If0/tLl3liv6ZYkIanL2ywWq0J/kqIlooi8sLDsgufp
bthr5JoSrfSO569hculUuYeJtJKhGyYtIsFCOrHsr85WSd2WG5tVR1JTvIFAziEQ
SG+k+6mMG2ZA+cBFhDIScOAUNYWnmOGYWmAhXG7YUq1tQ4uhPmcL2QKqZ5fC7OVT
SLOuFvbJdmOhE144vTJywiI79NkOeFbOFeNjfzXyd41oXCWJR0MZvcCpYiiTo5S0
CaID8EaEf6xzCKJ1fRIsQ12tY597E24Anar3zSAiAHYraUyQozSxMNhaD06cGxEE
+OJEMPdFckcWv/4IQ9fPUb5j9mWmufPXssRlrYHdetOGX1GHrKmNGgcfphju2Mnq
kNmPlULGIFlO3fxDRi2giDJG9YAiq6l0Y3YFjfsUxexQ6Z5sGDbyoAyLD/wd0yrj
QnDlWO1lb6J+KeEug9RuFmimRUQmlK364vi1C1A6AR9hf0haV/FMYMc69QpE0tYA
mL9b2zwezmFUsCt/F0EOtOaL66S2P0Yqyhxs3dRhw9LAb0vowMhf8HCVrcUTZDxc
qN7M71ytUx/ggTkT4dQb0+3YZQ7GFYcyJl/G2dqZl5F3vvKxgNWAP+CMGY33zWum
UmqREw12LWHYMKIT3g2nGMoSLJNrwePi0bltTBDt51pp9W+eXXmztM+4S2/5x6qf
EBYZTAFzQZOczDKiQupWnSlRvF5TUiS+ldqAjpZak3bmZmhuxLCeroOXPsULWCDw
wg304ePmDE02JE+0NcLWwkLrXGEUhV4reeJ2Rhg6fEvmlk2jqWQ2qZGOKjNhvPZy
oqiL6OM+oI4CYpCLO6bfSqyGL4ua8U86ErVfUsQR2JPXsLoh9IdhqIFMj5fqUXm5
tPF0W3h0UEdL9OPTkY8lq99WW4uBtnkW/dew59eweNv9FHqAk1mTzoKPWebUMDGE
71uFN6F4SxjgwkeRQL9qGzYkbewO8MZ4iO0KpcVW8c9yaEgJ7sBHnc74TUNZsSTV
XnbdEur/nHxafAWQkU74x1cJYj+19SxWNxD0rJKsAY0qxsgSU5Cufiyb3PmxrkJM
HmvEDwe/PYM85pbo3SJnHUFWqKEubopt74olF99tfeOF5E+/a0RzzW6fgqJ4Pz2F
PF7Re4nXi3/1aKMqCPHA4vQ6FVFSZUrwgy0QvMJXLWPKssgRXn7tWypA6iFQNxiX
fFar0Sq8lABwnYO5fntq4zNWhEtew1fXLidOT4gGv9Es2qdizUsEqtna4dwvfuZ1
i6r5ZPV0rGP/rX4RCIUWSb2de5JOEkACK9CnoNUEOU7JTqrfs+oXlCrOqSP3AOwg
UlXtE0LLY/9dgjq/VCTVEX373dZi6M7jTRGRTRzI5oEn0MCnD4ADnNaMJwXSk4AA
+/43Z73vc5U6EUkXt+UY0FwiJ2Apx2R1KfaJfHF2bM4m2O/G1kLVSPJuXYdpKWqq
w/Q+Qj60hfre6tuU2wlRWWq9aaGw22kYoqCKEgQK2BF2Jh1RhyM6I7GjTkXSSc0T
BidQsF2fBIrf+JSZTZAFx53aJ7xev9S3hq1g7+15IZ8ymbUXxeWjZTGLvtMr9Jfl
igXMroB2pn6meKaRxdoWPLCMzQGU1+Vz6hBYJdnBqlGGefhbXRaGlL7PM5CeJylh
RVVV3qCLqnjWKFkcKHd9omyLIcAqSXwCnyvXe4W4md0auaGd5oomE0ptK7zSaez/
I7BcPa+VIN+lNnOy3f9fca0KT+DwmYEglomcpgU91/DcEmsSNoTeeQ3EkGzCUyj7
qcelCIFOycB3jR/N1Yne8vMnU8bpAF5jukofbOaQ47Inbj0hJZORSUI01PqfS8lY
u92ij7agObf9UMoVLliQdtC6c0tKh+w/lWUfk20SM6K54Wt4WZzxf/5u0xoYQz/N
nXA9wvYNdU4qC9zdAyfnFflZwXtG0HGfnNMY3ARcrZN58ZvB0wdO48bTZlbS04KM
6nxJ3M7hyLlytiRpn1a1eEF77VGsZgWjyVsk+dJLJQDEEl5EUmQyuxScLz6mUzwm
sWv295JYXMjrWOUtVtWf4tZrtBi4SzqrOyrm/2VgKqSaM0Gom86fwHKNm+QVxHty
wXkilYKQLFv5Sf91W6oiRVufZd8rC0aErL8Heyn8WR+XYm6zLul10b601CpX5mCO
Kr7qaZCCMFLnvdzHNT8Y0ClQxWR7z8ufo/+1vA1G6b4UbUcG6DndWTWW9l455JC4
MYV22Qkao7NQrtupnjjQs4j7ZnS5mxRPncpOrhN6wXDMrEvt5pqJhB0iXfNZjVUr
L1fJ+9Aq5Tpjdk1krNnyS+PFPQ/nMN329IWmOu0MRqhn+SI/8H8EK9ekCNy+KWak
KOQ8ZXZkxjDv5FCO4EvNu+8hxXsSrY9r310BtFrUljNxKh1XWkjpg32CtkfQHoK9
AJvWzEj3zVa4EHHVoCfEQxYM1n2RZyluqX9bJC06Ym0ADpJV9/pLVJK3AQ/Bu/MT
1sHCR/ZF+h9jfLeMHVNfBHCj4nOjJOPqRl5hXtDPRB3rVlbg+nHe6p5jPjtb6cwA
QRmaaH9Et1pG+2ZK4Mdd6RqNYvgRad89kBWxGRKs/Swt+r67cuAvao5XMDVbf2UB
IHe065ND++JWxewd6RDo0XLHTaQjRxdPIxpi7pc4bAHZ+7BwyIV7wDOpYW+lvvac
o4J87CsVe3AwLidpsgzLTNwcH2qVI3wsAwfvIy46yqonuZsy48Vx1E6db2JoQSl5
uOwDjo9OTIy8+jbrCXlZDk3kM2Yk5xTqurxH9jgdteVKxQtVh/GSskd3ezd3Ko5g
gG1wChoN/d4r36N+mybDcak6YKHXnRTU13lQ1Xopdag4zxUpm9CuhDGV2IR2/WqA
vyToGQRUQt9mtI8/kvMFKSztJHZ/w/5p/ezKvSzhbvyB2XkvZtdFYGvYMHbyzaQe
NyFq8bnpo0szAYPYSI+V40gXg29Hbzc7LyxYB7buYHZ/TSKIzP8xAuKHGrBj4SX1
lZTfD2+gXR102b1RzIPBXfv5RwUDdyGUY7mrFN/8/1FSZe2oOkJN+zZjGN2p4BBN
iTe14KLmc6JlJrpKpmJQ1TRiReKm21g93UZFnWmI0Ue53eCH0qNX4DbSPdzwYYtf
Fj9sGpxjPxBKm+tfWhyxQlxDJ0lrrHcluXJ8ROxv+sWyNiV52AkFAwjvnQW8+r/Y
pq+95daOfaKdRf+UdDjiJ8yDeYWVBGC2ImjlMKHOo0e2FyAZbXQo83CDwPu9W5rG
Dl8iGJ0vaZw9MdMBhYxlvP3Uq3yZfouU1wKalyyl4LdX5JobHl81oxfV7s5JXMMW
WyipNT6jcg2OLNn+2cHqcW/3E6IcR1o108tPhY3Wyk0IPzCp12riC+Hw5mBpBNbZ
+pZ6pddN+f/QUfPY1vculuO5yuyyyqDKA/1vGsRCIVIXhx3F3egHQXU2E3HE/CxS
TwAxS/9S3Z1w0DiJAdwNeIbkYH3W81jD4511j3AQhLIP2bFft1GKEjg5MckiLVOu
bR4KsNWXgeuajPrSvmQwVRChkhVjJryrNMA3QsTjnLjiDdCYzMpYZRJBXzFdt/49
3zrLXZPTKBDXezehv+uqF0kY5MQ1QBQMCeC0arxZxW+3+NlR638TboZUUEN6AgUB
L0mKSol/hD3T/xc1+fPFrZtm02sF480Pzu2xj3aaC+DgLHm0xTg5YJtbSOAAn3iw
iLyO0wdfitnHyJLHlBVpxy1NSOx72yrNuM0bPefXjz4khHC1y9CcfN1x4u3pLcUo
NB2QmpKA5MGbyRM+SdlN7kbsuWaoBTWrePrEqyttAleskHSjRTVLT8Wpc7uDrcps
S+A3o7oJ5x3B9RGp0fquVWiUlZfqHzBwsgVfH3/Ba5T+Z4Zz1o7tsRExR7gP21z7
oYN9YufcDzISGGAF9JSLc14RCERQwW8/4Z5v947gaLeBHsNzth/dOESmufm8W+1M
Z8Ou/6p2zLcwqXz4Pnv7ELcQqRBwJdEqiIdshQAwGGwAUDpUJMVQM1IZDuv4Y6kX
kr+KHKDwSRabe3pN/cKBASujRhWBB2a9lrw7fwHXRL+p2Uga0Bo8a2ed/AvTwVvW
cjZRAZi4h5JsYOiRiq2hG0fwjaYhv1dBiBbQIV8YDzAVZR/rIqLU5SQcVWaHflpN
Yut134KypCIUxuvxXLma3s0XyFpAkByRj3EFC+ZyLeSvvN5/oDfEABhtx5sqZ8RA
Yu2DJ196p2W9lOmRfcacjCpF801mGk9WL8AhxWNmr04MZlJVk7oNGwOUvIsE2k6b
lWkizwCU48vQHv5U8yBCbbceHmE/5VaZLAD3aaxpHmauVlQi8QyCZ9m2l+6jYwX0
gA5qv7LufWBaC3HHAP16frBQJbMOFcEB42CRvYVNAP9dvxbJWPLHLo4ywbLAybcv
W6NG4dEDFEgCe8wv09WUY40dkCXr9wIlNcQcDBQhCuEchmDov8gPJri38CvwYbXH
GNeKI9khWI99NcqdzIv4cLvMZkWQ3xPtsTqRK/0mPkrmPO22q7ptzBu5esBe5Tm4
nEhWYFWAfMZnfEyJcYlVwpqRnxoT91s6cUR7y3daxAf8HtgXcRQuyR8YpIC1XSRO
tcZ5FmnXPs9SsKquiMpWzRCoIa/kmtkB7cNOfDX9sUtC/ZweWhsmrLORzIlmu2Sm
TKmz5bJgHjZbZDcWGW72afZrmPDnWtMT1on/8J3LJv9ALQT4HJWLMdxbS6RE8kdG
HW9SPZXB9AWvwOmwvQGaSQiKUwdF2Ic37BgvfOeif6dPpHBlmkR0Wwm2uHCllAim
dM2uGW00Zrh6I03zhEucyGLTkg2uXTCp/dH2hCulCCkHYxDGH9lQrh0P8/qQvTQQ
lUohrDbkcQHsQSX6x+LIoJjOEQ3fnmrHq3V29oQcYYQJL6xXKqNSXbHhVYs8sjlZ
OO27L4oK6nU3yM9EqTNJBUHbsasU7Enq7QqNc77AwxsTuwYLen0hOUSsWH0qCInh
FmB4FwIm05wZGUfoSqQqESs3AAeLyuG5nIJgoVSbn98cjMJ0Pkb53eCiK7BbCnzk
x4P4jZwnPaYPK0ZBC9FpxWSuUjrK+6b4nqlSfyTv/+O31BIbaAo9xu+gMaTWJbbB
guNeKenROxXr9Ug6ZerJfJGnK1Kuhunjo6C3ui37QdPyh42opwDGtZc1TpIV+0dE
dwi+3YAd5e0fUlMq1PS6Sw4Kc4PoPxu5dtZG1qJU44NHEWHzm7KYGW8qvdZJrVbH
FnZn8gTn1DUS7U/QYpeiJDSiXhABHg5/I7H2bMDREOsHcplTJz/5C9/pTaLUlWY6
Bha3VKiWku1ZQsb5ghMlp6S9Ebv98Sou/ST6agM4H5PbTJWqfAuNiwA73mr7BNUo
/hhRKwuMM4UXTEaZSIrn5g3CSaNhH4lH1mFuG/ldRDcGwlCMMvqsd98tNoTVpvEA
vOsTzuTRiuS6Unu2ld1GSEBwmJW7AH57EX2IGHy/Nsv04QxfkrBDld2e4zvUWplf
NUzK7rcuVkL3sv7VmpG2y4JUHmSfpu72++GJCbQ147NiPy7/zPQk91jbIkhDy89c
BEvE3hZQ+V6ldW5maAG7V2MQXDkOyOgQyJ6Tm4/92UIhVCvvFoBBJWz+t3K4Z7cg
B4rEsODBqnq84Df+FMvgXkP1mS3H2iBqEsMh4cVTOf1M3ze77iDByLDj3olwloUP
SGVF3508jVpSdI4jbYCE2vJAA4aBD2ERfeoGQx2bH2hwon2yuNBjukGqNgUuexcn
xas+lHDZSRY4YvGAANYxFo/TeiZ2Oh2yiDDRUCtnoCFzdGzrvh9JvLJ5kK3P3PRB
1WO09nnukH+H3x6US3GtPotsbyvBvk8EBBSIREe/k1su735s5nGgqOgzucuVTYHz
fFpmtXLeIdoCKHJ5wwvtgkhY91/tnlA0j65i9GDfWlOAdcOy6MQ0DwNAXpdwNbZ2
0B4LsN2eg0oWTozZ/X7EtrrLtGAYIIBmBqMEdsggRiKgVsUSS4C7RWmGifuZG1kX
HdmTtqe0uOiZpfM5j2a3fD/qYwo0lcqbN6VxmBVfZbpbceMOsVmE3xxIOxt++ilP
XMAIqVHDsfDxZZ+6KUXmIYzs/flqHvd1wI8txBDoac9c+DUA5tJj6OdWd58SReWL
t4MJH23vfH/PLzTTpndn7S4T2q5r0uRrokZEN6EcvUSi+/ihdVk0WvNTftcpJi4Q
uZQV2WjLb5J7dAxDXh4yldpnIusX38lTXFPYdRxFm6fsiFxUmOHBHDPOhWzx5khF
gsq7dJbqEb6u1v0CnQ4iTJy2tFHWfti+Z0OR3VZ5D8WtvyGlJ4jqwBUWRWeE0OvV
0V/8WakC/2oc3wql24U0yz4LDhdgtIIMMt1XT6ypYHTsFMQF2Vve1550pDNQYE42
OE5nfEwqUQH3cc7JZ/YWPzUJEy5MmbRZKBtE5f7Bu1g1pt2yyhSdDCeiClq+eaCv
Or07ltiM49UGF/xklkIQV60kR08SHDzlrTtSckKUpgj1lkteBQhjOKFbChU9vLPN
hxndOzNz7FOauuLJiT6dZPevkKoQNVd7WUS3A/aENNdS2tKnswDBiq2Wnf5S+1nl
dQk2kHkHiU6/cxzvk1Uw6l5UBP4FG4WPAFjsgKMf5G/CNkpJiBNcNYhPV+eJVkyz
B0HkFkf5o53SMwXOSD9mcxukCBKWDmKEPvh0A4jii8DhSbuzq0kWMqcoeWHfkkO+
FCKAkRnxvXlqLSxR30H/2lkX66bdUU2BdQNHMX00ytziJzEmGNmFgOxhq9JXpPI0
I1lPEd6KcVQNLTBKQv3ropexYTfJbVvx5y6BNRZ2Y3clBhgTHcM1rW2Ry0ljjA9u
YK6iKi60LEdm8tVMPR25/LRYDXbKMq0YPaK1bzOzE6rTH137ZuXbD3krbDuMaCqN
eGMCEnktU/cXVrDXr9hMrGdb/YyuqM6m0Zm7qwOtPWTHpe0Gh+qtm6vTJ+qu3Akx
k/WuFDFb6uUK+5kFKg7ryperHIDApo8VM8rkAMJ3s4kZFFNV/B4rzCvA8lxqMbHo
3500N23Sf+6PY7t+KHumtl2pqNvKo1WwItgTZuJ0oFQ7K5B4L+wUUN+iEtgq8GZr
yBGTl2aFbDwqMXePaWn7WXveNxW5/oNck+V0V/0i9f73NFSJ83kH5nxi00JlISI0
FqhvY9eloROGy8IiLFXGlUSAb4+/aOi0WzWCIRcJ7Yyqp9LkoQ0B4Pp4ELzUNGI6
H3jogW/b8+HkT8FfaNCV2BVMFG3ifxeNGVZ5SsXsJ6uqFUR9j08s+F2CjeXfRz4I
UDB5L3nxYpOiRXSGnIEBFLOBb1Vs+OyVrGgXoFCMoimW46abdCIGkEUJzkd4JQx1
a/HH3aC8/XhoZGrDpIoDbfUsRoa1JLLv9xA4dXUlngo9K1YqxKSGD3ApUoR04jLB
72YOFU0xJmE9RkJ1e5QjtHP261/zLXQHitcj+mlRMWYcxeGs/bpQvSaq0Zh/znW0
7Io0obR5u62zuifazpNzf17IPTyg5XrAGOO8yjAAhpyOzrrVS0xmsvBlyJMDYXXY
9aoxcPVFn4MGBbNVTjJmKsmXY48ovjSD8sOHtFi3sTtOMzqkhd3OU08OKc9lUYJB
Eo421aSbuWH5w/GdNoJU7Tq6Her9/zkzK4acZ6AHUVBWmRUc9x13dY3OMzBBiz8a
JpOhOI7Gwwc6eTYkb9h49gtJNQjy3uNi5Rd/dzF8/2TGf3a1wDiiAwnvH0cUfIMN
prE7yyGSqFZdkJdKJnxYnmgGmVmspUlM90StEyPlSb/R2udPA7xKV6A6W19KgUs+
5e49Fg3/0pPBYNYIE6VqPw5Kmwje9s33lxACYlgR+4tKZS4hFy9A5QqWCKoIIqlu
sCFevo8WwrK3rDqBcz3hQoCONs/QP1Ufa2ifzq+xGdStC5l3W3IVgDzxfgxC0eMO
QP4nvs8Eqf3HVU3DOAr1n5rlaPF0TfYhn5RiNMLY/YdVxqoDZhuaqdJTmcgqgtCI
8OF1wrOEeDZBN3+oeHqGFT3Quze7dc1cc/FtyKU9ehQDcmLvwXk2EeRP/Z9csgYT
mmQAORQwU89qeVwKCvO6njvdWv7SjA8pWvFfXfns4GyH9c5unFq0I7MCDzSS/kPv
prHi0IVeagLrrCD3u3lOGzbypt/K/7unajwcAEYnZQfNN8X+OVt5ccIuCeVIsEMn
91Eo5Wou+nyUEu7cdhkdwoFUe9jKlCcA3G8m2GOLRespKifURNaOUdwl6ljHGGzm
/4MH/s/MHRgmD4uUFuVKBQut08Q1rWSTVpePUUdo/zW/xLv+NCaHiX7+/7tdk5RP
x7F4wDkOdJnbUwVSxzH6bnPWbuGV6Il/yuImo/gALzdQ9KQEbm23FhTW3e5qJjX6
27apxfhY2zECF0+8/x8a5h1EJfzhcfbnk1cQSL6vp7PtCM3wx3NuNYqrswsQ1Ovv
MsVDe48zyKuLIx85BSZfd0pa/gJuoJuckdcKhK5XZaOr3ExxeclCIur1MMknUQgn
M4QrXDBqBjF9VSwCM2B2iPaJr5L3vQJHjRWRPlpUr/dlO1Iz9hgg/W+SKydKj4sb
Jp0jxv+rYF1M///42OikFlbig+xIDT3Dar9geesO5yBodYEqrDM7/eDYh2oR7J8c
gLcmCg7LAyB6Ud56gvxibXdTWh6vUO3Ns0vgYTV3w+pnWSBhCjV3dvK8iIdOvSjJ
ZpFe/uz0QfmAtGg71gRRQLgX1js+dkCKRMD15AQlCCtrSmh57OMKLcFuMMayHxjL
HQ8nLpbqRUzxZvG0ZE3+Ly12yDJOvC9fQ1RKQu9zj6Rn5Q+KUl8xs8CdA4AXNB4O
1qOvcBnXPei4Sp5HCXl06Q6T9ZZ3KvNsSzmxWDPGQkzWNLCtsLL9fvYvMYhecD3V
LS8yJpUOQ8fnLFo49KjPJnXKflXEdfX4qWP62KRCM2p/fkpcou1TlQxTPIbQ8CgK
olii2RqyaUU64ZQHBL0sYVLiiF2Xp3HTpUtt2/PxPT3jydZ1oSlLI6wkWVwNqA5b
YCjYE/Bz4IEflr6UPSp1ZHVbEieugnuchMCyIK4p6caEqOErcolJKU5NFlUCMzgq
EKtcVSV8H039YkI/zxqaoR44SMU7vSGTiqXeZ/o+oNWBbDVD0NmTdrIuafunJw+Z
tr3EYAEo4qjialhuSMQmZASX57rCehN3bcOfBCmJFJbpFulH56h4NIPSGktk7o6H
PHXtCVbGBpQei8tPavllfABnr7EhIpItYLpvcY9E5CHWoiPSX1EE/8ia5gEp1kOz
rg/q6/ZOYRiAMyu5CVgmenDQSZafMmcmhz1fVm8YWJOf01z1ETpeP+RS1AlFEm8x
wYpriKmLibjB4sXjzECULRg4Km9K9Vd8g9r9Nz2wPO+/Vc7uan4YoFqm4zbhUa8k
jPG5khRwA7DQaIDHQ4fYFSvXa1pIO7zraCOUDid7aJ1P1on5ANGY7ZcfWeAHdhKI
MQ4HEtxUVTR7yDrRGSt4iGDfTvKE9+6R3BeDuLgRUArTplAuNsfx+uCSRo23o+Dz
NMUsY4LKWFQz7dR7+vNG2eDkeONomYT92KMLF+VaRA6XrxhMJYeLrhussYpoLuhj
Bf+kJ921VVjhZ8SJYLT6NZ4hU7qUfSFLJCKh8o8h8xnhfkP4FoVnh1jgJ4ATTpJ1
Cw5cs+9q0FgqvJkpxCixL/tRKp8G+EARuUorohhtUwifyQ0jSOHGLA1pi9ZEyC48
ZjF86Gr2cvt5rrO2gavbw16+FmrQXjI3ZxAbdNAcXA0fy6bw5Te9el/7/CsPuzZK
inmHwiUJOXB6GKgUeK8okBoxZ2RZCm+5plDCan952mM24CvmD7H+vjG7Vq2HM/BZ
2RFFx3bN2bb0KFHiVlNirqKxEhgCcMVISdIF33+X/JePS0QG+8dWmg9m+7FXy6ym
WHrnLLacn1I8lJDYaMgqUMBa9NfLlX79Kw7pspOPKksAMNZYYCBNz9S5iQKV/dwc
cCAh6VnD7WOKx4P8iop07UKa8H3Mk2V3DIytCZP1T6L77Z431KC6nnyXxiTvPFJ6
xlkdF6NqvfviT4J4tbmQ07xwVER1f8CAWMQ8s2OxcMVbQwfIn82WFo9e6vNHZETh
YaLSLbb0upE1BFZlosg+A9nH87dEe816NKoT3S2JD/sTkeJ/JLkEMnkREEXdva+l
IjM2BJw1y8JnRoigvQYmrfcWHxUpaeUQgN4d8Bz+FVZxa7GsrWjnVuE1x6hKfYDF
PBgZ3hCV4YJGHVTG6xMP0qh9ENBEJZfCfLlZbYv2kizfeVPoNhkbpGh3I8EC7rCi
Hs4+ab2dPiFSaY0t79ZiAOOPbOqPnlPjMiJxyWGlbd3oLRwXIiGlJ24O1ZGAIczT
8PzN/pfRNj6yFJCDK0deJD4OSJS5F74vxEufuuwRX6fpEdwtb/cqNVbxllcapeIJ
s5K8yj4yhbx13xSrq3Gc72/hR9HhTiX8Hn/veYvONDLgtuIpP/W1Jq8JxSiBWl1o
VwqO/4QSc0jhrUl1gmkG6uBRfnpBiZS7GQCxpQg5SJQgl/2+QP1RZ2f8jLfqjtqj
tbxqbK4iZtFT8HUB8Uviyp+WdvR2W9d31pTUTdtQxSGpo9Lcp7iacO1Np5Ui6tlg
T2uUQvjEUOkehYSijleU8/3p0qoibEbhK82ntHrDNzsuh9M/qsrk26iS6B+33zzt
Fk1le9NZDA9NLSr+F/78l5VCjct3EzM6zeUCCbTx+ZvHiRITgaVEsJA1C/bB8X97
UlvzMcgSxpRHjFsx2xPAVjBLPMzOo+yGY1+IP66QbqDcDbGK99ANx0bD2am06Lph
dd12YU0QvIgiWk1f8F+xJud0NlIKGCgV+xaOFMHnVIwc66B1S0myfDA+HYX7S43f
oaj6fYURLd66zDB7Lf8FG7hYdK+RYi3mprCoUu2qxVuyuP4LMkVQLGBn7ClUdmTo
3k3o/IQWuK7VMJw/rupX03WqAC7MCkCJBRDQ5x/C67sftiijpbfLTROusdxfwAbA
c0v9/kbJM82CgwacRoYXAutPyOrBGZBgKsYcWO6yhqk=
`protect END_PROTECTED
