`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBLPmgb/Lk8p746wHtc+a3VBu49O2LdyIWu/0KGfSyZgZBeT0QL5S8Cxad1WgnvM
B3oUYAfVPmeSyg/ckqZDmPDJAwrMSF3xj+HZ1fXoSz9Ft9UP/U0i6AysE+PbYbn1
G0LoXC10e3mot5zyFBEFoKFK6K7H/1j1GnJw+kBn+8Er/ROZ9zBdk/U1c24h3XSO
`protect END_PROTECTED
