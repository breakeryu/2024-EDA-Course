`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/zI8lo7VbXMu+0qZHnYW9krQqTOPSeh0TwbTNnyFf0upKGMNfikIh7Q6i1y6g+WB
qTI9m1tzMt3cCwobrbjuArVCNdrzE+5hMGA44tnweTkrDMwG9RSBEKoA2vn3ycF/
h9mpSEznG/zsJxOonDaVMEXWed7AZW6Q068dqiisMd9bN6yTAOIotQ1b9vs0Riit
9hwbBu7phvvxyAb+BJyCVASqY7QX5wxyzgqWbqHzSuEyw0VHroXwkBYMH+sTwcnd
+8VQQ5DkH38+zFx2Lv45+C02GnqhOU7VoTDX1xJ8qmFhSgj6pQJeQeCMN0oLpbLr
gJZWai+gJKXAK3lAtEmeoPtGWxhWxQirbvN9KaU29+VjNbZGXYxvZRbXO++nJCoE
a/l9Oslh3h89gzojlaqTkCjUg8cMJ/6QWC/sTi7r8iwwmxWdz5/bFDKGU+ZUBZgB
gsGZZl55oXf7gQa4lVD+c7TbklRYHgnbmGou1P434pRMR+dpVh48J52IK4Staye4
xEscKvjA7Pxd9ff5iSRiMnMHtCCMmJs1yxoXlQBI3YDmimFBq4hE5OVZBDpHLzS4
EFuGY1gf4J3jEiNmBjwIBoHNrfFrS5Jhz78e316/R4VXFwKyv3265S136ajLQTpo
Osyc67TUrQdmQJLOdcdOlBBTeVR1pezsmQILZ503Dz0etnAEXhxaTLAcP4hEV2te
MYnJGDlUmBH4VeV8XYf2a7GoLx8ppS3AX5lww7Ym50UF1MVsw9PPf2GEAJ6EvqbP
MDhy0mXHzi4kmHv/BKHyCt8iIhOSzJGt7Xtf1uDDbKdAPVV2L6uveent2oIVox1j
avuQTilgm9evqVr93U0GVXOUhLYjZ75UGo+o4+CkAL5RsZq+5oRIpis/hep+yD9R
F+P9RIMl/9EBCpuzenuMwz22XajDfLRDJ9AqiGpQZ39B5nfAwE8LMrahslDCTAP2
j7Mm4mUqHi0Y/1eyX9c3MNRiZFF/yWsj9PLVdtnAPqaNSfWjMkEWsdVZVKd+EZqf
gDNXgNq1fwzTT6CvmbTDyIRitbclkwfjNkxyKLWoAnRL73heHiDwEV6CCsXOy1/d
q4FD0UJ0OHb0cy32TODBc2qITcNKBqVMtCHTU1O6K9Isoe6s/fEsEd/07omLA1SC
tYsg73uf+QDvapKAS9N6++jLUOejhp2DZ6O4kfm3+TTpmmPzyN/xKYXIqSfyz6Wu
x3qq7Oqbhb8epUF1DMLtb87wS+8EhMMq5kw2o5YTeWbAn2gWCsDbGnVk5ITHKOjI
1HAzLQve8K2uAyTFzAd8Cpn5J6WdDPybCf3SWGP7JYhsS6dKjnG9zmrEH8dzz/Kd
3X57xGUm86T63YXo3Ud+v4u3rFgdGnNd5dr9RIX68bULJtxwkgS5E+ZJrJHjIsz4
Y6ot7rVk6jLpudUo3FdpkzFCHpjBiKjhhYgvDru6+0pVK/v9+l70HKjVsFVhFk8f
fParZB6nhJ20zTaiauIs5PuyXnZqA74+8jRORh349kD4Kt7RhJbCzOchjfwieky7
gaWKgPG7AnDqGtZrQ8Hasj0CpKhPYBaLmTJRXDAnAYSLVFAXkgPNZTIE5khAYz+v
skawlRdlYvBXVrGxt3H2mjyfUL2LWsWLJcBV1lloJHq7YLYwkVoB0FmHlgHPyXcV
sNyZjASLFB3E/oCX+8n4Fl6avtYYw7DVDKXAEjCHLxxYVHMdHzyQClyJn0EW1NYk
Sq3CCnSdCnL0Qt8u8yWdAm9Nk/50acO90OdePVhvRcbNMRHdQ/Kq1t+3kauPg5CU
fdO2RWIYnNBegjA0SgsRHqoslxXKSsocVnYME5ulJC0AK6YPpGXuew2uNiv+nIgw
bFcZkQhAmhGneU2wM1t70dwKZUZbO4MS2aAQHHhHuXS+8Mb+jsGNQoqZesraKLKN
x5WPSSGKaDgo4zInUGboDB5j1+oK2uKq2myZ5AIZRCrAnedbkklNYnjDvvimy9+W
4DBatvXwgs3AfKkNak3Aa7QAIMVUPps8YnfTSJLL6sYUlf6GQ3MoPtp+2ASnBqNA
d1Rym77Kurs03pTEGYBxB4Dsqj4FXhCDojKtpwcXAheqrhcvMr9NXVSListdS4VQ
Q0lOYMgBAJH4SilG0XSnJHP5kIHYW6BE4gWlwavWO1gHCNmuUI0cLN4ZSj4K/aE5
ujeqxRC0yOJ/BURiHOhSJySJI0/esQ575R6yEoW2ELc3wIolBgO0JLJ1Sz6K8mrg
UmT1GXubDk2goRnXRWzebsJhZtbJufsbcXxPqqVF+95Jy3gr6+XjMWRAC1woJzDf
ICTk+WEmkJ4pIRGas3s53icfF/kqgJ8NaAE0Z9L6tsSZSVHZGFeM1adeONQKY/jm
eYyLpBNRfkqrkAUQQnYmicsvWL86sNEMCAdQnUNf6kmMUoMsViWsRpRGs7MQ9LhT
IlTUOwWYP7g4LSiEEZPF7kgSMAV8vZbRa/km7sT0HR84th0gECtLhVLS3wkNlBs0
w3YNvOJuP7fySM0eDB5TQXaG0uBVjMyfkz8TAEHFNKBnPUSgt9B/xgdHsfUm9B0U
EflS6ke3fh909hGY4Z/woP7hMbKXsRXJUy7M/JxVbR75DBgbNFWgk5thN5vp4rYd
7DfW7c/T3nTQduUg0pe1W40p73nphvp0iQ+bZKmdozt68TidmAlOhRl/RLlouCef
CXBCEKUEK3LVEXkw4ZhENUyCNShb2eS+QfrOKz1q3jkvweiIkx3PFd17mpRjhL2S
qDajiC36kCBVI9xBvtNKTWvyYgZeyEeEShLBwzlMEGPlItXrelOdMATHCVOwnceJ
/PgZ2I0f1uaMNpNmQTrl7ONqAnhf7Mt0ceHufaMZBFTLO4olWYdX7FmDQj0GfHRX
SChmSrfuCCvqYYWBqeXX4KN7wBFy7IrEIeoF9Lkpkv7RoVM/n5jdF32R3KxMRFJJ
fJLhfh6tJvDyOEDoyl8rl6xRWtCrxNOsw/anmQRAM97OhlVbXjltp8mOTgImhRTj
adI5qvG1N0/MC6L0riRH46u+2q2BZnGhCpbbq9x8er8CsK2PrXggFJDmcQNMjk9w
pHbshJ/xQVr2F3uhBX7zik4uLqCdkldzicX7SV6aKwCE1Qd1z8u4hdSVQJYHekld
US/1ywungqMxSK8tZRrUmRdby+XGLPAkXUwqeuLH7ZII1YAQ7bQE1IxAM9aYEwpZ
xaYgGNTIDywVlXXE5aayWwCca/flbRxnnuwJ/tbRiVeMBg/2hMfI6Crvdrqwul/6
JkMt/F2QkbeYjQI3ivWc77Cax3qmJky3l+GnDllwyN5xBsQHf1CrPFsBmX1r0sqb
WPdQ/PfauolmX8ae2MdvXkmlp7Ja7vpHXPgm91m0I9uoT77LKinAV9GVyN9WfOYB
dXIg9/xpC4yS+Rni3wiXBYn0s9cpn0A/77OpWGKSdYpFBX1l4q9Dlh3LAieIjVnE
QmmiDE9mmxVjBL5JqOsx1TWlwd0hQMRpp8NnRnl6OfkaiNIs7rXZc0aYgjNH0u9I
yo0YBvRMQl0HUJq+CHzPD8lMzVOWPaJf1Waa4fH+IsEjh0CX60DivoXv/BDCCjxe
unxTzo8rs+ZUkrw33/bH4qSc9t4q/gJhGYgYmOPsuPwfVhY+a131/36rhbsXpWek
5QDeHlik1p7HSaAadQOxBVWUnA2hmgcpNuv95XYoBRi/ZVCkPqul8FikrBLFCTid
l9YTX1TzgFI7/UtJUNCFx3vWtgvKJEXaJtyEAdAUjKl5vRHEgicX4h7JEyXDVcW9
pMgTiEgVfcxnzdTHoWH9AiFAShavIDYufglbOl7urZuC3UhNXKdsPhpl5AN9wn+s
5O3/RY5ol1ZT1YXiOKy1PG+CzybTiKEeHZIU6CE/4448hiqslKdqMHFvlGhmgVlO
mPKJNNPpC6D3yrm8L5uuBsGFANgHbR23GhuQkj/3FjG37ePYAcKJLd6O84/HvZrY
69G0LgXWnLieyM+Zlf3AH3HHBDI5W1RAhrb1l6TTJySqYN31oNbcB8yxWBoUYjDr
N3IMj3gtn/GV27wt/WEUxmX4OCkK0/QT4b8e/xiapo7AsPvq+S1PaluK54ECgmC7
XlId9aFp4hrvxA73q2cgZEhx2bwxvHZ4uUW2wcpP3Ij32jnfiC3lxT4ExOl29Fwz
U+yDnXqeR5aJ/OAHyqoikYDPKq2tKRq9ZaAsHOTDnU7hH5Flyoj6IrBUvsGyNqOy
I1rat+GjvIB8HQjvk/+X6B9+Ni9yVWZYx9IxJ9F86xMP/xtslhzbwG9TaV6tDL+N
Xr3rPeEbp4mvYAdar1dDYfAZv6SNehnyZWTSHSG9RDUf5m6dlpxiaUUMo2nFcvKR
beZQU4HZ9urt+Q5LKNtVcFKpmN6QNhhscMsg2HJqL1VeeYXNoN2zQimXsJyW/9py
660bcxdjwLzD3U2rg6HEGYL/BQ3IZSYvh/tyOKVMDdlbdKAeBvwFXxSXvnWUjQsr
ZTATFva+iCAybqmMDEo3UHCE1iDJFO2mfeXyd8kuw4Y6yq6yMFLa6hklvkFY1O9O
nSj1c0dQYqFoq8+TPr3EjQKSRavkk/C1qcZKM3vXnHXjJ5kgr9DwslJi6QcsfVbL
2BB32DqKiB8Nu7egSVPhAQzXN9GR4gwLQU0O5rANEfK26Z62gk8WzAfTP0MQsP/2
0AtA1AqcrW+l2HBJWcyS2ZFlOVDs/V86ZRwdrJmEVYA4siSpRP1ORfhA9IfqzVMD
l/J3g8Rp7ki5L8UDXARrEO7YejJixXYeLbm9VIAzErAKkwBChLxozynJp6YxKYOj
i0PU3/9a3oL57sqA/Soxr21giaLD6v1pTfqARsuk1Mhl2DsBXJTc1ymPSorCKQud
8C3Ado0jGSa2DrRd6bBTsn5nppY/sPJxP6u5d3Q4nhYZ4wZala3Ai5M7QvVdvji7
0O3LM3b8z8kNf+eWdkVVMRW3GwGfhYmEcNGHRbNRxUWUnwjlySnz0oXCQ2n+tL6P
eQ3wtFjkcmcQP+mDZt8vTi5rf092vkREPybB2Ix7WPkuwroFiORIJ0wU9AFkCsGE
P4U9oEbILrNWGakiiLM5UZ3S6SWI/MCrGDT0zM+O8NRQNABioCzqneuw5Gw5gpbz
ikBTnZCWez5Oze9I5khh5SCzCnuktj/VROGOF1ih2K1UvpC40/x+0GvYMlKrbOPn
GXYhj945494ceP4xd+P+jeAk9I5dQLta9yECWPc7Ksj6gWaXiZb8bHzBcxohJXTQ
jcG8/KHZRocatQwufOf0OjQiNRjwwQVcd3muRZS00YloNikI2UL9hjS2tpARcIlN
jHB30vNPvJEFg6vHqQHoZRKm/1N+qrjoRissVTncNc+AFndA33Dv2F/HsVxu9JtF
fZf2Oe1YpnsAnf4ut+EIhS+DADf2/9oxJFEUlq1wOMz3Vhqcw/P/DAjnvo2ltqSF
tFx5hiB0rh4H5lODyyhM3NClSq7SlHZVCdzo2ZYu8pndqApY+qEM+15d7D/KpfhP
rSsj2weV3M1QeO4VH1Ps6f12WNSfe6UaCirBYwMVZPJ2LFNACkJXXbt60l8C/5wY
koCLhWxHkOCynNXn7HA6t/59Xi4NttyhQchbZxLOUAil/ODaw/xGluB8peVbG/4Q
XB7JAg93E+WkSJYJEUxuQtgYOlhHnCS0/JmjjJ4HCbyu1chiO/Q9XjjEHfuIimXK
TP4WlZHVwKrdcPXxq7Q+qSEkcUydCNSfdCnZ5YJc9X3q3yeliIen22jKFLil1b47
YUxuRyNcXSGPnbJmzG2KcsyocN0jjTWqE9RGpLurireMR2+QanqjO99neen53Twg
toNMqG8p6BV7yU0lPtU0HZCS2hF/2oCYUO9fQoDS30QEuT4WS3L/eu11N43nUUjb
eK2mDl+GLuBSiMJMcuxznpnxRxPLCLiKV28O3Eox8M9E8ew82g/cQHZtZi2XzCwh
2Gm4lY7V7HJpyxCaItDYfv1Bbhue5Zsgm2rdmadjBVUb/u4Jy25YTvDt0l+Qasw9
VTOvILLnsQ7RIWvdJmkiiATZq8Woj9lbpG6dw6+LAJZx9+Miuw3BGlk6EIdRkZ5/
daUIaopwTVY+j0Qn6skyfmXZSG1bkZIGQrblWGHsOfcQ/PtzYbO4+jUAmfXRDQMy
lIBC8xI9Llnggd9U74WF2pwHiG8D19XXY+6c9ZL/jCMuGyoA8wp8T4sF6ONdNte9
Or+v2zSzkj1ckGJrTcwcR5iJf+cEA9np6R6eSSrcf/nqudPGq9VuqkQkNgexOGdn
3/bcdBNQM8KmdeU+LnbOXFZAcncY496ZV6MuASU3N4d9NyN+htH3Cd7tlLDjAkIE
7rSjaApvPTEc4UjEkx7/JF63wBLAEh8672lFlUiHsnP1JLRS2yknE8mnDi4GFT3o
+yBVXecTCdNIiERSQN0Nq8t5/+lvhJoJO3bUgTBdMGbltHJZxX6BGofrputkKc6B
3WWPSdinTlHF7Sb+a3n4VNw144qVeiOUoNJM1qBD53OEac/vPFw3VpJtBU2ItVIW
foEgvzIfI8pxjFAnGQMsTtsx164Lzq0KVsdegMZnNGfvmcLxqMhZXzzed/NaaMlx
kYkM93YBxfWzpf1tpq8Ibj/kbGBvgKX2a493zz5MUBeYvUrvoIcA87iXQexFpuUd
ESfhQq0C7GIDHYuFbF0zBjXskjVkQdd3C8dzr5Aq2CFXdoqnkk2sUr0ftz10fSuJ
oT3Izxun/+H2Khq1J9Ocv04vliJXDe/ePZCwa9rxdlSMmcL6+SjidA/0XXSijCFN
hoPlXKs+tDvCUFfTBCllfTLnA58QBd2wUiqSGaUOR8NDfmZ9PtXyb1FfiKO4mJXN
T0fjXvFO1+oNQb8vHeDAW1/nOOoBKBnoFbG6eGt6AMPJvHvqfMwd8D0TYPocfeju
Q0a4PmADCx0eRPo0uRdxUBu6bkv0MsBg3UWe4qoJN1lCy1wuN0yhWJ30b25Q2mmX
oZ41T3lIKCj+nwwmMiArWVFTbuY6UjZlw7owUTMqEPcb6xMxKULSha3HVtJTofpg
7T9DuHmuza639UdrGWPG6r8zfuqGT3dVge/aHY5vuSFIe0tURFebot9ibKCQIQng
UmpA5y0QRIzVyK77cM0GI+y4BNz2cGZKOhR8zL/2opHx8WV47fUjmoDZ+wxOgvdz
V5IfIEcgbimMG+XtWkM6KZver5ZII5nqjYr7suqoScUeHEpB7JhvkAbFg2sd7T93
J1uWnO3Brups9EX4GRywuD+rVPe8Rr3icXiYxGKatOgEUBKj4vkMpoP4rNtKZXne
PHiB3h8MbONGMh0q6DzbmqExQ4lLT1KX61jA5JbD5tt21WUuelN6w0B5+4KgRBUU
KoPIBoQmtEpiMDUf2SCbGx6FesF2gdgsjjheZ+2fl3lMV4CO8zhkuYn2xVXGLjxn
QRxr1edhGLFg54PHzKN0cTWYgbcSBKyy3Ih+ofSy/nqcK6kvcW7PgWXJlJ/LdvEL
8DmSZd8ejbLBiFxA2LbLpf0Rr6mWzRJ5Vh9eiTWJ5PXcU0Skps0Qu9qbqb639lfa
+iipIwmUbmysP2xtuz4o3JlHqEGboJ5gakm19OmnXZkxjpPF6okHMONND3yzaOo5
ev/v8LVGGZUakMqd1XQHGZpPIqeKBjvFKnVHqgI0IUyUtJa+3xPcofACIXhpdrr1
H+ajjPYrP1+eAfpZhA5HHoO0yAXFZJH0rcEbYfCXKDxvYo9GIja/r1o6vkduIxyQ
Sd5NfGMr9OQ6siWzFXRyMY5ZyoR5MqWD6sJRMYYn95FZDI4YXgTQG4GvzBPkhLFr
iddwRcRRzbRBzuQX/D6MZvyjm0TPRkFeNDTuMmm+PHIPOM3zhbfHM05epSUpt7Uo
lPg12Tf02dd+qOvcnxEKsA18EjCcPXStulyieExhAe+JqpeJulqCBU+skX+/2rav
9ev6Ux3mlba0TfkvqkFx3NvVDH4hjKQlynkJnt2M9k7IJ3A1CRE0O0lRtBBewYyi
WcLbhmXNLgT/dl/Av0DaiIGAyBKP36WE0aWc+jUDD4nUPfvjoUTHZV84hUip9CtQ
6iEgD83NXYwF2O4/vL6i3Gs/voS/REMyyzJQ8gDrAB/0E9YBBDvWRdAxXMAUlnP9
YgSkoY+9670rFvevBB64den1DrSEYWQVsRogqFmZAG5viLirjYewWd5uT/oDCM+I
/MKsNnYr1IU+ynmWsvScTdR7pRcXUN4sdGm0J1RyVb00+9zCG/QLjfIcMcsceDxv
xPY/e5ixWorRItbKuvuZhZlvfA5T+kX4exT3a1nXp/BKEbROFFL/UDZj/BHhksX9
7bPAo3fKW4gcTjpecB3gGWlgIhD7fegk0bCFPrZld2hHOY71RrF50Yw9BPqvOXQP
6Qz7wM74YRxBUou7i3dqCmHv+piJ9j9HhYtkSmnH1D+2N05qazgx0qHbDxfzwUZY
aJb4FDIdGe3XQL5UPzxVW1K/aMrEU9o5ZB6Xveu8xVfti1XL7ZpACldj/lUcTwJi
TJuNswjyVVahQ5S9QEwsq6Brq3FbeK7+hvqaFnOgBtkzlOqqzxiKbfZwllNvtE2w
8klQdOO2dfzxN1dmQV8wXKENKt9EmJ/oTvVhwuZnzJu9eFlMkl0g1enYSx1Yg701
FQhJexVmxCzubJXSrZT7CXogUxhwWLVbv+XdEzymZ4c2OJalWvO4enJUFbcrJSob
UrSAOQ1moWHAgF1EJTLxOgLWSNu8oVyGcAvtwPCb6qQo5XwZSpRgDL5cFCbKvZc1
We2If5QkOJ5wIcP8gttoLis1r/yB4R115aURo0pThagNogDjcyySnC1TL+9kEqRt
lCnOoP4bR52jWVC7Kyz9mrYw+ATNNDfX8QtCz+mOvrDWsxw0RQ6+1X5/Ogz+Lgey
XTXQqYJpR2dZRql3ckYmUO8crN9zuhWEGDo0aQmYZEo9VuIsv2WzZD2/03zQVYA4
ffpMT1cSt6ZvKHv1ycFoqedQgedIpoqDU5I5HJo7w1SPtUIBcv9YsX7ugmAvFqVa
KKwxnF8cW5sk6q+6sulKlxcsh6MMJeZaTeWvE+4pahx6K2Bccw+vNFgekXEfyCJu
SAHvb6Vdik/9jPPUHTJWbSrlw9y7LsOVTUAOyN0D6cwPr04cAAOwnYwCA+n13zKw
hIQvkAt3/vtTuW1v91Rk3ukjph/oJYBIt6g1cWwCWUPX0DVjFnX3q49kLtc+xkeP
eyfjvwRy8mSAiSNLxMnNKD0b08SbHZbngTz23uDFxtP4peZWWu6BgZQQXN1Pf/XE
LcbrDGa9T9KFKD0EhdNb8pH5cSiu4BnaASAntEVYN0qTc/hPJT1BFtO4i/ol/cXs
g+z9XGfrP3A0bi8mgGX88d8WX8ehjIBfcjdolGEBOKEsdVtDW4sqV2Dh43TD2V7O
MjY1HJB3yoI8MjgojK64v0bdRKrSEoDu6xLMVbHXPqqduwRByy7pynYrAYlLKVCj
cuDxqUJ2uD0BW13ChFOMM4IUGSh+QPHckLJsPoCh4HT5JafRuqZp7wkMG6HVh24L
qrOTg+kwy8+Ew+tLFd9pVL75ikXSpuw2yYk8WDokmykRkzAH2UoAGklrAIImxZNi
UI6PlGn889qc2Z5RYk3SPl8HzuhMV4bHcQryjc/3Ujn1i9+OQ7EswSCENZkHJjQD
jvrgm81LRI7Pb2Y3x4Yo3ZAUvWJ2l4CMmnmPsEX7NCVakyokv4UJM8FCREGnoTUV
ubVWjl/Gz+kxn+A1AfKlcfkqTmaQcJEDsyNC/QAfCXUWuoqFHLsqxTufdZyj1dtQ
665JcU3vDwta0yKqQEfOeWwp5ucx1usWe7s15gQXfp4NUiilRxxbBBG8Ue8Y3vJG
cfIfpUvyu/mdI1GinEAg4RgkGgbicfMUwIill5EQdHraP7kODScmTjKMtiRHaQXN
UrKeWz+FIRyb/qpiV9YtWGd0Fnj9Xjb/0dI42kPdN4rDUHbKQWKH2nploCOPb7Iw
mr8Gh4jhoFu0nTAkYiao01Wfjh7/KxW3BpYHj2P4R2AFQTfyyeSxt8w5v+Pgx0yf
vO6+qeOXidqZQ7fxeQ4stUo3ahrOIioocol2atTyn1q5wC87UJ5O20B7rBIy9b8c
0fjnEgScdmuomKIJiauC2V5XfO+GKQ9zkkmWy5d09ANLNtifpOP6jMGXDl55Gkwa
zSIjrFHebkuzWwTRHfulb9V0/wuWOpcT1nB5rojkk2lBvZOf1RVuuFIeX9HYUJ1h
vOPxiphgfV+Hm3uNRVtgj2gRAMnHqjFsZAWj0e1Kr2meASNm7wyqTX3j5IPz2vLN
f2O5nS72l+kCxFbzAbx2ne7SPjPv3zNtzEYwXSmdTm5fO1M8yyw2swL/4aSBL+La
kFk+E8rrJclNJ9U/Y/lR19++uWEDugAUPOraWY9288UVhjJJKSOTXnuoMCsDGx4T
orxT5IH9eY0l6lmeRczwsrOgNyN+Yq9cAAB4KY56azA+khtCtQlDFN1ZziVhUX1S
MawF+G39VYk8ms14jh4PKz+aLl+c+fU78k2Sny3acrFqydIlAo+9iHFvMH0iA6BN
XV3d+11Xt9bTpULYw7e/hue3QWtv2nYfSKyP7kX15MW5h9AvvD8egEqZG2uAz5Hn
i4XQfPhJeMxKYCuCAUkTd+TDRdlWfI/ydie0e/J7SgK9z/cg0K8J7p1NKf4cxf3N
9+mi+D8v8rtZ5ivglj20sjQtFFhQ3xe2AG7RMDS3oMNzdvigf/1i9DCq8ouK/wd6
oMluPnTXbz6M5wyk/+59UEgLdfdbgiHrwur1fhcio65h6DJCTwHWMobuHqr0kQvC
x7gfgn5JmF0VKjmeGsdRwkRI0h8gKZh5ev2zolTeYwL9LM7MIXfM2hKYwLNtK177
jjSvO07dbgX+GVXYV4aLLputsvMaE0h9nN1PjAz60XdlLtskT+ZT5UK6AgVcMh/O
ArHHUDQ5V1aHV5tARr9HuPEwtb6/8hwPS1BHUkWxYHPrIehY+4QfEBqZx1nY/kmy
gGud2HEEj8+cWYH3SFiL5Q5RPV0tZO4KBDs0WhRoC4DZhS7AHiRFomqKoEy9DqwE
pksXCTB8gXzpuZsyuWxQIacgWxqPRVfBHYXvcouPRSn0L2MsAQjOcI0hqEw2revs
EYu1ArWXsjRPJmYuNTTxyZmvLDRsMxoqzZNblVcz77lkOmjY/49NxPy2GDr5R+Wd
+OJAaifvOeWsVm6zXrYRmoyxTjlL/h4bGY+9maFeSOhcjiQsVOoAtwT9/lnHoQta
eTw5UTckSHoAKNH/uEOw/Gmozz0HCpuHlie5Jbf/w/mhnc56ZdAU6KsCZ3DnOpQf
6SW2oxmanKt3++Ci+JkX81AnTMXVOS2wTGodsBYGjD32YKt5IPzkhoR2M/nhCEN2
nzweY5F5k224qPZOtWAJ3jkkp+O9aAlwaVKrqtkB99dvcjvtYhT+wweBXLBc1AGm
lCmzpyVxgpxFCR7avinyJi4rrdKDoXUkj4vkQ9DaccOZ/VSG3+PLruFiFvtDfYeP
Vz3FUhjONoBSGYJKRuW/3P8rTkWJVC56cxhHKI/Mhg/gnfsC6TbtMsUZNRkwQmH9
ecr1wDMMUaiibe6ihKaYkFoHYOKeUDQmZVYFnQElG/hOIUGu5veUJKVzWQaosC/p
sbYLKp6wqu+qOmU4qiJHXQZ1UkY1n87gIGUfu3PkSO83FIc555xJT7UybTEa8hEi
5pAwWNfPrYZpF3TdE3NtbxzDNJrNpw163s/L+TlMmTLtupfNxKQl2Xg6/ny0UtlM
/igkJfGKfVoI4QlVErWjgKooEDOpP2SRelSQDJki+MlDQqE7/F2CN+9qGPXibhBY
xS4+leYAQk+kt7MyjfXS/c/5uYx2Si3lsQOMHFqFYA8hHD2+b0xtpKbZUDgC4d/q
5ZavsZvf56MbMhMF982PMDpC+BEFRwfQHbB/iEPtJfExXR/N6c2s/nSHCdMzma00
NM78E9rfzoy/nVVZHLsS1vKJTrR1I4dpEfzt++QNmPFFmYzUjGQ0aqY/MKwFaYu2
wPULJRHJLEVG5rA8NDCONgvtJPTIuvPTEEsuTU5WGT4Sx4TLimAucZDJ1YJ9xxzF
0KNfjxQDcgDtKoJR7KEGeDAz3gwsFu6vbJOBFpr0swialA8awqjbx6DzX7q5keUD
W1t+1rkpwYKiD2dZxdru+sjiNdXQzLanKP+WqoTOOPpsq4Ep6fNtY5RZpO8wGU0O
eND/Ff6clz7Y+R/Y+/ko+7W8PBPeH+7GTgOb6voOyKliPHP3gym4Zpq68rfHw2sp
ECAPUW3lAS4gF42Hl+LptXDbmKbvQ8sATX6JWqm6emqyJIC172YvPFkJ4n+nHuMd
+Ipey6h9q+dscsjL/7Fyauk9Z3Z8HKKUwa4qHatdiODmMLuiwTWpnybXkOPI7Pzj
MSPvJDwyaDqu//o168xGVUI9AVID4tP7WowUeOOw5a24dxx3KqvHhLvSq+k4RTEP
CsMAJ5TvpMNyRlNSdIQWlqb9U2is/FCx4m2p01gUKMxNH/zyLp0xmir/skGjm7/k
S1WHFjNch3F66ufdVLzqgvi2GFLZz9z71R06CrnBeo/NYs4je9CU2u+cuBIQJwQz
Lqd2ew2ytjSNkLeAbcm/JmPeYDXWLWJS3f6gDUi/fBlGjJ+i7CZQD/XwUSY8nR22
zihUXzZsbcU1yv12CdpQ3GJ9+f4n1oGl7YqIoOXElkqJoP0IUt/QFSkiRVKKb1rr
E38ObFtvrzwg+YjSykT9VHGGeszVfqeo43N5laZVoqZrWdgUlPniNPFFfKq+nIig
auHG6zrnOXkDjRh53Y90+D66yiOBH1PcpjtgB0YNTKa0rBvlL7pmhAQSMwBLnPuH
Q0fRvtSRcqGbi4zVlzkTmpuZq3KbQBwA5TgkAXYRJbye1u9kzx2Bc26kITi+abfY
96ZBJZxMqkeYxT2gpdM9It7fmlDwCZU5RfGBSjiw4lf1sgJryGsaE29yzehMsdQ9
xuo1fo3W3BUX0Yb/245G95A8aiNY8JbxsDdZ/lsQ6W6DODAfDpdeEnGN+XCrkoDb
vKpRpAMGS0+qJm+ek8XTGdcs2ulJF/6dDiBHxJ4GuKPVl51x3Ce+2R/4YClWooH/
4n0C+KiFxYcNc/4F1kYUpiPfE4fni4Jv6iObUNy2v+2wT5aAy/om06Pv7B2Iddsq
qGlO9oIzoGilsWmqYISTi2+wTGkE8LuB2ZlEltmXj23NoPjSpr5RDheFs5Vs9mXY
`protect END_PROTECTED
