`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ssxwSQp76NrK7SSo33G2bV9qABc1sptTzIzV0VvYKpNEPTo/jtvmDxY4wcolquRm
N/lLb0ElYG9fkpkzgStTazIOdiD9EHwxMelkM/xsecJUJRroe6dvZWF/2iVCiH8J
975Sktt4CcASCPjVqiNo5IoY5TeOkxoYs4rnleI9wvAsDw/uuszg8o7TXEQyrZxN
GfcbsYN+EnNMF0jczDjlP/t1krBQTbIi41j9Nsb05DQaqNlJ70d47f/Hu6oU8dRI
mEEDp21wEEI9zmchYysDI/r9pyU3oNOMnbodtsEzFK3v9XqqxQJiszy135/xExWY
VUVdoQk/p4zEyjUEcmRF6lI0YA0U82oCtsQYipP57zjqJA5hYpAqRTICZ2aAtBeo
YCAcbUj2VW3Qbw2bp+n5nmRDof5KcOvVUVHAxi0kumVCQJBMQWNOa4T7sft3p/tx
ddjx2vhqOoy9USi6urw2gM8w/cRs0QRtaYXsGBS+qGxPX1ziOlgvVxppEUCsWVl4
JaUpcMichi7NNqs5bCY3oh5BTENCKizpZnPvMohxZRr6pDx9m20Py0mCLzbjxbXs
jC8Dzk7GWhn5DW7oMw9tqSmprSAzJDY+A7cMAG+zhVSLfS5RGaFDjKIaQPD+mYoS
vDMLK/iHuN2xgJQq13kbz4XEMqAUnTsAvSyKNsFQ9SdHW6NJAYqYBBIBwrXNobuI
vPSdLOelkafYt5ho7LhKm4mUHS6/MkNfRdGDqR4y+OU2WyJ+47Z1VMIzGYc1ADlo
o2hxliGVDUG8h4Vd6I3bfP0/nSZUUTDFIcSHiG0TOq/fu0lRFJF8bj7TirNluTuL
zKgsNag3GET06V/cNS+BU+gnYmy2/3M5Nvp9Y3VnIBvy1fNdzPcP0dAmmAXHzMlO
dIVfIbC0y1vg1AV0+Gl3NtsPSmN2q9EXKE8LqzQEkT86MgVUP9TspMvkJeqP+VJg
lT7VXcR8aJKVGesiJEWdbGSO8KhowuSRG/di1BAU7b6k4wfSpugkLBeBWMGU9SQB
QF4dIarAZvv5OoXP7ocrut6UYTk4w66GacnQxA777jFEkxEtRIUbzVC0nNFVBgiP
zOLkSdy9nruKLVWgDLd8lcVPufIKecO3lDdNblj42KYvGe5mbkmAyqZMyI0WPMn3
24HvUBe4ZWVtaCobVa+ykkKPL5/6/z4ccjYHeUT4LvnDY87oI+kIxrbZgC2O6JCR
3rseBhkmPKW6lLsA0N4P96twPrOr9t6mwy0r9lJ0KggZc0SO3b7OdBji7C8seNEF
wd+oXgsA9ly46aF1ZLArcG7Pq6gVDxrnS76O8C1w2JCSWV/N3Jif6tJd++OB3A2w
eKsS38qA/UzEn9LvE9xpPHaePUBdkKRBNZ/3a4SZqMwJ8gNgf4+GmHVxY3QRD1Jf
Q46MjZe13fIen+c8ysULcYGhJl+FUhQUH1Nek7RqGMZ66bdfkBxv+ryw+zat+DiE
nw2GkxfN/nG4cdGyCYEpZvLimUq8pxbpV3AwkONIBzbH5ZeBjr2Jd6VbuiIm9/Ld
ty71NCPbRjDo1wd3wZCx12zZ43GFdKwdL++uRFM710Cq5dLYEccTdHINedEbpbUo
7U+ar9S8QlJh6sB4emyE7QaWSOS5KWn76EDWIVaOmwFGlBTrwnO/sn1Uvmniw8VY
/MNwiQM8IQ3Q4uOen0UAgqkdPiWNQWPvavF4vniMhuzvD4PufIIWSu09BwbknqxX
roIu/hJQsw40c2cDGpmcQsAyh/gKfsDH0sggyAltk+tFyDDa8NaAyJtBO2lvt9Ou
0B8LarHgFdCkEvkHGap5W4TkEQ6IixPPmHIuwlFXGRISxidU5MJJAeZO8PG4O5UD
kMpXRz3s+q+Cszy8HhiXqekb37+mHrQ8rVCNgLQcBrRZjbjhGUTnnzc37MyW70i0
Gwf1rOxOsk+M/nYiGvK9FWm6HtT0fK2YeL7d83WkVHG5QOXEJdU/f8Atf4F/dPqO
hN4JBTmSV+84uN3dsnc1E7D34djAZ7AB0BKiJZ5ocJMvmPgpghNQbTOfKH5Zmwpd
MC4XhJ3OsGD+i/F2a/cPOtwm3HRe/t1lpygFciEUAp1hBsSwUfapMTJGi7bAgzx+
RY626EXNTMtU+2n39IyMlvPgpafTPHsO47awVs5XDhzI7Fdgit22NWT0lA3x3b6H
cSVXft0FmlWxDcOUyCYymMLrd5QTzaGPlsvwEscgZTDcsm5PXDnGOHV7RuXIPIgG
he3vCZnJFrWB6SEwanHf+KPHGrBl8s7UfZUn9uRxpsnzQGZ8ToSDmBnL/vABQYSG
mioVqQfhMnMRTeB5VE+sfq6UyXB4ps1XfdwLed7bl0FxJG6JqqOSRNAe29VYt0ZI
Ero6Won8Qmkl4yaQD3w7srtiZzk8PQH+TvmQhdaD0VUk8qbj5NcHch9oBEgtIxGZ
JffNisItYnOMvZSNrlkT4opqZZWiFO40vxyM5wYoPImb1Xb13NMV6MmQYy9Qn0qM
Qlwc4UnWzJ2hEKBlW86yC2IrFp+2kOoWIpHnYXXyY+FRsy7Vowtm+j/X2faygMj9
6La03f/WWuO+3et3RKvRTpGn3HHB+/eWipoEv6xGpKlAfa4WVPe2wAMb9JOlnY2w
9Fl8GoWNscx9oxoG/nkuYZSRfOuFl2Q9vRT6V5VZBFkSMEnZhQGnXvNTX13zR0h7
X/Gsylcv1JrFiPURPd/ZCxGhpN56UGFWj0aTX0b02Zl4N9svqVSx/2NJAwIeTO9E
h+7zodpzScsLdeHxVJmuZKv2AcE6sDJ2oxsMfHwqqp5gpX5yEts4/3RTYldFgOhL
lgbxQw0dP/ZIaYA+Jwb1HZ0MTXnpwrEVFjDpmmYTAixWL9srmu9sZZhH6Iefnh1/
bEss+vEE4tAcUFv75viY2Jv8p+GTrUssMyqTJaHt9T704ngvB3hMEXO16IUh79ag
ZFyOhv+VS6i+OrO/4OSmHV4FmeDFi6Lukffly0+IHjrz5K4VZQXII7aeb1LsLy0q
uOJl9FaaCZlfQqGOh4LXazBqb5ojiTLUUhgplQTeTm4I80Xt2RnAhbcWDk1w3L0k
P5PcJV1w0NeHXA3PF4fwvL5Q/zZbOXhqOAf98A93hu+mMkd7eOufzcSH81cHZh7N
6B5JBqIRRaFn3LWkHQY/WxKvLJrV7lswKmTjO/y2diUdITCr+ejkryflQjG15xxV
+Zvl1pxkzsv7WurnQzzhEb7bRmaCaK5JH1Tqccryb6DicA8KWm0/TO9AHa0LJNm7
AFky7X5xQoprXvAACeRlPqvPnnDg3inYJ1tG9DwY/MbxK+PaTu/C2pBSbSMc0VXZ
BVEeJkSAqw1G6ksaoYUs+o96zzqZeQeEii/pPqiu3cuZ8dhT/SCuMDW4vPIpnfNk
2bJy94RYlKMJp1xfvuGcxbCljXl80YTcg7qvkpaSU8ZDJu3Ri5Y5MdrmmWGfO927
mCjDeid6lcQnZEiGm66T6xbdHom7bNEnyHETD14Om40tYWWJX75QCI0vi/V1FXuY
SoT6twr8k8XovZkO7oPnq+xRNa9pckO8t/VJnXrPz/n2bUETt1g54mpTAgbdJdmP
O/HdXsk+hrlgPYiDx2Qp65wkAGzICbQqE5wv3wYh0GdBUQfb7TcaquVkYe/iayfB
0Y0gCEZzmna2dfXBI0WNvtCwSK2+ZIQ0dOMPYXLDB/FvSLndzTOjlklyo1W5ib0Z
IH8tsRJrghMIiw/iLVkj+bKHVu9u5S+CWIDuf0hVKYUDZOboieQzsDpHW6TNHuBO
Z0TTexNhjyIrRgJd2FEjJnzXy8kLyEa4674ZbcC3nBreSMe7/hMB04Q+FAlIqJKf
ycW516A+LkVzwrNKCdtVVr5xD76Yig7OWL5qJztB1j7V3Ng2EnQCLTtVsqoBRN9I
eSKZfOwF/qpe2PLzlG0K1sN/kmlp9TOdzNFgGG3GvzoDXe6C73DkpZIgcVNM3bYV
xvOgf7lKs2PPPnLhPhCh3h4f4sEyl0J7xL1hP0ke5KwQpshHRiK3aS3K589F/PQc
2pRY3pRTsDTsQwH3StTcsFXoFk3pJVmcXINSaWxoUKZVa9KIbyo9yhhz88DCGMlC
CkuhaQhzcRN7EGONfNkszi1pp1NqGlHi+G786UqYaWJaCTfl0M9ehHFGmis4bj1b
VqsP7rHPqLEUZTV+cloUAl7JN0KveYXnAtIBWHHh72YmcxEKUOd1PNXI+J/vYy2M
sEVRWkqmfbpv03TmM4aUGaEP5RRIioUE51jEhcR9Q+ZYKj6wr4QcomM0yJ/dCXXL
ZXgrY2dhC1ixs2VQq8oiTgT+b9L76KZN9WtdZ1k4qOwa8+5rvd10JvAYUgx2d43O
0obojy6zvoNXCnCzUol5q25jfk9q4rVvXq6Nprs831nwhRytqgNPqHoc6y6AuuW1
gVGC2jN477KsAHQamStOVAeZhuqItnXUyai9aeLMOVOxmJybUW4Lp//YUsWc3/oN
KbRztS/2pEtx0NnaJqGWzjk7dCbOTAFDIHjluM8lnG829BEw+YOt46FDN53NGT5q
M4ai/a8/Ufr0oVpdlw0Ki+G+QiF4dvExQGM5r196tbVL2zWpOiqrPnb7Xy4cYFmI
FSOxw3Mh3XugFarBtsbRlzljpXIBqU5WbhfuJOyBP3aFVsfPneXUmUqaUvE1nlDz
Fu2enKfkKEdkEAxt7YfWCZjathWETe873AF97VtkQZ8PUgDZjpC/iSRtQYt6ZphS
k1vbh7JiRvp0q/0H9qWIK4FWWmC0BL+yLNPlzMD9U+BZ/7vCKhJ7QEGVjJzANdBE
Gxqvb9FE5qnIch3Fok/NK3/mAqoh6TAjK9nFxJbWm9rXiuqy/Ay9zfANjCrYgYYL
BqxEeYip6/mgkOxPS8YXEyrS0IfiIFUX8o5cD4R1tJIM7d+hwOLnyoYtDT05LHay
vG16GWhxtNAhljaMJ0euTyZcoshqfybIVXi/V4U5oNT0KMdEuP9A1bAo+z7YgiCr
1+YnJt8SBnBrGJlZZEoK1z6v+Q4jPX5PJlBwkwvzD0RHHSjezDcMf2yXOW9RRpru
lVmFYa6nukJKkHlM06Y/GC3Fgk//HQ722ZFaFpWRR0rvXe6boTQ3AxXuRH3LNHT9
ZqbD8bJi9W/y+ntVH5HJ+GUwabiyTbAW3o+JzSxuG373IDEqtVkK+qV7wLRD6TQQ
V9Y+BkiFl71KyC4g9D5FV+Bvq4Hfw6VIB3hgklBz0nfEolDedmrG+Mceaw/aaIfp
q3dajmo/VM0+BjbVGjLOkl0qpmKemkgC5jLi/maBX4yvjKTPz+S+PSSPnqccg5wY
59vJo5RGh6R+/gKomn4Vb7jd8FZ8srHBuPIyM89PxlMjaWjRgrnYFgQbntjeGjMV
V2JR4ERs0DZKZaHBXJNc10+bhrvXIW3P2VVIwOmockLJ8NN2v0tBYMTAak9igCYl
XSyeNkCPKbnaduiiCf4QJAU82L2pfnPnXNO562+a59z5B2AaaJw15PfH92sILO1s
WTGnM5DKjovw4V91gbhDG+N5W0Q7UuQiw1meTBxuWs8mKTFEqkQ6LYzUFC02FN5m
qxLKhOfu2A2UhY+9Ks11BeK+dp8lnii8Fvzq4JXKd0A+wqQ/dRo3S4BPIWmpu4Ti
P9gESk3056+2lVVGGweO24lE6k47XnwM/Ad/FU+n5Z4MR2ofHPXiw6Rk79ciS680
2dxhgxOtn64I/QuOVSSI1EWavLht1+EJdUJ03brvigfkiULIZSL8o76BdJUOgvzF
6x23r4NDWwH5VWEGlBnQyyMNNrzJpZh4+ZGL0vxs6TykFWuLplD5M8umpNvo6N1m
CcSbOy9MRNjK2uWROkvdkM2N4SstDeWRhyMWIL6FDKLGWhsawqusbEX1hv7IyVbF
0i9bf+/XOS5a/djWeNTP/jZDlKoYR7m7xiGX2RLqQWwJiGs1GuFA28jflHQxPqLL
qVSJFZLte9Rf1/4YTl2acoPGlsJsT3QcmBqWWdHaPF2GtPX85WYN0Glanh3JFRZh
gLgBfWjgwVb+gK+YnrPgRpOJjH1lf46ulK4j2k6F7+apaSjUHOpqdu4p2rIbDDcc
OioPXWK3YPhGZGu7+O6UFaExRaF32AeyN961Iu5kw6Knj3WkhtmjEUUetr5Ox810
svzYOdXT3CcS3czxqZ5fdpDgvHVwhv9NMjFkwjh0j06NLKka5pgmb7ii5Ll5YeWq
N6TSVzR0bwqF0ONocZoEFmICDLYjxMVP04PZnIYT8V7ldhLZGgK12nweLbBy0hrI
d9vUGpCdoFps2rWRkK04GvP3kE5z1B2f7+DPJY+xY+4dCXyGtXuTZqvCYrI0evZp
QTDLs6WK3KSGGhlodAZhW/9ptoq20J9WoMxtg1onGcNqjSyYpoybeIh9rEN+8hFg
uAXLAsiU4dm+swO6LPp5OzVi7A/J/w2a4zuRmuo7lpBQLiq4Yf5eE1aQModMK6Mn
gNUicr+Mg8ionxdZ6AjuiLTgEhw3O31cgHK3rgW0scieXL5VJiQjVeZf6SWrcv4a
L+OHRWhF17KUAnSn3C7htk27gbD7gTG8NL8hHYxvQFoQHgDt2RAI+5/gO55mIrH1
VTLgRvF17lvRJJiCLt3sBKLVMtIGrGLSGy4xX/TmuTwkBMrJy9gQ7bFPHzMwmX40
3WL2i4ug0E85AUDjrP0XoKWR2w44xXOrq6Iu849p9E/sMqbpH3aqx5xY9lb62V+K
3tMlHY5G+qFnFivTLRmh8JIacsJ4lAnrh2hwf76GKxXZQAvus3h4wg26lB+oEk/j
z/gctAtylBONiAInbjsm+ywN15rElTn1PbA21pBWAHhGPLHFSsN/JhTS1dMiaBen
2qFh/8arfKGTSq8rCkOmuOf9wM3ikraA4OleGwdGwmpfypcvLXl3rw5g1797bpA0
9P+Bm3Mc7mraWE7vcq5D9FkaWLfKpvRCQZKDprBr4Ud5aLEb9rUL9KyNteXFDAYD
UJKZPu48gZVrE3H4LsEOb03qgRaZ9kBXutOIit7S5yOmwlvfps1Dp/V9zTwRBMot
RII2uy5xx6M9BCZe3sVXqxNXrPT6Q1UAH/mOt6DUHtKTj7xa77sBdOVpEhA8LHsc
3c+6uLyZxP0M0gDAm49I34m/ACs6brbiahsmsZDxz8OjpD1cZEp7onZX88fEBnQM
xRo/y64OntZ60lPvF0OUVKG7KZbhIRIwnf5Y5iJ1jwKgsRdqD0Z6M+fsowz41Ef0
EufI5p9KOfo4Y/wyGTZgNrX9YfkRVtEoIR+IZLX8Xq4/K3JtPmAnmmzmiez2CPlE
W9Q2W0wYPQOf1epCPv2cYH23Llm77D+b2BVcULJI0CEpcn03beSuJDquH54Zr1VX
tZ6+puVgWWClnWJW7/yc6Mm7tUf7k818/pH8RyT8nOtKwUXxnUogbhu0HXc93XBz
CeH7L4Qlfn7stVPU2J02zy7Z+Cq451qV9t3L9yOZDD95BWlN0M6cF3znY6RCsW4T
Dg9k21H67Lea7+Ewlb4ga1rv7EH1vNEhU1qGg3EE2CYHE1ysYPCiFcR+3R5BnmjQ
ErjdUwpJfFRk0C5uK/1Frvgs28IYDY+B2lClc7w8P+ZTKGK1LPsVgtzTEeKVrcpD
vVPncuDDy56aMSjh46YEzzw7WdKcXaFQ88/5AjfdSvHb2mAj48MIfuXesPA9CNlM
vTbWeN+iLOXD9w06gnTHxjLF0JzC3gNze9X2aDIfIVIx2N/zfcpHWRxxAFYdJfDK
yrWRiIRxTB52QICzCejhNCJ14cFF1bSi+vjo0mzU+xOsb2mMq0iXz7SuzlbnVOaq
NHh+vGPV3NTB4YuxckV+jJU7d6p6KIqv4Y6jADb5+TuBOBdl5FBqOVxyWiA5KWHA
aGFwO6UCqNaGffleprXhRowUxpe1actOFryXA4mpQEy1itrshO1fmMetXT51tWT4
XAvOzablm17nTlu1LSACU57Jnry5iop8m6ht07BUhU/WS6Bjj3mGIHewltT2TTt+
SD4V4bOnDJHv0q4qfeNhZhRS0KEi0YPsdhhMDYkvFNTGKwH1tgqCHXU+9TOoUFwB
lKcS/Ygam7aggLCrYNuIR/Sm4vwcLkd54x4zq8z1o++am714vJ+jfu7euiveoOCq
7yHs6s5f7EuRGRIh6i2p3N2Sy8R9hlh2tEE7d4Zn1m5zqlbwAd2ZNTCzBTg23sQa
bwsUs8OkXb3pGzZ0n2mIxf9r6uK4kFgmuo1FaKBL2Sy9iNOKfYDwSpUt3clRY6y2
HPLjeCJC1qQB50wIlmBcgTgtmjmNblhPo/m3xuU6jxXIHAt0Ebz0K592/+nQhcdX
JOYUTqqAKDKbsrf7MSafQp79DmpKqDYKHRSL2JxrkNHXEcvMOMwliZhCbsq3rOjU
MsX1gZPfzDRyA0SIjjQW74U1ZYF8CI2nom7GXt09m27957bHBA4qfC0jTOhyNQbA
U8se91IySz3uG1bGC/W+fvzEJ0lcNxG1KEDS9RZrK3MP16XFCsDYZsNSj1i46YoF
iy/DOepWlgbBDeVdd4TBL6gB4cpuG/TSaKpqILUENrSN/P9x2BdY3aVGHKjAf5Pq
tcU8cFV7NPG3DG/gLHBp4pkA85Pi+0yVSFMJMxY7xjbs+4uAbeBuaA9Di1vyNvuF
5Lmk4FLpQy5mVdpwRMNkcYqOnpWzm8qVSzQ1oY/p4Zm0swRoTdYDPwJZ3j31vnq9
B8uqNf/1dWWlcwxggJoymZrhtpoRDiCdh6U1+MOv4qfR82JCUoC/+ckyDJKrHf6X
AibRk0/46WWlL/lWIKRrdCM1l9dehfCPa1eWU+eK+Nlbhu4FA9KCB8WAO3LINw9g
60gFrRfGAm5Kps2Y295+Lu+PAsuuG8Gc1zTOGed2amkppMWtdp6indoODcUhME+Q
r0icWr/3Jnn3azqQaN23baSG4aDCb3CZ6x/UcUav+4p1X6t30J92fymBBHQBE4Wu
pDOEq5GgM6BmFECqtbO+kiBKCYPMeLNszlAC+29I1dXIDKQHpWs5qw8WcPMWyjvh
OZ24H+QoQ4yoisfvx4Uf+Cuoi8T9ze+qO/iVP2vidMeb8KxJI8ZGjlKcTorMt+20
oLC/rZDiD1cMS0eXx0zbrdi49uzHpjaoPUyLo1rToaNJh6DbQ1oxdsDimoadm9q9
hJ25aIanj3SBexxDE1Ef/k4W/7XdMFU7eRu+oO8fmkLAJIptVUzwYTET79sxQJko
g4uAuO+4lc1bWvnyI7emkjrOTV1AK42TCnJc+elO80B8qWfWH8Rk5akJZhSKjErE
963WHSKlreyrl54QkOc1cinZSah6onmGSj1doRRdunfo+tnG0Meh84ASDLntnaHl
Q7WK1rJAKPHand7pRDwI2dWX6Jhvnl/rvtvK7ro4l45DzZYAeP2gJd12YuV4+jRR
q26KALw8VeJ20KG3b/utv9gMUuro5LqM8D+J7NkbYj2rl9drEtYeaMeG9tB+4g7v
xZYve6geM0Zvyt1/jTWBTw6+RcwSEFo5t6ggC0KR7FFiH1NPNRQmUjDPjKoR7krd
a//tQ1UU8o7DQBfRd7QNzCNK8j+mDHWP0P0DSVFtedsa6A+zXPB86Wenkx29EpbZ
joAA/kBwmcOn1Vouj6dGNP9UHr5j6kp+ZL5CuRenxWyodJqE39xHzVmqBq7hYeeY
YUUEw5t90t45QZYBsXMIbtZjeyfjdn9AqhHvQeZMywFzBw8tbdvzdxqlP+Zq2Pss
omvr1T/607KxZBxc8ppzpjXnL2+D0gB3DHcc8ZF7tMi0yVCDCCeZCB2bKd+fNR87
PIBhIZ85zyKGSKBhgXTVOYFqcZjk/TD8/bSPM778do/LOo73GX7pAdPUmXNrw4o3
Api0EDd3F389X6Crfg5JTHDb7BsP5Q64sqLxF+t/i7SMDA4uX0Gkxx/6QVdt5nUb
2Siqs7rtbiVUs6evPugzbu6W6VkcXCihs0+s5Zxy7dcoUkAyawzmo0fB8D3sZjuo
ovQHw0KtVooQniVXMdG7pUtHtDMI9puNSoJ9iXn3PH2f+NJltOxENy1LtRlB3Lng
QgNDLaeo33wPByi/dUGqUMUxEsbjh4FssF10AgJC8cV9RAr2aQBu+EK3SLtxib2m
HXtV/+ivMGKR8if4EAaM3YEuDNtgG0X/fqM/8CNcvdLKL2tfoTvwCukdm9V4e4eD
7ki5xa0Zfkw/oSjY1Wbhx+NThIWv7tsdwHH2nKrsziDFcaUTXINVLF7ZVIWSB+Kj
XpXm156R9ui2dr49K2DNXsg4g3zrd49dvVPelMmhCW2RLADABymg397VlOoGtw0z
msEI6Ua9fNOk3rBX52TTuXaCfhGC8YT1rWa2VckCRGkX2FAAifDDS0jhth6hzBq9
uTt0jpXMoqpYy2U2sW3Ys0rj8PkVCpkA8HZxM4ZxduKehC5jGosjXAazwX/LbXVU
nq4wVuf8PLtdFY+sXcAghupGMeJMRjBL9319gJSPXaeLe2LwIs6+DZ0X334GpZgN
G7QKm6G0w++bEOXOyr73K3Y/MxqjdLNRivkY4aZUoAVISf9QmambuvLVdVjyJf+G
J1dNRxxay6bHifW4Uf5be9kIMKlVwnBO1efDTOZWqpUvW/RUakPSWDW1ex+UZLfZ
iY9HnPB1nDsu3YA50qNjWN2Wy+mURlbHW/Yx3IvAvHSNuPSe4qf7EAI6c/4Ezg3Y
Zf6xpWY8zMw8ZWqjzNFXL0Q7xZ2UX6cMGSbunnFpeqEB/ZTROR/0PNXXy8G9yfHp
OGLDAU6D4hchjTs54L2xVTIcc7bhX8MIWXRYvma49J9A0wKcxe7il0KoWpVWNHnq
zRPeR3+rbDyH0CnXHHJNWbh1M+4r2MO5srYresITLEKckH7UgGJdfsB/weVnyM8j
fIk0irkZWphvpLWOkkZGMgnyeLwlrNL4YwEWafuUlVEWaPSJH0bXP8Na4NTlHD3v
qt/5/IbpBNq/9v8XT99YsiH3pp8ePsBHVKend4BiVe4/+Rj74SZZ9UjemH0rCQDH
ZVZool7g0Vz9y/Ti5zYmIxgIoN1YUFWBtIJzirkJQ8JmGI5O2VVsylPvZvDV6PUt
jJkFyPxkluj6/nX2isnVKosuxqqsST4pNfczSd6ls6PO37rqQqkPUOOiFSKDf/Sj
VaqoX7g48lu63jzC3kajmfqkUpRfWNG/9Hw+syPh9oCj4+R57y5kfEjDmaIpVpmc
YQbnNrZeeWkllacwDxGcUzjegpgp9uygeY1hX11arcOhHVojY3LPZc5zgSWpVkpP
XHMAWJO+Dhw3E2TJ0xh5DHJrJsOmuQwSMu/hjhnV20OiTzQBydAnJQKcGcR95DoV
payHyKidGtBTzmbdF/J59CRY3QDpXknhYFAiJuLYWPG3j6VDLcX0YQ6u4OBsHH/0
dgtllfVLKPdPm4O0Cd/PlzwM3jSP6ONaDcFOw8OIa/vJgjLrkPazhwcrDrPZxi2K
qfwLWiBBCdvjiTWUOhxmaXh4MnFp3xytAFMctM+JnZXjbW42ExzSuCFFl/cziZft
KcK1xOeMh0Av3FleH6hgF+we167noJ5eyvG+i8BWy0VALyspRKBbrH5lgcsJ/Ysq
xuxr/l60tXvstGP/4NURtG8onvWtaNAbiSEWubUl4jrdKoEQPKeqyjBnCZVvBnxm
BW4l5W7Y5o5LHlB4Va58jTKEuZmkV6iOLAzMf/dbKDPPaE8tAiy5H3/jEO4aRhJI
O3ZUo92RWPOALlQtVdQRtlC13eTUOPWsK3OgkgWkf5gC/wWO0nl/xLykYDspiIU5
jp9xjFm0SAzj6pK6TCLYv5U8DrUS7uoKe6YObYFHsyDeXgMRN5lVI9POMV26jyRb
7MC2ZsrTf805IAJRAPkhIGV2hOU0TBOFWvBBE1lKFHv1uCdPcuHpSF1vnP2OUT2n
6AA2oRcwvaGV216dzO7y4eP5t7TrrUDSh6f5XMMlM/guE+ITOOgdo0ngHVxwL2Fv
g54SNFUejCBtIGS3p0EAVptUcmsKNfO6wCSr2tDvSgUY4FCA08rbiiZ1hsNcaoyr
Q3dW8rXNuCn1rKqa5AAjw9//xYrzYt/qrY6VTf+MmQ/F0FMSITR1JoTPAo98VWEL
Jl/m9rFJZXCRpvNyr/fjyklWxoaiHDTvsxzVQsbz7fmy7EsfOoM30LOiRX5D989V
HZ2DydRthT3pBc0PiCd1FLpsFcUclCyH6zaVlXPjcXa2Vy614XoRcXQoRc6N5ehJ
YrrvJ13YLPfSOQwV8bxTewBv4az4jK/MlGg0I0WF0gU4wYrMsGgG9yzvKeSmIZta
8cXzxfM4Ha/qlzheqEOf6YAjwbNic7QuRFl8EIBoZuKGemh/oiHk/4vVvkBrpGOi
pvfh5h2G8TDxITwwXHzkgWNqL00yjnzLhhl589aSkXRjzS7IhcIvV/SzBsg5f0zP
nVB/0ahXYyiVd8Jzlj7A0QLNJtYWnJrKpb0qEENg/f2hyV3LWFiHHcqDIbZC6WN6
ZG5ySU8FqhoRaUVeGh0o0bpu4pyK4Vqlxh+9w+1oe7XKtykMw+qC1jB+hT5FK88J
U/v5gHcjFX6FmKfTH2BQ4Zqj0gzoSwRBLuov649CMqKqbkEC3Bo//uqbIYDrUtbY
qNNW6KrxJhtEQefpFEJ+yRRhJFykB8B1N4DCuOkm8ke5xGf/LElsJ/kH9YgwJfHT
MnbMvOgetJOVo6+mwNa/QzRsRO+8tlHz5A+5bsSZmgpWRiQnM6Jlc7mQEbcvXcGa
vqv5sppvN+mkIfo3vpQznz8vNcpiYq6mv2v/inYXyjYx6jxIuPk8RenSz5IuqD6R
fFC/qWtSM48Pnxt2hsZ2wOPIPDTtSJ/qjKGqhMRaNyDpRw/4CgbHjdMq0TR/E7rD
+JLiDveIusdC711jiDOhx/rEQfNHyhz88wv6MN8/D9cgwX3RVZGX4zexZj8yRD1N
kmHOI27FqMPnFG40SwTaF8xelERChvFBKzYMDfetgH3buiiuYFC7qb//0fGg8DMU
5agdt0CUXgERI0ZHU9Xhggsgu2UiJMHO3wUH9QmxI/uQkJBiKdW2J0mkYfK32IoL
HhMTQiLI/igqYTZ1hNc/v2i7wH8SNbt7vK+3kD2sUF6tz+1mRhOgIBAudDMcjZwT
NTgOWZf3Pj08+CIv2IUY7Ew7Cvj5NJYIgoGCdC/MLKZ7uU+9xJKgsTnEUd6AkHBe
4H+/jOiE/xQ07wlIHh8mxhLLDehAENPg5XItnrfmePpCzydbCiBaQ3tkrUFPbIul
2hsnVVKGbQUkEQwoKqs8KdEhZhG5dY3bjw+nP/dk6HtLckx747yAn/KC8V9WsMPC
5WAh/sUtjdwK74jMy0RI83YsV0anJ4tOKoOz95rlCv0q59J0B+IX7O5Nn02p5iCD
lCwHqtCAFA5HL6UqHXJGrCmPGrfKLrvrAVU/HephwgqzWvYGH9sKZIT2Umn/Nl35
gwRrr7S2OjPUUSIb8BFfW55d7on/p9ei/y6AtqA6LZ3UtL401VswnPkoUVrZhD09
3DkigJkOQMenubBwiq3YhVlvjRzGTHtmQUXv3DyWvqes4HDsM/fziNHlZRje9pYA
iQHRwCVq5/ldBSTjgx0ycnrjfwFbNPRSPqc7GonfbWuAywGg/luqT5qP/mf8V9Rg
MWpR4lnq+4M0D5ibBkXz2u7LLa5kQZUOLXSyax7qZQXpgJELXCnaMEkSpE8EeuPz
s3NsVbKONh8mInjuD46ZPFN7qPkeo0qYf2wNzEgW+9zrbHqkb5O71JX2TYkRBmod
uqaOhV+ck71WwnfOikuQ1FZ7ECkExmjLK7nrvVrVdU8yOIlRlV6J4etN/eB5X0ct
uYqKYNXFAOpB/z8gKkPnWqw6YlQydcCqWv4PQ9EFNBSHd/o80PJP1Z0m5cJjkfB4
sZnj1QuwhCqkkWw/8QbmCufHs6hofBA94cD6NeLMZoG9CNgHv8AXPHEppBEo2kw1
2ieFr00nomgFLmXHVlOuU8Qtoy5x9QyuCQLwb4Qf/iFJdv7TAE9+hLMBKnKcuJj7
2qQMHjL6oVnEy+iiW+nawRUm57whzKtwkzy26VVNgCU4UdyXy/x8hFvuvgX7qk+q
ek43fcFqt397wLGu4lvOuD5aWF4mKKoWw6ocH8Z2NIE5fMHZwQPAFQbgUMUsoHXZ
rPwF4+SujGt8mo/29/KugBqczz/PTmCAO3XU84Df2VwUnfyq0sG847OMTyVk83NS
I6LA4sb9LhCGQkkYkCgLsuLZkOKSz6/lqz9YSAwm5qojn8GARRgdEmSInryDhgpU
ehowjK4dI55/1ih6UgE1IdEfvBMJkEr9xKUEDjAt0FLVawDLFHxe2wHV659UHISD
K7d8J4St6NbqhMDGiOFrjZ0teTtFVjydhdcyjcLiqHc5foaWuzOpZrOhVslW2VwJ
z3HC/RJIv0zVGN1KIvhgOfudmIKgmmZbzSUH8JjJZLHI7N9KPjVYL5kBHpX7gooA
Yo1rE9+tHsrZmBF/5vZmStepQUD0Ip4ru4S2b40Af7vSYSGXtJEuSbTFo+aGqAX+
Ig9cMlfFhZP8PM2RphD2rcriyZG98MSp6lx7ZXNEqnpL01aEvvCKIghfcXuKNHbN
r8bMGX19J1+1o57CmvHL6OzdedPDg+quYb4Cw18ZhTwPnRbzwymlFgcOcglMOEaD
LPF1RXpFdDwD0dqzxov6Ec+0beGxaJhEzSGn66YGR9VXJ/2c5XkYxH/5SaSihvDW
DTZbuUC5jahUtvkQJKCUoWkwBu8HcFm9SO44iz3g2tzaZ4x8sd+hDbR8O3azHTX+
0bSXd78uG+lF9rMNUM4Bt9s20jr3fE4KvfZvB2WtpElt1OQ6AY49veP+K7bOpkZ+
1rX06Gg+YuX8flLCt/Z7DidqlWukk4SKBk/kGjEXlqmY2eIbs3tM5FwIeBoZZq1e
+9W9Twy/MPzVq0ogztmFzAFteVEVsBMdVTQsdZvwpVfI3/DEQTVWEqiFjAQo1QR5
QOlCqmAAhTcxa3SqW4fl16Py8FmfHHGNya83g3akKw/ZbbXl44PuUzIf6zl17QaV
uOh4smJVFvZK+Tp7cQCIWF+Ys4rjavENgC4poqaXPKFbVF/SRU6G6ft4epwzqYCv
HLtw7Hm6DYzZBC7bijLvh1a5A1gCrpo2bRnZENc0lG3AICorXdp8EGt0eyUejrQc
hHq7xIZPvxk/VwTFK7oULZ59DZQN9b8MUmP/NkncAjyxBr1yhfzPFJTXvEzXsOK5
Tkd6wGwXGNpEPRwzgG0ouNsWM4ZfBaLRJJKF8Ja9Xu89WJ+RktjxWXxIcyZXMGfL
IBW8nNRt6TimBeNZBGyLbzSWm839JGmKCfI/NLcMp0a0Rd/R4imXZpPOw3NDGsUa
hPkPBr9GePHECyNcsHxTaHmbNAwCA49Nomf9h5BIVCh6vxpX2UgdAxPVrD/1fB9w
Ddun4EyIpuJAaS4Xvo1j0Kf3vTsk9zvWWr3rAhMwH0fhvavK1KPaOPYFDKArAMgH
O6Y9CHDli/QanGhfFqGZuADtgm03/Rsqmvsg7h8F3wf0E7flcbQNKhuD8hn1fi5y
E5NB2wHm+dIOgDD116xfjuw9RML8IhhIfWYTp8k7gtN4n1ntWqcmqx5bzIHrQVtF
OotRDvcu6B0BJIJ3HbjLnWlpjysJ5Q+rrIIS/tFSzOicsN/66PUBJm8iPPamZwcq
sBbglq53lEKdFnbwU+y+QR9GkKeCT3Rew/Pvt8W03LW+gBqbBeH6F8qUF/n+Aq1T
ogND/0Ex1MYEe4yeKurZRg5NQqoJ40A6Ed9ATjWJ9DEIGBGVsOvqqIBNeGu/FhvF
bR0vBYKShhGHqE6vJQfo2X4wvDUJ8F9H3z+yRFY1Jlp4ujso5XVCtMz06SUyHzo/
a6iGo0nZn2YRlaKV31sn8voNwFK6fzkurjpW5bQkl9Mfv33YkCvQRpA2SQ6GXYEp
bYdMdvfC0GB4FeiGI2dANU2IbF3/SsZ3rtGJ87++zFNCLHAWPGlvkUNoQkhksZa2
/S/Vdab4jAC2lbL58rtblZpyvr2ZktMdYxKnYBS4J6JLOKmnHM+ymDQMcVK4PRG7
WS00SXOEKj6VIi2O/QyrMqQjLw+f7XUr2DQRLTq2+z24LBwWEiP2bTpgqFYhF2et
OrB1oCzX9kdNhrO2lsw7ibkxK0KMiwoBY8EpJ1m0MMgijaoaudGq1rMqgY2w0R73
Wbz1uOk7eiSeuHf/cXqfJcnlTVBp6p4splPXNs5G1BFpu+5bwZyG+1g9kv/kTgZC
P4Yud3dX5Uc7dONQxbuwaq2IeY3AIwghJbRpLK7OhI8XJoNNnBFwNjLs4IWUdvRl
gIx7ceNvG8M1FOyYMiUe8NWwOoQYIdYDB3nHc/0KSSmamtZVrxFvblXRK0ruIzQw
/5guIrjUJpSClB7yLAHVRiL0rTVeV7FutDz8/84wMOMueEi78xIJmXVChWzyDt5i
3ATktuZ0p5K46oUgsW6uE43JrXCH5tqyrBwi3FTFfp/YowrYPac/3TjfkfktTOvY
aYUlbYa2dom+7ElNaF8AksIkS23vWDVveURePXjJNicaI/wKLwtTIk6Bt7oWstOx
P1EnoCRJ8HxRutCg6EaBJ2ed4mijH10+TVwPEHRgF7WMYV0FwGMpVy6P/oqHevqS
DVkQQ2Qx6yh0ErgduQnywjegMPUXaCL8EnxBtgPitJCYUWet2B4Axe/0sLbuAvUb
cZI3GV1Q5VOwH/MCUFTnP71eZh0HbC/xQW8ZnsROZD1nkhgeQztldJn3DDLVNDrM
0HI8sNycxY2oKWvBsUXjlirNgpGc9zU72/+q2AsXIFv2Ssh9wSirQZnO9mjqD4N7
fdT+cGi2x+PRRx+iAUpBXILi/mqD0Tg/l/yG7d5xVN9F9Sun/Zhs94bDSCUqbCCd
SKPN5PNLhS0zAtIggyj4ggR4OM389E6zhlP3ULYezZ+XrVAW1Vg4WFUAbr4O66ic
wFmO3hXPu6npuSc/qFKnmcf/o5GZzkDzj+C/dM1JI+TohFhjG1gw8/wEGcRm1NBL
Ta24wwiG25kaY7jFyDp/s/xA7p3yLtm7dfk9KQ1HmpCLfWS9dH6UdsXV5qKGdT/o
04m3J3FQe9N1CqwPmWLwoTU/kvtouAOj9bE65i1s3J98/CsEu86bSAqoLV4S2dt+
m1+3UG1xum8MAhvJkaGaGhJ0Hd8rILc0mhv8w1oMl4+ZzB5CIIB99tEJTHDXSFz2
Nwr4lblFQ+Wjcc6mNwCasLF8AxmtMISi3aw0V8KHVfnk0KVEKrtWiNtwBvh0LoQU
YeJufZ/+nl1ccP2ZvEDZpWbZQb4vRGPeMDrcl9ewYuIzCJU4PAaZxYbGbBdhNMJ7
MZtZxcrBN9H8DL+o7DhNSQdi3QdZuR9EEwHF70a2mlc4S1x5hDEjF2aFFNZJg8Wa
gJyWJ0NSniDPfqlE2elGW7PRxLFGR7QCvZCJpN+YgTMX3M4b/55DbZXInfWh+uf+
xY9DxNWXrzn5drFx4shF3rnwscAkZfZzBPbpuF4E/01eNVb5jFY5xuwNKuTpd6Ex
mihAQGtSjnLQSt+Za0WaC7L3YjDm6xLAkfx/KQ4F1/s1ZfZcdKR73uCDkW0WSIfC
+SL31sUXCuHn07aXqG/xy9fZ5KzCJ5LE/uiK4998QiJLhh9T3Do0cK0OBl6ht0Gu
hXATqVkXnkWK/8vuhdq/8maRaOs++e5brrIS3tWSaKnJqhf4jw6/xvZuiNolsEl+
4fLZ4c3xDx2loc1c3v1jGeN+b8qJqted5W8x26VmEN5bUVUUhgiDheE6fW9XoupN
OiUqxpl8xSVnWHc6BMJ2Pvgrx5pg7dCJFqXoBGE1a6cgv9GY+FpaKieE1vwiiMr7
cWTRSRgahtiUf+8z4YgT8Iy1LLQykchPZmsouMrKzWM1yR79EwOpYJAmnsLAb3bH
TEirAqfEdqtpw1rjx2asDIOk+wWLFb/RM2c8TtAinqYHQezqKqjCsrMN/S1GRH5Y
LpynI79I2R3xm8qGpE9G+iFYq/v/2z0ZDHeTXJq3uOG6jEawRJQCmtNBmK8I4Z1H
d8ptqjspcvYF4tr9YSa/hSgRwxBaoDbKt3Dvkt8PwUryk+H0c3OkOk9MCR6qNFeH
Csr6QbfV+qyV+e0wNEzKBlRTaLs5su3NFkx1g0Gt8B1FFfD5/G0EHW5gql+o/Yb3
c6uw4iWTwY+XaUcMDuagek08dJgxBlrtBPEq3O6/Nn9ycNqEe78yut9fYt29tr/y
24DaqNCsYTz+d7x96X2M/C9lSGOX/1IZ+42naBQeP4i6o22aewCYBrwV5pd8DALQ
gDuD9TaqwIHBOgUe8NjT1P4RTURr1tSAG2/FwAAslgnSQn+/Iady2xs4scYPzuIZ
ufUV8c04Kk5NS28Zy20Wzy9gLMSP58ixVD6ffMUgSLpPOM5+EYXsnynB14j8YUwJ
0SqhEM5nE5x2IUdh8qrK5cUMtjTKGFpf1rlwpbA7rTuCrKnEqhcyLbVdWiIAIBJ/
VSIvLDXbKqhy0VGgV8iJzYW1+PkWTWMdQYyN8KMncRhQn1nF2VwcWPP0pKH0arfp
RQ/w7GrtEiiC1glCJBiVQuWKU2oYDpYGdgY/Wj8MnWDMhoW3AVyzX9Hol+E9iWRT
cUqXUbN4g2WPz/X9el3ibGvV9uwyAjtgP57iJT3ft46/Riqaf8x2HAP7hZtecnMB
ycbHfZI9JvCbjR+6IOxFQfSfesUCN1PZ8+K0ZTZQSvfE26riAnP/d24DAz5zTnSc
WCDC8KeELxM4ES58nvujIZPk1A9WipA3Dam0HuAvjsMhb01pxC37PSwlUC7Ar1ms
ABwLZsobcIplJSwlZZXRfezaO2np8czmjcO921mbQt0mHwORCy409OBuIRKyDMok
7R1sQ8WxPqvDyqALn2B41XFQznzyVAms08duy7sWE1bPHt4wzPgoJsYzRKwqSXBV
KfCa9KatLJrQdagNu4QwUHrTeS3CRHJMnacPuVJTfb5u4WXt+FQIskuq6w10xATX
lmq6TVz0093iFp0ndLaWmYbueHzghUyl7YDWSde7RMxXYsB00S8iMq8IbH62lSaV
qjFtzMf3hSvMKiml2dPg8ntgCITK1044h8pIQUunbF7DVJBdLxDryKcXfCU2GBaX
grVOlhLtWmLB7+kcmrYFUBv000MttZcJZe+W0FGhvBAmMOrhbTribp2B372MZ73w
WzaYbl8k3xXzdfcKIAgdcN3bommlFAih+syt9609evGT1mqqbzPYnoycnApIPA74
k2KY9xQndcpt9Ju/MmS1xO+Tvy22vDzLv18yHsDdWMC6lgpSukV8Q1Eclgz5HuDw
A75f7zK/WEM8kPYcaMar/nq2cGgWfU33WUyUrhY7RAE7wsbaotlWw22YDTMYGhln
yXLVg3za4LPUd/kfiou06J9luKIfZrFiScorlBiu7ueAevF0u6H/nMql72+ZBYkM
7+ObKYJuuvfH7qJOK767pEx1099nbskrnJuqRXTQ7w0M51mzVUvJptF7mh8I5v3Z
Hqk20aYTZmTMHsF0ep9ihkFwAosWaxui/1Y9+aZ5wVA0ztudWlsfvTC8hwFEA4SU
RRita/f8/6i9m0HEh9FZ5FB5a+DJaYT2xiZbcX0waSGDa7Rh0uiqQrwge74M/doB
9CWJhCcCZbTLp8mg95O7slJIzb9HgUEXIOeJCqqSWwBl7zDNgJ+PQz2/6EagOtNf
/UAiWy1OnWz6qTFsWUK4hKPSWOzGE5Vo+DGW9kg0zCyGsXe1PiBQc//XKr4aFwnW
ROfZU1AtPSvRsJoX30GYTKBfI7Friw2xHI0JT5liE2JSM9tRNTJqRLE3e9umgDvd
dwva1ESp5X6ShOdL2hM12B2wzQjklyPU74HPzTbdKuHVIVyiLUpdX8dO5+98V9/m
cIVMXp1k1Ex2wTfqMvzGuKUXzb/vv3qlB2p0I61dbKWl9nRztKqci4HKVjWteA57
HVHIgA6Ss0wHJE6D7Z+kHcPMmQ1pdnvdpiokiGsn2KUYghgAbKxZh74nzyTMKFDS
SbfOBupba8YAwavgkqlTQ9iWI7sPQzLbOb12A3vf3biUoy13SudT6+uXBeFD+UFM
dYz5hk4aprDzRI2GmgbWInT0mDgL7XMlWZtNNg5q7VgYaBLtdHMMi36pyolTJC0g
Ip+wsbva/SvubdoJmdRByQCfZV6H7HqMKM9t/qxfqhOm7eAoIE3lTPJ/J8haMb2y
7wDQ83QusE1u2doG5Oydv18JSyQOPQYXPSoi6F2k+vAek2HXOv3xTp2MP0GboUlh
gprRHcUzbUv3aKq1JGyQ6lATBydCt38HA09N3CwryGd5L0GKbBwHTPnDnYz5AU7F
3oHrZcZ4ZXU5jNYgTOmrhxBUh88AjzyVPsDghTD62Z7xoWI3UKp+xUC9qdGFaMNz
a0OVEc7yrHr3dITgdNiKTL58UKKh/vt1ikHwz1LlCiuWO0tekRPg7JdqtWrcYjlA
bpi/NxRAW5a8KUV09kMmsAiRnbFiCMuYUEduF7WZAbhC7uBIhmePgC48rYdrxIQu
WbCTJQzKFPXxWxtTArBvV6MEIPSm57aZldB8heQsn51W+J6bQJn1jEsdG7YxhO+B
zQbN6GtDo6LqEOUDLsxATqoAcLTbIU3n7VGF5z0ywIVgBWvEp5t/3hEsevsdnwFZ
f27zd9Qz4aWKoE38gOQeH8cEvzd+BM2yjr4Vha5j75EvId3PR/cfuAnPC/qrjGOM
yNLmBL4608IA7jNDwxjtB7GRWALl0jaClM5UmTU24fxpkG5OZN593nIomy0pEXl6
7tccHP71LvRMXEiBwffA6HQDNv4k+86a2Grk8KuF0LWpf9eZ+BtvKjWe9yIq95+W
HR0lnvWbgShBdNwYPuoW/JT9Qfr5sonTtjYUT2iKqnJLFYCVSriC4EVdd1aqBRSq
4q/owqKYBd80Y3Huwj5Npws4bwVclR8WlGVS7HrFWze3WA6/Zw5k0Fdfr/RN4DQI
Yaske8v0h8epG/q3xQEZYPbRNzikmXjxEwpiy6RB2fktart2NEphOKJtM1s8GfI0
u1bvgvMXmLMMD/WSjzCaYmm5Rzu3G6zkPDs2pdIt5Rq4QNf7xgda+ALO8R+5T0hh
z1mXhAP1wSixYMYs/WpGw0ARRZyJgx3cnh7ivSJP3rJ6W6CWiVdxVCbmdRjgd+D+
RvY/PIwgHbPRHP3g2j6VfWpDAiF4Vb3ciS1uhLQF/sBXGkS1IGUTOz1O32dQ2APr
S/WGoFgNMoScXfzvY2bu9gTcuiAs/b4JUhvEnY0apXK8S61R+71TvkGh+dswAxhH
6YmDKq53c0iWuRNpei+MPjCSsVrZc/Yla3Lt2O/+2N8uqpBjU36QwXMD9taiHVoQ
1osI26iK13hpOGJ6SoGwSc3qYIJlOCA+sACkhFZ0t9pPu812To15nDB34eYqNDS9
2GLwfZo4EXy+fZyg1O4krwSM7goAYNzA5LsJyqA7+JuE3JUQJ8djX5Du/jnQ3q+t
qSnlInhRsJ+HpJILODXmACVr0bHS0tG3E4IrLCq+BtBg3gUfq2VUvhwMUqYHb6Pl
9PRiQeuRcx87JfqOCinUrpGloRuYV7G2scuAAsZkHSVC/EuIQuK3eNUyakF2J8ZL
7jSbXNXyLLGj82vv7orpZfM8iCf5NaxQQ2oN5GqFDbNZaa94TqKG/7ja5ZDL4R3l
pCR8PJOt1E/DBJlKN5636xmnsMHhPJ0C6irbCyi4vsqWC1KvYwOiz+o2oiUjie4U
SslHNL1k1l9XoMmwmkau4QizAA5DpPoz046Jr5eBAqgDMWr7Ke43g5me4I4rdWi1
bnwIXdVRZCvPAjnfPH/Lm6TTbloQM8mWVU9WcYtLSqA8YMiQ1IVjh7FlCyRegU3j
UC8MVN+n+0uu8MVdT0UtrK6XIDM2RbU/E8vgmXI0ahUqysP+6aiR6rQAB814Cg1F
dMEe7O8iV6zYoMppdzb1GaDqolB5v/IS6EM41gCBIkpRyrjN2ZAytIwRHMg37aXG
A74w1YutEDk97oCUsSSZsWbo3ptI6PAR/+OSkNIfaeX8zVsR1OBWsJ9hL2FKTxYW
nHwvnx9rikpMl7KbjU0pg/0zDeWR03LEQLsXOx/efqHb5XZCpiXTvvZZSvI8Pumt
iPu4Qvi1KOw3UAKQ4i1F24tawTt94VbobI34PuiUaq5XTGlFoLJmw9SzOcONKF2K
QuM1BFDoWCKEuO4g8RZuwx9FHatNDCciU6I2z8u5l7HNYVvew56zWXR3qh+hpFem
kPoNChcOL65jZQRXyHa44KaBSbm23mOMfJrjaoRya26OjrH/3JxlCkBrtQR9szt3
ksk4vbbYRxtqw47PDw5ORiXiemi7cmLCP/st6iSsdQ31t5mYmoYhishVqwAWIt93
fhKK0paEGoP450p08mKAa2cIYSsX7rvlUT/14R6DcRIKlGz1EQzVLuygzGbEX3A0
UnEwHOzdF39glgl9722zacmhRuPLKKU4+Qse3wUlLN7fHmrm86O3V3nqQXvWszuR
RXERD8cgYBeJtXcApuBh6mB403YQ1sKzIfK6E+Vm0GXb7Gy9TmJLEaxtLPxDRuKB
d6hTl3DsdIwtUIAdKjKh1fIujWQq8E92NXecEydSrwYSkwWfheKtyzRr3MDIcYEZ
X0ScXjWv6MRmbxMDHCjEr9rtsfmATtjps09bLZvWTDpqgVZ3rBXltdm22tFrTN8e
pVfZvg74y0ajMxStA9SPULFHtoDIl98DDYh3Wt4JR4/zekTtkhS1hSRCnCfgM+y6
IS1N2QaYl85X/t1ErBLNntFyeUtWEnNxPJRcD5glaa66Mh44DveHQV+q8NhTLUQn
gWFtpwxn8D/IHj2rtNH0oCACz8q6HxM45rlUqHQVe1SvlJYNLmu9zLLgSeEDO0h3
z0r3fInsUktsfvxwDG2lwOAvjjOv76ge3ZyL6mCp1UPVmeTf2ArI1assQPckxPnC
hQ1fLStjbTu7HisUBQONVFzLQlxqCvpZJ5rsctEPS0aZQ7sqKNSJn7AgY68JrrO8
gHEbnG879CebBZUqSZqOdTvel2+FnrGLsF3p0lAa7hbtKcRa4Rhn9zjyJgCCK29g
pgldZUt5asiWHa9NlXjZLg70TfaNbR/MMFLRxbDpJELZ/B58Wr8Mg9p3SXP4kpDG
DMRARvwgl6DPb62VOESUdtqJPUKlxzZGJQQQGoliTIDepBWwDQL9BdPx5trrBX54
LUr+t51zVfIaGpj02tsy4TWfGdQreYDSGCr/3vuPzukpyU6JW3uOrFSAD05x3N+C
UVfgaNW9rPOFweJbgK9F8PAo1pAo3OimR7DWZy4ie8H5OLGAEXPJhk82tjLYuOhw
iGgmCdPvJ1tR2FQi6ZiyVPxHDcEo98txtdRsJhhyFzKOCs2SH/7eX2tdxQCDkUcc
bECSUckDXQ9uXJvjFsftKuswV+vabGyjYEio5MaxPjJVY69MJXfp4F58HOHAhHPX
XGunLpu9sqK4UyyToqlwOFYfRojUtixFHS3OAzB9Yh6X1lRp1yH4F45KlKMPnqrI
UxDl0Xp/gbzuz/oTiRlZ3WCni7V7A3YY39DmCl8sLZOhjYVBXFRu5FVax+VOceJB
jCcq47I915IJTUZp44+myzoXXwMxW56VH4zwYnt2K8SocXYecCYZI87IynzkiuKM
GG2OiNvRyXnPzjbRv/Vy5z070kpJwu+baldRerohB5tYPMTeM48kMJItiiz/ggp6
yC0o3qi3SLmz30gbLutSjRqcXX9XBthfaW+hwCHf/tMOmNzUQWWlMmhUQtC1LIjS
49k2pne9uG0mdbXWaoBIWlSoqFOajUXFybsjSKxLaIeikuz2/oFM8cBlzokme1sK
LpLft1SzgzFFu5tyjLvrBK5d//YContFzLQGquc1bVgTlEJ6PCWLy6/uqWBkAaAP
xBbVgnPwWitUabNpb/FEChI1yXVbMXSBqtAVmGGujGP9uRa18BK1eBSayI5tFAlR
X5jUTtZc8S7kvMi1adpfiOX6mB4liaJgdYNmOQSmmE+/AAFmKMEj2yRhNXojcN/X
jHTd5PHOwOdYc15pqzOG35tETVSHuKyNbI9vZcFpsYDs5A8G/U+eZdT1brqqkkgY
C4PZbPqLReTvcxXWfhQkMXg0jP5Y3RiFjgscMdIkHu42JghYyxSZPdkyTI+iKJgi
ZMi9G0ARsK4DKd3Llyf5BZDmPOKxkiJ/ClzpK41gyQoFvda9ylnLL1RECGA19LAZ
4UcjMlREzRMJuvk3iunK2RsXDgooiOT7/uPz4JNyjUGgL9xjyETYD+HywUUgq+5c
Ac9Y+BkysYSXndk7+vcoc1UyDURjGooz3lNREdKRknD+gBuN8iVFONB0xFUwdpyd
AyDckiNfKE2OkvrOHsyRegOP8j2DPd98s8nnD3o7Lj6ltX8v0wItBfSjUR1vA6zB
GBS6S8Y5OVoXWEw5di/eT61pCxunsARiTL0dQKRnEYILgr77lTErkwbQc6XDkh1E
h7fXQIXHZCmnKERhTXe5KpXpfDgfW3yT5YLM5ysIhZml4OYzd3X8bvg+hlVHtWsM
Nxqnw6Noriz9CQw1nEoV1S9knCwQgSnwVY9OxKGfBQuuKKV8BqnMG7Yvw9xr8JNt
vZQOFoTJetFGt5VsnSMERPAlvsx1zsqsFooiLyyWIzHKYeJdE1Nhj6dHpyiNXff6
h/F26jQbxJ6vtMtGZ1oL9qu28JzAi4wksmY7DWhadQeEPNtLtIWHE36ORa2GhUrF
WFKtvxIiDLn3WSESX+D59K3JzIoaQONi3GKCJQ76s15HfA+0eTVLamWAwQtz5d8l
rUn4viJewtaxd/gV9TyiwjftCbtb+TNRU/h1GZIAgumsIE/H+JJJQXwe5jd7kNnl
uFw08wEo3Zmxg4rALr+aQolSp6erx3Iz1Wh/PTrSTMEM79z1YhjsnN8aFIxXax/f
V77mVGOYIcs5LvZBuqCkUN1dcWDX2DUq0OvbEy5a1/6cK9VxoNj/CDD8nZcTdOc1
LXXOaAosy79/kQx6QGnRxuLzSgenddFKQhKrf3prZQCVt4USDQxzqJ40BZVFq+L9
NsUs0GU1qbe5yXyhx3P+2hJCLAM3Sm8unB0mCTXNgD/H7lrTIWZfiF6Gm4VyJ67Z
T9nVUzk1+msnOjm5Ehb5PlkRVYaUyr76xT2m4WN478BYFU5UG7rjPlAViqMnZP8c
4EvnNqsbIJU8XlaNRDcuMDOHP8aNtsHbnJOz1r6j3K38ofHgSvgnLrG+Z2CP6lvH
HjpU5J2OxQu2kcdL7lb21jAH89fHHINYgZonrbQfsIJCMUgTZan7ek+ZXf7945wE
kHgTn9NwvfSjdUG0RgKdj8PIrYmmpQXFxr2sk6aDoCA/KOFhHE0CvZaqJkOEv98i
dDmnJGxRHQgjRw/PG/yxpHPecIkYVF55WjqHeBaYn1FgiULllgv1vngxZYyonR4p
sl0DNSuuQwR58dJBEOisWk2JA+O416QdFM0gVuXSXhrFJ2+nfQqNnobx0/Hzntnd
fuYCz+BCUzXuKK2/mleAnJpH9yKNfctTjB9+La6k8r+7SA/9r6BiCQpovgybO4Gm
xtgjzDAPEYHIaWL6LK9zXjFWmwso0N0Wc50IbAU6NxOwQBVQ04MN3ElY1FNFXQLH
U83s3x+1YKs4HPA5kFr2TYOy+BIhPBlyrSvIOoclmJoCr0uRBGjDWdEKx6tgS8rY
LAlIWXAR6BoaezmklIRouJBABcZ6rSWcKWc72sXZLaES1WkB+WmVVW0jsyDKEj0D
zfJmxtz2GJ3QLbAhO39hsPwsjcTCVukfIbMevyk4EwESw2sk7SjhVO0zyCpqkFn6
9Cr7I87/QIN6Ne8pNYsIgkJDNNtNGNeYtZHwgxq9V3ej9AwwuYy+em4DfYZhIcNB
OFvAjfE0gNQxuyp+wwHBK4rmb46S2hQpZcV7NzdbGT4ZgvWJu6JUcsxJYGhgZqz8
juO38dtzl+dRvPcThRH9xAkK1ysKJMBHma89NGr8VVYWe2/M/cSCbPBtsPK9HqVN
eIvsF83RgSGaPy+8MKDpdvHmhvNtuBI/w5V+LSDeiinX1zOLDH8IUw/aYKZd1mdq
b90cZir9lU7X+4QEM7W9MYVTxflQuV31w/tknhbXTEnEmKYtJmyUPkAHu7UO4EFL
wT1DpUPQ9uD9XWBkh3FyN8tmlLbSzBautuFQAPuh66ZYCnVyCPB89nE86+m7hD1E
PrsmqqMHXhNiZ77X8KnVmE8dFY1B0aAYKOClSlB+jjdXH4l7CaC1jJgRszxHodk5
KUF7td4snzAgwBCfSykI/LGvlM8/dZoryOJJdXmBqEfAeLmVHsxP6JEK0DhJCN5I
Ic+SkeMNXqt/0f/rRjmggriHcSJrE/NCTUnp9FdbHjW8v1cse6rfjZgl4mqaCHP2
mXtiUiM+N6VH1w6jpWc4G1bD7J789azKJSp6nlc+XfeoA7el3rbpKXTYJVIKmVeT
DLg2vUXMI7hfgQy9n83/di6fAHKR+0VW2fYmFrY7csHBkVyYu3nizvQZ1rdaA/UE
oZOfkMr+h2oBB+DljDwc2tV5gm33i8Q1+ujKA+09NJ2beT3Xaxf6aidJZvWH5BNq
l+gJXDVRwP55p23E3bfPitG4vzQIfLTBN/Glk+dTThK//Uy4UcrhUNDGe4zg5p8Z
4gxM6gsUH+XghozOALUQ/HDwSs15lVDeK9nmPqXbnkzw6qIKu7WEfXPeg+nIciKF
M9byF+MfXvnT4IaPC0Pq/G3BMMZxH8xAFd0WpKat45Em84DX254p+MTIfYCaxlHi
s6uH/f8AuqTC0A+i8RgaQv5IjHSZ3GTYH1+Wpv42vCI0rHsAP1/++RqwsNxZBeox
bdCrg5dwYK9xjWJXVYk4WEYUy674N3SN/x08xt/juloFB3X+1VUzMZ5draH30YtR
sVjokETiQ8IOt02qdm2pcSlz6hFZyobcG+sXRaHjmauZKBVCQyFMNsUvistmnBxj
0D10B43yrdFemkbzMLWf2+fUje0nvcNtlDRIYlCyZEHk/FLVVBP1+XAzdB4M5CMN
RmSc+eLFH9eKpPnNSxXhV/JIMBR6xUrnBXiIWdrBVGh9O7ubV06zhlPDHftnNdy1
btr8k03AWxBv+J3al+qz5JbquxQNLvzhYgYa60T0sQwN02jj1DvKmvNHjLRSZ4oh
1Ndg70mt87Ir6DsvERIZJ25zShWr+CwO+qTSYZb3cNrI0W1euALnwNC+uLKa3Wci
Poy/Wr7ltYVNsN9P6+2udbepCr/fXmIlfeFl2u4rvzmvu9Mvt76GHxPHFsdth7qy
XdTd2DIWE/1pHGhvalycOjPsfPoRrOWBh6Iz0Yie/77xxsXFqbtILQOCbjSY+UqE
TTy34r61Pn0ZZWqsfeeO3B2rjqGqkgZie9faN/ycFDfpbXTwyssK2FcRJ1bdm1VH
NdlNlBr8B0z/5g1WapCRKXeSBxnWpnQgy6bCP4zemLRvpLTtwJwWH2tqHq9G5CGH
/a9lF+iP92Kl05kuhaYIKJo0/brf4W57pY6JBI0JPOa8KxjKmkxHiBW9x9EEYQ6s
lV3/L6XAd3K5D5kgdstQi6Dle3v3mDL50FgAZq4+wn/1+WsJ28mdwymivyU9/7rU
3RKG/arGMBYcrQgnHMYc6D98whJeZqGubmIAbi1O5z4LTIeGq/Yd+3j6vEvnadoF
JF8vSkVzI38o4/8L8TULDd2qeFdBWqqGXD5saPX2dlX15/Tb6Jxq6BRCcsv7ctVc
oWuVrRs99HDsevilqNbgWjImGUft5737wy4UPz5lcUGxt9XhYHWamGLaSxknU2RM
NMyR1C95tugNEKaN3lcTXt85LK/v9NqpDlYV7DxqGS7E9Ocn1Z1nZ9QfjZdSXBxK
3iUgKJXhXUA7PBbXwfNwr+Vzx3k6RlFu92Zkb7dJ764rnCNdfa26WCYhCdM4D+wr
zSHLRAs1NqgqSHrM4u5h4fVIZ6lPQMgXcYHW/j/Nx+acwqdJQ2xXPNgzpO12yCE+
wc8gseFbwolQ3Oy0Nh7UgID28uFMtyGLaXeZ3AVymhIAt2vdrz/4DFJ4id47ysBG
wm8ln49J7KYYjE8M9A5Mdkij5rP17Tg2wghpGcSO3V56KcImY+y6rT++KFgOSErq
yqOYPX0mU6SDBMSQVVLgAb2umPbfEFqVyr6sMmL/z3uyTxrwF8cdTwWxp1IZbCXx
oWIaqV+g45dMOxFikCopIJDFY4dRaoxRi215CKCtfeO+2DhwoS5uNZrdd8yPTgiM
tw6EfAq5uchPZK19JRyWlbZ9TnCaCPaxWQsrOiyaZJgK4dRNvT0KMYTTOCVmpn8k
3SeMNecVpyMHldL+NAFUh6H+aUJ8XuQBN+cwTNXsaf+gOXFFlGOLReZNvLz7pihB
Tsh3IvXNmp39BUs7fUIqlx71smhVEqoviWn8SZB1KjTlipXdEKytmM0t1A5bZkgt
hUEKJCXkSLluKxs/qaMLExGMX4TYxA0iC0NPFHFSQicpCrhcGta8Pp0rbiNKf+Db
1fW7bPyYTG5UWanWKCGpMSZ2eWA4+j5DOWVpW6xBzpxW7CEikRzYq32AiWTIxdej
XIpPWFYhxtnn02u39Dzo+vQ6b5xtkfe9c1R8mI2v4aw+yS/o/eZtqbd08DJLPrEa
/tN++ulUJjEw5ar2PYJT32lLdGYAYjguR2PujEo1/r/zJvgMJB50NLzY1qPkNewl
5fvjc0TQkuw/5X6HSpossRZQzBQoT3j9/j1C1ThOOBcLg3MXn1bzEfhYtdaZJcMz
sE723m2zx+FT9YvGua5KrNlWusOjzLY0rlh5HNvYjX0HtDHhSgVN1KGrk2fo8pCC
sHB73mNdKLE4M5t+Wi0+TAKje13O2ZEeTWwehrIkN8qV5bDfjN/oV+H3rc4cVEg/
ztoSXH4LfnRPAry0cv75xxpJD8WgMW2XZXMnKMIGCegEbwuKwb5A7ZULCy271DSP
kXq0HqVyklSRERdx+NtHWDoOzu1SKE/aQ7HEJVuqdK+bLqARqbhcvpfpyPuzdkTQ
BL29Qc7xUz8yDltVSi5mumLf1jP/rlISAgzZUytbv+nC+gc01AiX3Ii+RRCn5ujb
dhUS/1hlMosB0QwBW0qkUSGEaRgX8FARTvQwj+A1gz5820GbXjMxmQGNA1j4XHmh
kGH79rT8ewNT6uaAX7FVxuZkj2aieu0LvhxYM8X/4ccrPCuFv8uBA7t+bXjZbRcE
cHTSoc5pdXGWN/rjxZtPlyGRArGQRugyzQNNJ6DqGzLeBRvOqHGp/VxRqBcCBYZE
WjzVz40p9+quodZp7GTifEl/x7ZegtRaea8d3uriEhB62NNgw8J5K980GyoamJgK
7O8iJPn46WQWaF2sViPfXaJLojly/LPw5SRIvGg23Yj1BCHFWRx95V4HFsOz3jrP
pwpB4akjVJ+gP188RYoKkTP6sTGP9b3Epciy5Fkeqea/XDnX0jNsa5HEijXaVhHG
BBsZcTnQT8Y5k1jYZpFxF3SURbSYtcEy/T80ysSB17hi6DLYDMKMVjOGh1VeJp8t
YHLdwP7D1Ihl7fmvTofkwRI9Cv/w1jfICZ3jyOZ97o3k6Ox06/DpGtBjqRgyhpzD
rUgBtixCXMBBILMxOvb1lTbP8naAeLRzkpgm8BLwAAF5txJik4qShHObKjbitKAn
YNK6ANKmeVnOHumgrT3mXCtwYUrXmZsGp6Qn52fdImgOXswh6beYPW6ID2z+Tw2B
p/rlPlEPOqhyYAnOwBRJ0GF+DBHhLeIFBQ9BXTjbePuauxWdHin/bNACYg/h1utk
aHPXiWxVhqMhhr4/f3y+hUjgqp6TKXWHaqa4YNY758187CvpX59CQ6GJo1pvzMno
ITWWcrJnUKTTnKtjolPpTWAtqhihbrkuwnv259vxYQ7YnrBr/lYR+tE39ZFq1ouY
0pPBrluW+Fy/MNKZjGL7pkHFX0mAdMtsAYLpn/QT0wPf/QSrxhms19ThzYpFmyig
IXVah7XWdHPSZeXvTdh/D37fhr8m5IvnFZsrFwH3qLBK4hLzgqzwOXSdVUo/3MIj
yMhh+Ln8UfE1hIpTflY70wOoj3N0Lfse52x6q1LOCGEt+HwpNLmUuQR0XRciGZda
6PyCqObswGLe3Pv5qFdi+XZi2O9RLq5Lw9xEBkkonDUqjW4JvHpE8OVGP6BTLJ6Y
hND/mkDu4l2NoChQG98rEF5uBChrp/8Zqy3e4QcBP98+Yp1CZFIaBntDCql9fY62
rmXZVHe8NJNotSMJQtD6vK48mNLCq+P95NWCJeduXoJLll91ya+yEyoO00a+vRQ4
D9Hd3QyoL+lRexFvU9VUOFOFyKmsMuvUbSExQYx6+XnUEw8cQmtJY0sxjnj5OkkB
JebCWgMAL/myOajN/pxBXQY4/ND4BXRSga+YSFDAFXHr4x6lvhYLJzrrmzpwdPQD
mywo1eqSZ0m3OPSPC8Q5srohRl15Z+nMMYRPZdt1ej6fCWiUky197xpXunYuZJ/y
Y0w5cYKcCyi9Q2pLfKyjx3vd3gQYvP9zKBc2AjtJiyK0lD6Ohvxoa4ylPq18zqUk
RKN31P8h1SX6wjz9v9YODigA5Jpy8sWYw+GCDYHO0Hd26ObTa1Sx41NIFOyDBlO0
kCxa7Q/1FV+MvIjvNXqF1uRQoNLAJDKZ1iFEvdiexcLoFeHdnLr64AwofLEAJLmB
87/e0mBtdITDjMeiuAK2kyLNXMX5I4iqT0HoMW5/QPZ8xZtWTvGdyX2mgd8f3vOe
KONxt1fqlqykOW+WUbjnpSZxjBlLUyCnegc7Mzg/swinIM7Ok5lN7rtD0tLbvIpZ
8uyvRSyqH3jbBdNvvI+Aa3sHr/UqNFfUk9OEk78IjjXUDk7Qe/DLQnt7txp4CCCN
a5/7+O6+EyKOOx4Li1PPSwrBz5YiI7hXDyHz8cGJlpYvp0BZDndjf27ep8aQimcd
sHAK0lvKs7oX+C7aotpV3vHMCNKY3aVfrYyDl+cgBH3poQGYMWPxaElD2HsehwoN
4WwwHfPcGtsP2/MNraB+4tRWVlhYIZXd2zff1r1DSSiUUzENyvwSkoql8DkEUTul
rS9qBG2/W1BvOS/6UnMJmhVbfNAAAaDboNTcZaGuCVRU3UW9xyT/7ukXt5uZoahG
wVb8Zm+TxJOwfFU0ATENJhpOSOuvXTUb5TsZM9LLSwGETMO6gEGF4yHYwEU4hE6O
HsJm+o/vPA+hqKw4mPCvkmA5h2+2ldUz3kFJVEoZvt1cyG5UzPPck4R0e5B1/aAD
dRTmAvfEnwOuTQVCKpd9nRzrgxeicAsf8iekzK3F7e3UV+cOQ+bRA3DHhFde4F50
RehiQ1O877JshfMAVPWZSRmOQhgkF42hao+510IGD2OvUod9sTfobSxwEOC93d/5
onT3V1pfc4cJHDX9Xo9IJnUsU6LZV0VTLvQMg+yEvtPwm3pjvmui5pL1zlgjDyqd
m6Tc5bquHrchY3DuyjwRliS5nFOJPpzP4wWf8YGrovNadQDuyMlZ8MDvXWBOOVoN
jQcT5z05CMO9h/HD5SZQ9fA2UNQJ07BieBIf611chn/Af8x/eGYzPDS1sNzr8SY+
K7MOTBJaABny2KPQf9n21HIQV2HzC03Gy51y3IS1uhvg04wq3sLXd9IOaDedkPKS
NP4pHKGbBFuouze5MlXAaNaixD5DEepVg7wwphZ/Fix/CLApp8FPi5B9A1b162XM
E+3QPwuyIG3vO3yjzV+SxlPbQBomVpgNr95RmIkdKQUbcMiWyN3687vFDhWusLJA
ECWQDMD1RMpzy1SKPCQM1eI7pvaBLPsd2kSHWO/99CC3ekU96+PuO9WQuVXhORqZ
BYN1loghbv9xkK9mZrLIngyzpqLt8+nAtAOfCvH6ty7nf7hzuhlL1Sil0izSFAwW
nO97PWGhPilpVtT1ayUypyi/2shPY5dbjhx65sDWRUXZQQUgaIx+BjLiLvrTJrk5
bfBEVpXJtd11uLYmqo9f+En2GqxCHenZ4ZMQd8mX8BPJ8+DHkLJbUi6vSqYq3dyK
WW1NF7Usbr8RnzruhpBhXUVM3glc2o2PaaVtJp/kT0uO3QB9JxwEfR6aqDPIYXuz
ghuTz2Gt2nWNJFti8Fp5ckxm+G9t/DBCAsknJy1ntPz9HXbPgZIRbG0g43kIq5Z3
vQQ5Bz8yDnuhwZ2wRkuV1EOy17LgneIse7GbeWRuMI4NMCBWrzK6c4xz/IyQkaDG
qnRXG4lEpN+DQ3zMyyWE7+wumGFOW5kJN04C5428DndQa2il5VcbA1BRo6G3Z5ZH
PRet2icFlcoMZJisiUXPe8wa12Y438Mlno3nsCihtYDoNk6YrGvx0NOswcmt0ejN
+tSmUaaq6gEnOB2bTGopPE467sJf2L0D5qDpROki5+zA0Y8IGjGh/NRlIG3st7zR
YpaUnmQi25KQPrd2QTKPi9uHTq7ErerDyb+JjOGV+9lxMrqfeAY+REcSJzi1/N82
QCwcwFIds0q/jfwcf14hHfBUbMdZfRqKkfAf7DwPJWfbaXavwNB3aXujeKxavGZm
VJk1VrG8wLGhW4Eti2/v53cFOXVZY74lcKoU7XJ7pyvRrBFfJ361erZp7OnaqBF4
v+/iqocGzr1qJ/KuXWwt1ig0yGX3YlAvU4/6VxiuA6YPg87p0krF3ayvVR5mBQFI
iqnmYDLiFrn/E7EE4Ml2Ya0ueJmsSqAGxHdhHPYOk9Z4/oW5bUK+vtYqgpTFWpGf
p1f+2AGdlUXG0jHMc/UwcMVGSvL0nIKAQOpfNymsu3KEDuLlCsBdxbJA5IXKAYZs
miLaM1mzQLBn6cF2MdQnJ7q5XoW8bzda8TG3B8TD6o2jKpKsbSMaxv8YdfWVURr0
DkTdbk7RLQECnBeUaySJfp+TpOWevi8ryBlpnFP1GEfB1sTybfoaGfuuxYrJkthj
UiJ/UMmbndKO7UuTU1lkm4KfhNHOloOjcCFAihcpgb00vS6PoFLTaKYpdirTbI2A
9sG3tDERsYLb2J370dU2VLalPVKXcYEXu7O6wH2PQ9wQxL1u6M9P4Na6M4A+BEj3
HWJdgs98GmJgoGgeVXTbQjCGSFCT/6hCG6wZWlvK2XBM04LZ7RIEdVRDAPtjtJNz
cXepn3f+0vaBcxn6lMwQuBWcqDc4OTBL/1sBk2qkNCjjzkoucVu9wAk6obb3BM90
p35dKVKTyYSBVTgqBgLOGbi5e2Ja8aNkjdag09Rkg7W6jykxmLeCdd4L9Aupdh0c
cWQTGyFR9872/d6JB4OMwQXjN0VbmsabceTBdAyOz/tuXk8lLaDIRELuDFp2B4/H
h7cWrVKlr4MnEnoFK6IjrXTJwN5WpT+ODzTkOczC+IF1nRnzW5rU0xE6ypwXWFIw
Thw2Ko16ipIhMldGs8mE7kfwgP+Evnjgn4TCnHXuzR/vbhz08atUUaB+OOBkZxmZ
pbZnpJE3xuEs0XzRUjhwF5z/9X2LE8hlSHBFHxhE9InALjI6EmlN9bHD78QQ202c
OHRlZZK/hyGbhpBxWoSjBCSt4PksmgmHstzyBuA6wGptEefeyqDHIz41F2MKkJTN
QiBJdTrlMkzVk1bQ7MAUn51sQRrrnk/kPjQkJsCMYwmBOaVkwyVoNgvNESgKEiQE
0nYTSysnr3DCrIUYKk54Y8ZykSOroTgf2SCT8UOcpomH2Ok/uluPL4FNmGEKs7mF
jgU2xk8NGxjJiY+PfpTm2a912p1OyvEfsaImdoBsus3UyMXbytBe3hPyOXpu0riF
DZC0CqX1mo/P10YU08sKaeM/5/ulPBCF5x9WUXI9fN9KdSYap8fjQU/lIkuhbzF9
s4UcfRasVxhq0+WqeWskAOht2AGVp7oFu7m8mfgoExiKcimm7p2TUn1PywTxuVlA
WbpVC2GAG+VVSjf/byBWRRhVexCRJ8xulwvFOAqiv11S9z2LpubbMhcTiHzre2I4
bwm9pAavvbYdZ1SGISO8cM66TtvolftDUSz/5gnNLN95SnLIg4UL3kN5r5yRDfh5
DJfYCLT19EKzJgaOXIIEyOQDrc8vsCT0QyrjtFDpTBZ+SDVaLjNM1PZE4tahzJyh
NT9My+d9aQklXrEHjeEXEQRkJLXTWS/a8Iz0afMENGj+Twzw9gSgU77GgyeBUCYk
z4ksalVG9TiZfesW3c66vE1rX3ePrl32X+eEx9hFiKaxOOMhP6qp94TAAZlo77HK
IrdlEh9+yfY1jsvjnQCsmFypJVs6CqpBWOyTA+XVDe4VF1pNN+6K+j76OPzwz75n
V7q0sANS/PXG0x742nY9dlECsGyBylKoSaWMv9XsSvTFelAJ4M8BOvEi6/1O7pC0
ipWsN9BCEWi/VM2iZJW6Jn/kLg7B5H/UKi37rGqpO53ZKBCm/qHRqZ8QFWcPnS58
QPUrm4kMdmDv+QN6wc0HWwcD0wFRELpJ0gVbjVgybCo7IgT8d8G2/fKUGZ5x7OCf
PyYFeHJ8WhNkjFIjuMvFMq2mabBs2RD1wR5o9DMHqfesI+HE+x3JsesBbqUXcOPo
1quBpeqEKC/f6qGOmDf20OMiTfEnXX/lYPRYyEjPs8/jNly+H1Wq2DPT8mrk3v4H
YVi+C/J3AJStO7aJVtwKvWaYX5Mbzec2yN9m9ShV+xsaO0EGCFXgMw5IjeE7o9Wf
Mw7PcwQNPAmtwb2S2rikQoJWVGipqbrGXgPHNWMqa8BwRvKAhgsETHTRXv6wi0rx
FYEWQZ1ni/tMRnCqJEM/shmXcmQN/Rp5vy7QuuRMVmB2XhXGVyACS5HrZTSmzQst
rkgpjwknOxAiIjAElScb9bzlEYd8BEHpuTwEF385ui8vFT6H4SzTOzetGxRkWVbw
h6wunc1b4bwGgfMYql7Fp+fG9m1lyCn67BweiZAAF1LEwi1hDTDWNr0Mt6WyuofT
jjGzjmzcWgt8iwKlXdqtW+dcq+R1F1A3eLtZGespflrQv2meDfCt1LOxVQNizhQ0
Kugz/MOTzvTxL9VeQ87metrm3i6z4V0ap2F7xOgh8lseJOBwV9qLuHSlXCn/SL2Y
Ra2a1EpVMpexighD2sbheuKZSsLTjcBtTHue7cKcA/mYeeKjDtJUlJmhWbt1jQGv
WWzntGDzdgxtBvVD/CwMoxsQCuKBKBaew56aJC9ETX3/Kb6OYtq3gj3KEas9NIc+
Cvob9uC/SEwSxqqKhBzR9gfWCT1DKcuYt3NcOYJBZsHZnmdHLEkXm8oXLaFmgCdR
m7Lyfoiw8Hd1NHC239ygMf/w7ZJaYiRE6wYJc50plZ7SXZcmHaTegozUhmw4PPYN
S9iJzR+H2FiTChPd3Ljq6zpfa1rvPDX17cd2an5sUVoioUMOyw4Dynh90ZYAADS0
miVWVub4sGUhbea7GxGlJc9ClUWrnQmZdA5D28gukmuCHVqR6RTQmsIWGPq9Ql1H
8FeIWBEZd9/CSuGWk8XN1XivK2zGhmRvS0983+EW8v0A7VycvdbAdAm4eMK8HQVq
JTO2+5hV9i/6ClRCVrznNGCEcM4do1DB/HMUqYog3UlrGd9BDVE4dMiRTtAm0aR8
z5DwHaP5ewyDXyFTfvmxmcYPt4wxr/fNQxVz4V1gbYmCo1mADe7Kwh21xsXe+XSP
xLNqp1mFhi8BwJM6PffRd5JQXJq22pu2n+WCoEne8gkwVYtcdM0agWG8Ug7t90yz
4spmzHyWtcE7m8x70sqB9uHJqtAXKw7gI01/zmRjg3E5JW9QVwVul51utvIuAR4b
iTO7JyEIUn/udHyb+LSLoIAOwwmkPPqL/tvMjuw18kY3YEpKHWwtMf6ZUj2rXg4d
zXOtxVy5Obe1MRj98RFCVKJdFIc27ITyzLu2vat4PKYQQMrpkkDmN3Cz8cLnBG+D
GjziOsAfV7HJ6HP6xdez5ff01ibibOVQLOxt3F+dXufXf/kjticUbqlyXTRFcuhA
gIgA3rYyolTCMkqeP0/jB5ra0RGKvRN8nL0ObrfbuyZ0CwlrfkfYmhjDxMbAYXeb
84Px1ak341jvrYWYpTezTYTFuh69MTRG/LyQ3wAoMM4UuJjAolXECRIj35XJYaUt
vrE/EayfSZpr+YVtw0sczcnOdYjXAQqZDhpP3ZKEpLR9e+/4CwrIpahPp3dycE1I
1t1jh+Rbp/f9MC8AaX8fKgoQx3dB9F3Bhy36NauyokDKuLYeQ4zxI/aRre3ER1Vn
5KfD1pb1zHBRJhIZMr1FF5TPFD2svcDDvda2wrs/FBN1ADhXvGcesIPsalwQTk0L
x8VycqRKEqhpaMMkAgXfLbHcKLDQtGG104ftAy+HzjicLuZr0B1cKNKPKgt+PW/y
ylhEbShYEKp7mOXdiu9+oXK5GgdjIAQZqtjtQHBB5tybYnpWFIq4eW+X1t06Inmc
fGacpGHTpo/8mXTSQ1btwsFz/JCeaYQXYiITpEvMZ1NBw4+Uv+5GW5Ke45B7RT4b
LlXNdzlK981yDA1Tb5Cq6zU+gQVyq0GN/1frJWkDazQR50VWKYOrx26113O7rlXk
oGHVFkRwLco/CUb0NX7EpB2Eh8Tkulq74UhJuuQ4drnnw+7G4g6v0/HfHe7/E4q2
WnAk8nFb2VnYp/rqm7HnQNIVgPOwY4uAlz1gp/KW51+1sfbmVWBJYU7PajSG3bgq
LU14cqgJ7v5S78lQqjiqJri7S7VyvmXuiqs5JMlrk1EQC1B1RWuWlJBFu93h4nkw
x1NAn2ga2ffbBGKBpOZ/pwDF9AlosMXkNcmDdSrT7gETuYyq3GfL62CcdEPDiAuy
inK1a1DJf7MQrduLsGxSqAeMvBcIVGWCLliou+g1Nkxu1YE24RyQ5QBxEY5iL+xa
uZfOEfnfer0ZIN+f1C6M+oXnWGg/U9K3o4kkHCejI7jbK630vpHHJqBw7bvCGUS6
Oax50Z1IZE5dVv6FemSqCtTPNq38MezXSezvvWxY72O4gUjG9vzgHZ4Kv2H607ZH
Zh690vjIOGcQ3RY7EelpySwGuu3+IywjtDV6Fny/IRzpJ5pNTtdX6b8Rl0u+C8X5
TTcEntdi6VtTAcmrfMZ+kTo59mjnAaKWf717wmSmnvJqIWubX0kmzcb4u+7FPLhK
/Zc6bPowi/5cUv0AbjCc8iXwnxHCWBy10Vu0BNVfT+9k34xvir2wD2JKDpvYtefi
mYJNvCG7YKds+h+d0IikrC6TM4G79/VmYabUSUB6K+Gmj+n6WZJ4JxnDXMbC2cEp
kMkC6p/hNvRBeHMvJiVlS5XrAOLo0kadDMWWWSLC328yS+vfTaxGY0NVqp3QgR/v
97/Ot7YTxwq3UDRbRoyF3ePO/828ek5w0RQQeHNrSClmIP9J2TdUKIEj/R2qGffQ
JCnFyqHGTVrO2LVKdRTj0Zl947hsZpxWLc3yG41XZXNmRHVMKGbjg8t1LdNw54SB
a6TJyWD+HaCxbJ/Kl6NPEORoy0NeaZVC64BDqSu3pJX7ZPVAoCQxpstHjvKaafiq
6rAA4HjNTuKC55a8lPNECUNlK577mGx1g7vYeZpAZTDzgwkf8gFJjLj6CEfWxNYV
raYWEadeC9IJJUFVLK/joKqnYH+4b9zE9SkQmxWf45eyWonSgyc/urGrAteEFWiC
atr0fDFxzb8Rn/bmhqQcHuCrUEz62fhuwHfFL9apkZUUlFSITtMIrKDnnoWNzf6o
r2uUygNiwx+azpf5uvTJKUtGmt6rQ7CAeAlaj83qtMBupbR92Hvlsby7OgRnqFCn
Sz6jX9VoZITXd50vi7Nj0CDYYuTHYbl9FZIRxiiLA8Eij0Xj5Ej87bLkPyIY9QSS
2XorSoDNtpX9EZoFbx5Rmr8D66dxrBi+xpHKToDSScDxIIZp+8rniPjjw/xTh7eI
Ol1pSldusph/6DRokLg8yVs8lIGRepfchZkvHYSjnnu6e9g3gwXTFgFSboeBA96n
2jecB6L9HdkX0j7xwopg4KiUZqClHrrHVVExqkU4lmd2aXcjb6lOZol0b7Fr/MTa
mJBEhaUFY0thoxr76PTI3lt41kCPmnqXN8b/qTuo0wc2kF6pXvKjlz+7ZrNg4Zv4
UxchGrIN0rJbMRj+GFjl8nszCOROGIMHCBMWfkboNdsoRdIEwKRNEksKHeJnjuBz
fzqMeVmXm9Yv80oyokVloCLX5N3wonCnPgtb4qXy+2QpPOecKBpAK0GIz+O58P0k
9E78reTWfZGksIOmDHKNc1aa18TQZtYdO/U0wGYCeUlKTz9eVnZNsf1vWf0Jme0c
cMjrbhX428PHg3WyY9p3O8I5mgCCN30zXmCFvDZ7Zlo8FwonVJrR9u/lufIzzwb4
niYMmFFZqqKJTxqXUO1UlY7Jruboa24I01iti3tWDfCJ/stesQlKfHpHek9f+Eb1
QAEaVbWQxgYKciW+7sP4H7JQ0Qg58fI4nufIlcBd3jSJm1NXNnj9a2+02lQ/jbCD
lRzB+nuUsCijO0WsMTMjk8joMeFS/mI8DG51H6IfE1wZfGNHv+9UP8g2FgSLPM8e
qvnulCQfOgkgetT8y3U/1vYki2Q+iE6dLoHaPbhFLp5m9ahDlHXZnsTqwZwO0Cz8
hsJPoqTGRPg30PwIMA79sOfyIvV5zUExAJBh+VfyMRDBVv0t+88Bf+5Ync40gtB0
bl0/rW2X+jqVrz3zS44AvjNS4R5NGtPxYJs6RnTm8h3ND7rpSh8e2YjzQKnyfQD1
qQgJJfBTyOWCBi7WQBzfbX7pfAPRLpTBi4pg88oFRBt/iwAAXZHBAI9rJkSOnpkV
PM+6gfWWNiX9YtLhAhYhq4nN9cdEvnQX5g7oyc1VnH34LQ7DFd1pWLiUtDP56iy9
9n4GrRQP9wPjZvhbed8V/FAUbclc1QPJI7kb/ocA6XWPuP/Fi1NpKcP0A24+xH5t
XgfW33XTvzU63Glm7HHRm68aXiAq4+4Rv4s5C5oyO43yuzzpLVcP1/a33+148Bxo
D+jjxOCFMyrULkGuqAm/RLGbUN13L2IcGSrbwoariU9xYEvzyb3ytLvuZDV//cDg
8V2xex/4E5seNsbR8CvP/v377y0GIM9pUELrE/qHbZcwTBcBnn2gRLPjRu4PV9OM
FpN0wYyG1u7ukEbmEPLqKUxGb+Shl3OsgYRm3nGDt+CaZiY6LkI8y+RVN5tjOReZ
HrSow5PcZ6868ul3JlkjRTbVwMu7Ml/tTmGybhUce1LV1RlY2dSJ9jCUM/k3oM8p
FawFIV/9gnNnKYgJwGvE9KVHleamtMT/oxi0IZRvhRpSi7GFA1D5dR63n6h0YHCy
uwiOcMtXdPbBPGRgSXZzVzn9M5z6pdzGgpPYOkbYuP1h21pH/di3EONj1JO/psrp
ok8gDnRu0i5S9z1k3rXpHcvlW2P7nUQln2ikVsQVpf4BQYVaEqiB05Q2RjLRzESu
Zns/N1BblyyusrhqfL7st8cNpo9RWBoos+aJkArTBeOe4EiJ0MQEh9Q/Rxu4BkGZ
YpSN1jymXqpsrYjKfJ0PqkoqQdl40//fPdfMpw9omSfwm2rh14cbTswmltaY+Bui
ZIniETeglGANhTWa2529Y2bCi4htqASfnUNdwOAdHKGlKterjesszDhjdsOpCIVR
hFDRWK02UqM7wvuVljGy01GRbxPJhNAwT/XHLGXqdHTUzwSPG9Sl8DqMKR21/qFh
oOwrji3P4tqT4MVXpgYPH6Csj2R6HQ8tFPbPVG4OcX+KB8uDwQ7gMc2NrG4qpQU7
3fQqcrTIOgw4J8QpmFiGBR+Zl/a9kB7bOPypyHVnG4WU+uUwIEZlR51upasB3K99
6kTSwrvIbWJVS/MOfAEhNnHKrSCFBLC8El50v/HsbXxikG5WnKAWEu0Ixg/S0EVg
2r0cuK73Y00Y+cv0p7BDVG78ZbbUsiC/qGtJ7tyJOf+AlAD2Ewcmfx8uu3JTgNa8
KBMe3JCv/CRVrn/9aAO+QbXNUbzedQ6Ye6Z6k5zYGpc5MuF75CvxnL7tEwwiqT7u
vdI2FnEgnUB/VX4zo8wPxMmAQBNB4fwohG5pv8oqLLGe44YpHZPzD/aBI3GVJHN0
490mPnPX/OdZ/top10uckXw+nHFTk0hkmsbKApDqN+kdd1nciLPgEdZ7R5SW1udQ
5Vsi2i++QbxYTjm3Db4i5GFBipLYhZ8yHEsWW5LO1bsypdz51QZC+SS5rLnywH4d
O0byEiJM2lbFD6ktjrMeuNHQskYvcs5R26D8aNwvqie1xLDBMc/yO1oXoczAewMw
ITRt8oZJlqK+Lomfv8GGVza5Mtnd4laTeu16/vp7+SKIC+sbIEGXG3/SYhFru2tS
sNWB9kJ/lqx+ORXNVzM8sDqtftyjM6WyzflPaO+yb1hPpxAWv6vlONm3M6/UaSSF
1WH92DqN7GqfXCPidpDMX7VH+uWStG8S2nfPmsFeAdSASmtAc04l0iN63S1Sno/3
WN9U5FPkf23iJBcQXJ6lRaR8JAZOGVg4sPUUnszkYk5wEkAR1ZOkcttApcyenYHb
BVWPEx4VPq0PgLrWVb6vR2M3JJjvD3jZJGTvbLP6YBuuOkpemG6zj36gZBgQd+oy
GI9DV7wr5CRYf+2iYa1ZfMzuKvq/wQ67Z+BloxPfIHO1bKtDuNp3a3xHC+Y3mj6R
RisSVbJokfd+MqMBXSCMAaD6D90yCojlKR/5/zSdUTHVvr8MfIkeDDGqZEIkQr/t
8WJOn+Hv8TWpI7++bluVSr7K2BKdhzVrJeFXMNiDPlk29ntRfR8OibSIqrxxEO+d
zsvX1lDvXCSlyqkPIdw2xUQbdgJ55UtBRgFyBsVRaZAHWaBOh2nw48A3FPmlDVUe
sHM0dpAQrXIEK3+VLas3Wj89AVE6k8MkEFtrckeAzL5ywUvdlkgBClLu3ePWvweh
cJWc6HiywCdggHM3JwM0l1SqT0ptCJsCFHDRWvXn8DEpuchZwHZh2xZKJp6VD2eE
HxU91egojV4KLEPjj0uMA0ezwsuNTauToTfswodvmN8jrfKSTs3RYYpTcl1py4gR
d+e4i/ypP63OoGXZOyS7lMycqlj19g+sjMmQsZ0zxX5DziQmjjBZnLH/jXpjFAKR
OkBG7Z4n1ZAjj4cc/8kPnxkIxoitodaRif6nf8Nokgzlt0zOfj3X/1tm7f0XEycF
c5cKdTBU//GBCpXxX4qWPlRKRTNBBSLhmYLZLO+kJsWdDzbMU+Etk+e8ZKik+k29
zWnZAmC6JQtN61t0ytbLRal8zI5+OS02HQwRZMmra1+AobXIItfxTGUI79z+SB08
uNR5Ce0T60/ElbtBKlsU8A2bvst0gjYQm9CIhNkxpf6FOmRpg18CVOwqlizYSOEn
OXLL/vZZqNuKdykF9E2GFTk9965OqaHyHvrFj0esoMp133Waq4DhciNHxBLTfld1
KXu9MfGhgoUotIunB/aDwDj0N60YmZeT8RqG1g17Ymgace8Pj6JhKjChY8Z+pacE
YFPIKPxTquj5bySjBTtckfLnasJBCICKrZG5dzudMYb4yPQycfC6V2U5iqO9YC7U
6NIG/B2PXn+osCi6SlCNNKR2FIEgjB7LSfkmWvoR1zSJL+mJk9EPJKc/YTBXxG+F
2S0rueGm+DntZ/ZfYPlwOk4Mi9zhiyiwEZymn7CY7tZLEKMR4cABEaHvaeWqOQch
JCETbtddPLBjDNNAuAw0BXPhzKrq3aRaBuVVHAJrMazUdI+elsyeH/vjrZWlZzFo
vhPOGZ5Tl9x2EsiOWWYsyKEvQf+mxPX4oW93bQFhPxz5/2lQN6/+lTZLEdTHw2ZZ
Ego4WYyUfG/dfLtTVhdRRNAe5AOizfcVZlQcY1JQUPRWVPADHSMJvlsN9q5XCQEC
Kkkd5xapfNw+HFGx1CVRFPZauLjztpAs/Z7r/K7j+rX3oXZUcKLK6MhDmff5xVki
kNyKC4Q/mDQd+vyoFw0MJTqbSTNLskHj4X3A4VXdfuoOUhYXLqJMk3KZcSWcJdOA
llqgvsKqNHEIAAMpaWVoaXNoVnU48PCCJAZRKOnbo0pA2lXLnD6njK84s8SFiLZz
XpM2jAa0N5C+83g8pF/AIcw4nu882CLzhhG6ElO4NT2Nc4NnMUF1dpcxtbSHDThn
UEjCECq/9+fKcoJ9afYQbC9JIIPTuuu3qOhxRFrN4HApIVgpiphhmhpy76g5SjGW
uK29B6tCfnpW2GgIZz9zyidb3xzhJATDHbkLjJ32okEnnZYZcpExIfqaIiWyZG0k
iDRFetpONceVJQqO8BwiAkvjIfMIwNOvWwNJDUPYSTVWaS4i46XRJ7THvBOPfghu
luvAIRxcm/IxJw258LzW5YF84o9S9sZIM5ib0IaSlQl8JuQdL9e91NxSL0ePnlCy
6SQrdQZ0L/oyJbFMWZ3GSgRKt/4BD1TSQ4gtU8Do3R0H+VYmnpQTBrLld+F2HiYI
Aoa47vZq4Two0yME9QQRmxDNWwDtA0+TTdxdfW2A7YnUp29KrZIDXrr4p7G3zl2t
apo9LKHd8ErJkhm10mkYqKw02fThYrPeivvKbCNW7bp1u+B+mDoB8RkIrw4j/WSz
kI4KXc+6OWqq/OSsXAAu7iQXQ/Qq0AQy3rIxeVnmrcbo/YCv8Q3oJfb9cdZHgBR4
u/HMLIgBFkM/I+cjA1xxxWpkwfxqGq+79B4+iCW7WSs7bQWoSoZQZ2hWwNdPJADp
4YmDpV+mzO2pvqvM/Ts5zQUUg9RwLBMkUt4SonYNOdYBi4cYU/fQ9G/pLa3ekgJ+
LFTd/ciwzerkqxa62RwI0HxnS4Nl+SGVcafZInlqIGdEh+8iE4uoRh9mcCp+iS9L
ImL1Tll7Vk+xjC986uQO3TgmJ7vcj5amn4hZsHBcFK88V4Sgkf4dOOoge0sBLqXW
5aA+2ed0YgboQVvzHW85YHaSwigu2krvwWV/n5Ggqxqs5siAUB98G/9vxWzMmlGI
qgo+eQtadDgkyw4GpPaMKd1okOzR5GK8beZmFjq2eYY5kORJnoQwgX12PG7i4UYA
1pIppCozJs7feKHPHQKzVt8Rs90qyq7ied5D6I5l46eyfeQWFffY8EjpaO5L3mrn
STOXgwqu6HimttjI33EmDx6tJsPNtbjfT9sH+pxELvVuOrLnpBXFs33lYK+vdPK5
RK7JaXed3lcWX2F0/js2NhpS2bHvw2xD/pkLrY1TZT6LAs3P0RDcuLrXE2l3Uggy
VkIWzCH5P8/pUVrs8I+v27q5ct/fnuLOhg/tjGnaRUNYMT23IFitB4cYg3g1U933
HDoUFCYJifyM/PAioGQTf9ZXuHpi+qx8OwFddB28YJ4VTWl+Y+/j60e1pf8vP95f
iINxsqPv6djeA8P3CnyGMZEECMAsNVJyMMBwGIzmq6v85lO6qzOgU0FXC/a74WZy
FJkOS8sKjSGn1mu4fEJZImSdmD8tuVhNcvDf2QxWAVFpUHXO32ZtONHrJvn+EDTa
W0YuNKazsXtOAhpdrVJb+0unpYbPg6uod9xaiRwwdavb9+d7eRBe3Fj1IqdRVYAQ
bwBveZhYq9ebqoNtSN0LO08P03NwloqSKdwTURG3N1nfodnGRsLwWb5OoT0yciA+
b9H0GNvWhrTUChvD8XXqXU4oZ/yzU3hVMP2MReVE9lvcrRnGbuhelDJNRTrOkkP/
qIaUJYEjggpRgh6x0bmU+sMSOH5QevDwQHQk/T4231I1saHpnoVAnCxV+LZ1+YV4
VNoP0CV1bG1b7EB0YsxCNNiPSSlz4VgKTspkbPHkT/5GnaBVTWDXJarHkMTEHi5x
Ht4imNXY3MpgvhFnb50YtExL7+/N+EgJk8f9XHxutrhVs33+LKxMJ6kBNM9+JSqY
+OJjAQDXG5fiWR/i9UKYMeJtGX6YUqcFyQUL0IHzDR2nna8xzO+gOmtcnQ5+R9LQ
wiSt6PLGZ+YDsFSE1+2266nIRUflCr/F04IHibUmmhaO4uhm4rpvHc52tNEmSwDV
HGjNGiqI9AzED/Mc/fm7/QvOI7rpV3mTKsz/3rezyTHAU+/Wqdk5s0Xp58dbqhQE
fJYJFTSrdAqkEAPjQ2FwEFPszFlvC5QSW1j7dUhU8BuQBNAWv1svNoB4tX/UvjfI
7Els5yP2+kkBWdToOYhFaoombIS1WwlkiHYHPAOuDIfcUjgcj7bwRL8OEOJAOh2B
bJNNdpvUyPGsg4MX7sOMO9/7ZWbPedLb+wWjTL/Do6XqD5YArQvsFFbHh0d0Evr8
lb/gj6n/cVHcRKukVxC9oSVVpP+r5OvCX6jfXsAQvPwZ8umWDKIM7nqk1PxQ0kkA
xY1maD4kOVI3M+ULduxz9MF0lAWp7VxZHRp9IIEU9CgbIss2AeFXwSyzrM8FC5Ag
9hABk7lB61M0oyJPMs5ywICR4o8mFmfxgjhy5GTVfhYqI5osCVumdc1V4bn1tF7l
uSHfwSmlbBwxxzU+O7JuiVWG7a6AOSsgTwBkIyfdbIwdymF47BBY5HsYndBLzps3
xMOXwQNvfwIJHmmsoKKwXFSj4bBQDQJE19OAGUSNUo+L0UUqhK3uofjPVASU38lm
UPEAaPKADXiLTfU7sl2kgOX1DDvKC3PUoq9HTm6NAWzNo88MQ3l0gp7srlCgE5l/
P7RcwGIyEc/JpXiNadfc4YSrYIKN4CQEvhx2Ot9u5sdfA1Jibcnvsd3kgd3UX9Xg
V+AF2cJTzVe2Cz0nRGdHNmCHc2Lcn+AUiVBk1QqROZU1Wsziy4CQGx+G4hu3/qkz
FI1YlL0l+ZNYwR+KHiGyny4t61N/TMcjEhTm+JWcPgAwJRLsBYkYhMV1cTJTUYLN
umAaxpIW8Srg3oW7lZ5fUEOn4fE2aZUiNDnOSIMEjMqEKVUUQzyEeZ9h3/ODgtzl
3Nl6K8+yciZJNDF1zGkLslSXUJuoOgyZoxlqMeTJlX6TktOSuoV1c4KV0TWc0iej
mubvmjIzq8JtSUFVRLT2hd+UXUCfxkrAQo9xtB0bWzn4qOCeI3N7XEjmzdI8XHdi
/zjRZuPXZ74mKIvoFTsEBGNfk3XTKZL9GPGn+roiVVo9VkzFAlEpuUtV6X/WhrGo
VQvdftY6oRd06/Xof3EAyjU4w3oDraH0j3MOQfHqeRbetORumGzZxcrkevWs6y3g
71xTu798CkTNtxw0WHzK/82mF+rEyoh1GTbg5YL+linVDB8HloPZxHuP6vgZE7Gl
O+rMCUtKOL3uzDiWOKtEvup+yw7jlfuX/M1SSfPc7VdvJetzgEpkWKRdcueDUecd
1Wqz5SSaTm+Rc1gUXYQUgUknW0ma5QI6YD8qAgNfmWQmZ0UBiSGfWTmHQBWXWZb8
4Waior5kbPMbW/hcNkJ1YOaxyjM/HmH8t7O8HO2HTppkBm/g3bxA78qsvwR/wWkI
EpfnwOSUm6NRVPSaJF/VfbY5nUO1WlCcoA2QR4RU/YfEggECGz2N7cgOdlCB5LXh
wurKMhFXgo9YjkNao5VtHjtfFk3mGGz9aTc8T9V4IeBoRufY1+CtH+5XV4TVjFUt
PFr2T4YNM6q9rtzmLmDI7s9vC6D1AofKmGBbPmYa10dLKPTVaokL52Rr9YKkthrX
UpaQEpMVBpRDTvUhUu5B7A4SLzb1kv0Vcz+a4BNimopi8/vBvmwTZDMBEBK5Xo2p
LhYrmsyht+N0AIvv0rKMRP/0I0RaEwnRyY08NvXSW9Ph5gKtwk2PDw3RGIYmn7eQ
H0akVtf7+SREEPDTIN8llaXQNNR6bRzm40xSpGzDkHrrvtsFRjxMBd2M5rxcPehI
Y/FGoezez9jdPjYv5QL07TpLxYL+LOBB4rEfLrzywXmqyUGzMc9luMtO1FBXjeFk
34qJQHhd0NcGmBaHMLGfzkiQxu77+FDW29ieK0CMSqIoymtr1fTuXPERYed+GxkA
EHgHcrABN9LuBuCty/LQnB1NcEOE7qg5bK+Gn+LAQ3aNHfawgWR6CUpWInHD81ll
r6Ud8JWoj+7/G4CWItnqVohnMnTRSQH5sIaPVxNQFbq9MbDl6gpIbMwWxPWkdHGc
8YzOjSqdWA9YDqN+VLW9GynAvq62gouUyT06vuK5XF7ZdnojPdwCp4sCscshzdrA
98JUEFqdCTe3SH6JKz4ueB6xVrITKD7o19LkPUL8dSA3Ekx3jyeaHvr/y40uKKr2
tJPGAwxXB0SnCBoaNZ9jkwIT8/yHptmY6UbIq870QymviemFNRIqmkSsfDjRlEIJ
1JNfNv7A4b4JRXHhRPNeX+fIb5ibnVWqZcaiOSom2y3NtJGLkKmO3lp90GcUWUrU
XuQx8TDDG/luSZ2+k9IISKn2YzPN/JOFXpycfua/Qfi053uRye013+Qwc4uPBo9M
M0Eptti8idxpBoAnu0HNISQsGUkco7SmE5+JpqxMHs891ricubMUbCeqx4LvxlWM
VjXlT7SGslrDPHyoMUxUvuq4Y+BSe7xfP/tVS8uj9LhDCBtfV2eR+JpVfflV4IUJ
UTZi7kYUEX7h3kF2kfw9tVo2hof05xrmt1A3bpjTvStG0T8/Ro6zTnSJwQQVd+xD
8SyKE0cX7Aqm+cl+52fnb/rIDKY9XEI7FEyWwIS3eEKfVu3QdpaOc9zGGS2M7875
2N+yZ6NTiHGsFwWOjeGhPtASaeDsK1CS74RGLhsIxd3VVD65VyLJUZes1tzwxjru
qVfai+JhDJNWM7sFvoOZtfVMQfkf1ABsFBDqXhdg7Zf/IluP/YUNGUIfepLLcTfN
eEJt0EWI5baAsZhO2hddKnkALaR2aOw+Q/Ayoqze28v9mdaauW5IEIgrdII8ayDD
jMoKM49gcOg9/gmmrq9H4mnVbOPfJIWwgsLnbh1zFcAK/4OKQ4/c9Rzd2DriC8zb
+MOAVK4QlguQx5crR2ODXO4rM2eVzsJ8QMIoCyZpqxqgY3G7MHOLXmsUUQWlZQrS
DK+KwYd/k+gGRyjrp+USrPeHUkwh1m4Ni5UH3a9/oDsLEV6hUqjkG/STYjyg2G2U
DiH5t27b9dQqcDf7Kz9vETCfPc2nt9naJFWHPRZf7aJQrT5ZhUU5muLyeOXTj48F
sT4mTeJWX5DzezNua425ObrjfY6GGT4Ap2lbPHj4Ig0XqJbJx0dNHG76jujnjpdD
hSjK7icCyz6R5zhqUQsLNpH/fCT+Lvq4++VC9E8DWtx+AhO0C2xmhj5/DlAJP7BT
VVE9WhG8Wq3I77IJkCP3NTV+pHhr1GQXEpNi/EIGaftSvcEUMiXuWoAzsZny98fb
omMYvgixUa4G9IBx7istZQeGFxOZMt6HP6YTF5mEbWGyUQGLRa8tlBeCmNdmECBC
CKFcZILK17tcSKKIeFqP+fhBIeR89bGAgqvZpsehop7S4z+SznJs0Xemxga5+89e
lCbfw+KKeXJWRMDiaZdgsZy3C0a+4lvxSISNXHQXQ4YlEmJkm9yF74/fR3hxew/M
zjNOVfE8DZnfAcakMGpZCg9vIuvQKXAYiVjPkWQnwm69fhsgpnOGy9aFAlV4PTnH
wijcAIdJs6Kz7CoT36VR/rdimaNCkZM0tK85tag7AHidd7GuXfHSs8+gygbyWFPH
p6Nkq6k6AnDyTpE1BlVAuKY0SbQXTjqyYnZUK/rynpZzQFJN0+UJivJ0Y+F1qo+F
yXcha9i8ob8EaDfW5RRAfUywyIeWi2lLgsYyPFxo9XFlscyZAKghaCeS9OvkHHhq
t8WhXeN8lovI1TTT9ZAKBsx5paBN4I13laF4MXA1leXF3Ph7P+yF0iW+LOT+kQ4g
G1/UjNtQFiheiWFn+ByV448vcD2QhPAJfAKnlOzj91jMLMTevmhU740c+6Q+VL6d
bSSZSoD3K+weP6BKjyRcZhZMdqazgf+ldqz6K10l9eowqGdwPpFsXhW0XQ1+KrcL
F7lkif2zrOmVm1g/PpR7RTH4lO+0YW6vCk6VbeRjLP3XN2LLI6qwab2ZhMNWcZbb
qKonQCiGca5yFrrvDjsalxXfRsiehE6UaF3yI4HfDAAgkIP7RX7wMT4UrM26nLum
Vc0PgEDYF7ptnHDixyxOn5cyTfj5g4BOyASxareE9pOoOrXl9vuA4D3M8AOn3JVI
QkWTWNCchU90RFwPZtiBwl4+MWLIeBKR0bbfJhjYUl7ifP2MJSCPBOeYEtMAZY7R
cLnBljshYWdg4kvBcdc9LXtGEQH3j24NPTSVlLce8V7K0FxTOCxkdWbz4kFsMuwA
UpaOiYDT8PP6aABODIhENj45bhFDgWx52Zk//orfZBH5QiDf8iWc4oTt0dJAnBz+
QcyTqKi68TQg/4GYUeb255NgBEtMs23506kWp+RmTtWhzi7miprE/omNV3PjHhpg
G14garGGxMqmwi4GkFdfkVvaRdkZ/o4H9sWywJuxnkVfMdzKVe3r6mXGZ/mOtpm9
eaTorRAR1Bg0GI1BTdJvO1HsLsHB5sxQirIvDiqJxOqmSjQLrolaGkCKPcqZpm7J
fFE0xE0bDSWkKP2gzwvLs623Q10inCWMZXb5SKY64dvys1IT9jWhZARB0woTWtXn
XkAo3JZKyUcg7vgg14RnBfJsGssR0SehTAyh7OSpJPPOk/42LVWXyqnj7N/zpF7L
NmjgS9BnlzwNzSsJRnaBdHWLerYRe5iPruAJzN56Kiohb3rY/grHjyallvhYN6Rz
RayEXfjJ1pDLHkC1ZIKjgIVJRq0M167zaX55NgGPJpAS0WdySBnNbSkndejaCa5E
Qb7zbVzSqlrWuLIFkSgR5qHe17TboAfVzmUnG9yik7LdnnkoNgs6hvgXIGa1qSC3
WUcXstE4q9okgdjtfNLhWJJksiwPpgzJnvm1b+qpNRmbRNTG945mkMAtk0l8X003
Qm8+DjkgMsbyStK1CIqiIUa2SGnGVNg18xlDTwcOs1v+54qNCLK5R+P8izb0Tc63
cok8t9muSuhYQnwXd7H6YvN5upWJKPSL5V51ZWEii9j/ltJeRaVxy6umfj/+AsqR
yf2sXUhQ9QdM7WYfVkmRa1AjefCMrlD6rEWF4EWW+pwj+d0dmbmgHnRhPhX8B24j
Rm5pEiMhh2A0GONoOgRl/KXFMQsZxOH8kiawesPVz17zQo1i8EUd9qmWjPloU+EV
+J3medVNuCYB086tF8T8CPjyoF9tceueiXWq6NSnuLywYoNFPHA9vHxm9Mykqf8V
kz4LG7CMngW11JzbO0Z+YXQTZNJ3orjLA+WyHlyiF2R/HocYEwRMFYj58TyrMbfN
UAEwS9Y5ay1tZICjBohCWUDye7ulKoOH4NwrNzLVTyM1O17rmTgcAmZATg4x3d5w
wrxCqgtfcv1n6/VM5RTcmhjm2+jbnC60v02a9viAKDbPhIrqLIUdWKgpneQyBm3n
QKsQ/My9oWbWJ55Iyk8ydTjz9w7/j6bceuCV/VGWDSzLLg5167lhGr87mB1p/DN9
8R/6SpGQ8c7IgU+Ill5SB6sTtHVVDON+lxR54gl0ylMj6JCu1CNbTjnKoxcoNvHP
jGWjgmEV2dNXJw5S4QSUCeNMUiwVbnk9SUHV1IrwILKoOjNRt4Qv6dwNT3JBufvS
2B8P4NUPvjD6AKE4RyZSdXLP4rFJKE/KeukjFrKk5dQRzbRANWpI0LEhZD7c4v/n
xFY6F4z++XzhMpPBDR3+dzVdixAeJcjMi5lpW/yfLnkKU7nEaNHtHd/ME6BQs+4H
LwjMCQFiP5m6HnXcBt56s9aKBFiLXBmBpAAeZWCqqh65kyL4HED3qoJpATHlLeJX
sDOvqvuGmbwQiU6CRHvkzDzW527sv2vD8wYmSv5KwnYztUJh8Bn9u/Us8+tBiI2F
hZfyuMA0d6C5QwGW6Nmy8F9Q+BPoTpjcceS/Xy7v58ub0/IqlLNuH+z1Oo9r97hY
n6peJuOZlYP6OKF2NyHikcKPjI0QkRYdti9ilCqL/PdjEHVP+eFsn8t2onsfHJjn
eAxOnSmfGA1Kq7lnOLbJtn25th2W2UYJMTXvwoVOQ3kzminSJMvdcTPI02lHNZrb
0vO9L4ErTH6JCmvdfUPwdWcRRsBz+pe+T088jOCdAUTmgf+JqAX0j5tJ5MnDvjXF
2YP52qCWZRop/utL6W5hlvp9QiLUtUL6nFEDwF/I5rVnn7AlNPRz8u66iCWCS68z
ZXiyaAWA18hJo5/mubgn2ZJ2pJcFFtvlToqIQkb0FlbF1qVbBSwm5uKbT81kjQf2
Enrd/HxIlNGeQXh7gDZb0P87dGjekNUPlRakDFOiL4K4u9/UvuzA5y8LeNTdHcjo
p7FD1I9EWRkoY33YL5oxzYa3+8TsBLY2BZ1Y+A29sFI/IMdrDgIjPUO4O+m9oVTv
JkShy4to0BfSe3RNa1C+QzO1xd7SsjhTgXiA4rf+HhbwJXiE0MQWf+ewtF1ZuFO3
h4JkWctRm+x85Gn7jjSBRRW82jN9EidVvGbKCoGekk6IVDbFw3MGEIAk9iifL03C
VLIkWtzv5HTN4cjbm1Rv7J5zpF/him5iRYkepU6V5WsCuWqcnh+MFo9i0/5Y00ho
qH2u5k4SCSAnxrbQsLKb+6vA/s2U9F0mWUeUaunKxZy8khB/DcUGdxRmx3EHMBCM
MISVKjLEIXBhp0SNb3mhKq0YoMUiCJVRNtigRqa65LGQ/7XNR3BOm5UB22byjyk4
JszJC6KKtL25JV1lBcbUEBljeBD3J1x33E5HbnSHTH7x7iyhUyBEAAlfmbE0HYen
L79p1NSdWQwaFWQim3Ctr0+FZSWWZggEHTXX58BNcMhlOGqIGNhKPx1X2Ynr2TKS
d905jg8kz807jqdTbGO3smnGXEnE0K0B18I0C0DTxlP/8PobPE8RveNagAFIna3n
tOrjfKY6FJ2NgyN1NzPCiIZCUm67IjQ9Mr7HogtiB4eo3G63oNy0MeJhFkB6GErt
XPIasR82WqVwSj3W+zVQLlCC+9D63TwVZHvhoT2PC4nsQXIPaBz5M/dWsiu15Hb0
gN/iDFjwse1jMFni5qnlSNdc+yW0m5AzzYR/13X2ESDpqHHRr3wzmx+/glbrzGaL
WOQME7UTdgRtTFNIK1NVowourPzPhQr1El5h0UmZ3qXlEFneKGCM938nhgeEd7k2
OF/Lvn9gUPGcdCH0OaGdFO2SQwb8BM0zSRGxkL8OfrHOAlcp7KFHHFzANhkzoVmi
eJR1Iz9FRQQxDFAHttPTA9gnmDwmEqYHdY1gc6xCwWoTjj+ElnjbC9pavfjMF9X5
m/oQSy1nUuxrosUP3IPXtkACAIG2SoPcuvP3F0Cj6cWzJX0/jFea/FxC+4zANRyv
QsyUusPm+vQ++p/VSaGNhnc/T7Tzul1rKRhKJyG9QcaEXrF0jAIFVZZgjfooGI16
c5e3UR4M25bwACoFX4U7AmA+1ruvktC9sJmRZrSE7BygWkbLXEEkmrFvDawBzjJU
FcldMGDWLYhqS24/K3LWSahTZN/mXmeLst6zArQbSsz/7odmRD3Iqt3sL3Axqnfs
54dgh0TlNTxZ0h0uCcP6FJkO+otXz4JZjBnPpE9AoNgZm0aikaElpQMwIDQe/2NT
rVGLBa1LTvY42VqndEUtYaluxRZd8/sXtsz+CF8V3AXdANZqCy7P7Bw32qugnmmW
kp4aJg6JQYZEX3v56gRJ0TuK0447MKirKbljvAxqHcZXrPwH4OjYvTNFCQHQW/n+
/992SrnTewRF+HMxKRHTEYyJPzdg1pUaH3Vv2obqU6N+2a/FVLS2M6Nby2UcQqXL
+1jWMC/wMEElR3Y+t3AzU1jkvK7JQFER47+8w2zvIga6G+XbE/mEjkgfjPFZ07Nc
NTuNEMJAOeN4kbyeUWsrOh3Sm2PITskevcuHlWowGdpamwKAqtZlmzV0PwWbEYdb
KE9u5Klw3LrF3GPzzOs5wo5ELG9BQ0hSfuIettx/KE9ONSK/heWqpuDU2i1WgQYe
F3mMjBLvKeELUnOylE8ES9eGTZuddQ2aVXE0zafZg6zcWb1kA466vOC4oklR7ygt
UXpVKctX82gBOBim5tDlZcQ6O9r2xTVac3nBEjpHWJ5hPmxInWjtLmjbU9kFxDHS
H/yo6McIRBhOLUxm/CnKKIY5WVLPJRtDjv0wQcGqTWf5X1NX/0WriLCCyVns/WTU
ulJ7JQaozTaQ4XXHtM3J3ncORl9U8gKE418MkXhBJhQP48EcEbrjyZIyjpIxVMfW
vmU9mECV5WWBcpmYEutW9SNrPBeTEBNrUTuMjgkNzeR4OZX9mKP3XaW3ITgy2Tyk
WmSuv+pFLDFowficMNmAk/R238ym8wRzTFnqo+IDSS3/RwEX8O9UYwDBWRAXICgA
wXQt/GsW01NV8r1dn92hshgNUCRHcY6ofnQsp/20kfVn2oRvM4masCbx4MXfgPrR
CeJYYIzuPeYCnKfFLQ7p7Rpx6yuZT3y76bA+drTxkyH6INhTOIIFQqoRVtunK/Vl
bkwkAn3k4CtpCz7lLF2sMJkWDu23A410QuN09A+Cic9a5qTzFZR4tVtlp2v+YKyo
qpDGFgcZYpOP0vtutNGWmavQhNeuO9EfQ3gsVPbXmEkUnf6xL2eJh1YwrhMTmdjS
wgdkrFR+OxsaTMwV0azeSrpk+k2tnC00DedXjCrMzveMZFpQ0hCtQqniAZ0EaR4Y
RvTWL/KVewj8JRo59bWjnWHG0rdKFDFTN9wELTxgvTOKdcUKuUfLkttCXx/rEdEf
V7+ds2/jERqBoe2+0H3BzbC6eVDqYm7m4iyK94ZvIFj5pQjfPTZ3T296QRY5j9xa
6ff8lPh8wlKgSb4On1DNUU9yRquPKHzUcPrjuqWeG5SgGwALjfl3OD1gDvwM4OFN
4Etb841dUoUlJ1xHV/zV6ev5L/kGqV+jywQF9LvNbUeSuNx7nZOmOaICJnJhPkRK
58S1vT2CIC1gZzFL0j3jCL7b3VCFk70Jo0qWm3Sy+zO+ffGf2cbHYu1azNHTaOCp
9jDUrv/9iJY2AO/sxVW72BcQAR/XnT8/G9rgxz+yg9NfIBwJAIYYpGvSHhVEc0WI
9USFbKPhRroZbpz8J5QFXRfeVwuqSifnnpmVB8K8wxLxKVUGpg/X1ZGouD0brA8f
CpOfIEhhW7O8dc9dPegnfNoaW/o95dxfJ7LWUwrAIGBU9LRMd7Ely8n+Dx0/afaR
suQ+7Hn7f281OyiRAjY43+YWbPGqSaCVEsblOPM0o+seN1jHzZFE6RfMIRuOggnK
+cYXfj+Rv2SoXY2XvR2hDaqvvLVr7KCZ5AN0+C8wXVHx1LZz8oU1F5ALbb1xlxOQ
J5brrEaWKEkJV5jQwzYuml14oW1LnrK3uVnx12jc3eAmO4ORBu9x8f/6rlcovps0
IJsjuQHmmnc/kLTpK70M2rkrNPG5xvSsTQ00NOVmGX0NH/B9HOG6WNp25tVsN6N7
ULTpAag8gD7NkFuQkwWbsF1nLWWq8LSXsDl94fkapM0W/zEsUmcfd0afXCamfiUi
Ldh2buNXg//DVKvsV9xJsk2xU8Uq0zV0EQpNciaR/d7HgFuQEtXJfxmNybRmRPpI
CsYOocSp2WEndg6H+PFqe/8i36q5tdkx5xiF3atTE4zrCePtKaaHdlbUdc5v6Tpf
xSXchvE2JCchI44dUA3veKs1AOVoQRPHoAfjETY03zTZWu9SeK0rdDssXPuuD5jQ
U68L217YQ38Olls3d9EwG2/Zg3FFpSUnnnOZrK5Ona4F6lvWI3pu2sn7CqkSwVE+
FL6TIC5d71L1E9NgvsNZb4qnd2TFT+1kpQBLmTK6c+GWM3p4nvCDJsoJyOi1DRSM
IF99HuHldRDrLcf6WeTWKLmGeL3R4ycAwPw6Y/Rduv0qWh4UR+ulfhN/4FoRdOjo
MNjToYAAqAvTIMq6vDMDruyPzi84kGbqnbYKcj+Nd8ODDqOChU/GDY+ndcaJIW+Y
cCsHet/wufr56rRU9qQRwnWLp8OCOwiPifxvFzIMMbrOb4qUBgJgDPdOl+UYeigv
+N9z+xNU3cBx2BGUoh6GmuCxNY9mExUtkx6powPoM4shS5GUHuohOINuc/AAC9kT
JARJGAhfyAsi6cXzIomeXPS+RIGW/c5JTZO4/KknYhVXOGPl0hbBUrcHaSWEjZhp
mSVNTD7jiXJA1f3yZ5djDNIVwY3rrZBD2oxwTI2pqueZe9HLUyiuxDhGKiLUmhRb
xQdawBjgKeZNF1jNOBkERj/oBR/yyXCYXUWquNUuQCUJOrX5cU0C72Y7bo+kdOxS
HL+fjUsK39i3XTq/Bo+tpIeUbWzZa5EMBXlOfWoVUnNrtE69isO8EGvxn3KciJqF
77AZll9o57sGGr4TcD9VzcPnGnYE29eQSYjtqM81fHBHl5W4NmBYbZucV9U6vFte
b0ZJ6TYLUUB3NcJ4logI+33NIS+WBNAGf8BzLw98qxfxW4SqAwLBjVhbizzadbQb
LwjuuAddhQ+B+sBAOtM6/lYs6FBcLb3vx2YJYroGD5ZS+C3B0vcHZOOhA7ieIZDS
FNUgWSDe7gjTWOSbueWapylP3mK2Hx22hbhR5SXn6m3ESethsP03piZCWsbNtLqM
VyS5/WF1qob2vJeeon0xEy/NQqWhKuNPikgaWVz+/KQeJ+rfgz44lVSpHs1lXqLB
XwbCiJOQL3OYgTeYVjYGjKJR3tB8+1Rc6hoKbW2rHhD1KDEhk2KbeNwUV053Kotf
EDM0WjxVCBNUxdLvLcakK5gxEseMxbh8b3dI8G8EtQ7dSVJbRJhqPZNUN3ORyCYj
wovIEpYW0O5ucGxx5f3q4f3RAMNbP2HkcppXAQzKrxRZLI8zwDWJPHVOiCVtfneU
qVYPrFoLGPdC9IEnaCCW54XKnrwMc1NMubgDljRtnaVTtvFs2gI7nDwZ/HgErhY6
Fzera7h2bqedvcEMPx4lomwfRvd4MefXj1IV/0yknj9g/w7loIgfJkcFwAbz1sMk
LlMAvRiu3h7CcCFlMLr/3PaswP3e54PDWLCOT2HqzPewPSBY4lselrhy1PYa58cL
LJb7uQXfNd6mkt50BqOAGbvoGkr++paHgveaH8p8lMPxyW8+YtE1V1HcgRlS/Wan
Bo2HKRABeLpik/niP22HNnfMsiQDnqEC01mxiVOYc5szJPDe2w+7yHT/OaZebV15
hm1/3cZfW2O5QGXJbD5x6uMpnWOfm69Y3CMje+VG7TOuucajs9hghn/VZETlpaww
PKeAMBNQzkDp0UIVNRu2HpnQHV+HkpDcWfptkOZNaD/DjfeCQ17aeymXE2O5Tj6d
Kna+JMixSC7jP6w+jHvsRXiUs1cVdfTLWLZCV/0D1W3uA6ldoMfEpsMBNh4Z+9SQ
QUwxJVLxW7kDPUt10b/tMuUmNwz2sxtebb9U/IC9TLcUiaKgRjFjrxFQQKDMRqdr
/RSOW3R59oCeNCMVzqAenT4w42KfPVy/CLH0rpxS/lbi/wgZ3d10nU2ijsBjSzfR
SKdUiRXHng4pRkrccAXVvSLxBV1VugPAnDhLspn0WZslHAQHqO7HvfPi9VbcCiA7
0dxWDf5pxLt7c4Ms0QftcHV4Ej0o6gf/AYMuWVi3qjeseU+bnbdFv1JoNrhSSp3M
89a19xwfSya8Seo//LIsFLTe0orHI5WQ7Sh8k3Qo/v/cBZl2r/AYf+clWa1FJSkh
mk7OZMELR/dpC79ZbnEu9+D3McWONeASQnvfGO23yP9ZW6DSPb3v2tGensmT1hut
4N0OhnoMECVSFA1HIjSu1K7WXPAjgplOyENkVR11brfhsyIEcaQIVKhMixB8r6bb
p3mR/VFdW0PTfpD/QXjMgSmFYD5KdM6MtxdSgSbo7+UPj6kZrklqR4pKo+YVAdjh
/rXiw/6CVFyLBZbStPjYO1dvcpQRFPZEPG7bAK3gS+T8bUeHunr4W3JBmr73Y5EK
bNXThnX1wRRtPDGI/ilFaZIzPiPooE3DodRpplxDnK1mWU6qDEsmXiILY1yoFHH6
K2B8mO7Z4XY9Mk86gN5hVqiK7BY6rNoYx6lGTmbZdKQ1LLUyLw4Q9dXoJwHtT3tt
qkXUjJUCtIQdmGXRGk9KrWJV/bVi60uhltTdjcnn2ICwYDWovj6CPIJfREvgKIaa
ng9PNzeo08hSd9JI3uRy1GmtE+JvjUOopRrjfDHZiYq9UrQ4cBRIWveON+gQM8Yl
FglsuCVWs6MvqywDNOrOaGfq8U17PArx98G8+S5X+Pyw8MCJSTC79eOMO33UhQYM
jQQqWDq3EIBjUNw5FvkvkcJE4+//if6bWXHXuPx+D4bBZu1YWc+6tJ3AllqRDuDR
vwUQIY1YromtJtYGDPjx43CIXt7UW9NxI/4/M480me23k3O6PVDi945UJIcsMzmc
jdWn0BXJ7R16u8PQvymtrDHpD0Az3lCCZ4ir182brBwTHPzxn1GKjFkRrHp8rXNW
O5nieObwulRJPQMPwF3OlNA49x6kz7GEQ1T5jbqf9f2iu/5HOAkEfw44q9VJZoug
16XCjYKouqIIV0hqp2DxELb61FnruDsbVyImgHZ317vxbIj0BpHSSarlST/ZDmfu
r9WvO+mT60HrUH18z4WUKH8iIYErrMBqdDv7pSN+W1vm9+HqsmrGYi+V1/KeIW7w
BXaDRnkBOzGwgs0rE/HIIfrYhwEr+t+YU0f/94aPdJmlNcoc7IBrxQZhQ4uG65Yl
lYzzssfMwts68dCrws2uqPS/m4b9ZWnloDqJTk9KXwKoea/npgqkUo95qOL7UsGJ
D6M5ivTijslfClQ1I6VWrsYXDkkDTIJ3QxCIsJ1l21em/9eahL8TbzbJsjNAfJyv
j0ernKEeE8aQk1E0si6OBnh0QnnjTjNOV3aPwGey1BGfVvoHVZQSNcjoDIcRtbJ3
t5HATrtySpuTwZpU8XOIwxRB3nQPJJ1E4vnjpEaaWjLndI7Hiu4ide3PPo5K5Old
EEOCpnQRZKlwQhJVpCcAJ+aVsvqeYeF0YBhxgl0u9zzSlD8+M4eUfwafxaHT/Af2
4WZem2DHVaOixAYT0YVrheTletIVojYsRxyZIrPdhKBFM7gNXYwGdXndJoYEfGmD
uX1Xy1DfzHRjE+iHCDTKpAvQ1+t8Nfq/13JTwcvc9xFVu2s3D1wsFFv8VDk8jRuu
iZmf3AFvINBApPVFTFBqT3Clzi8UfeZTWDgkCNKBBfEMM6v6IW4l4gcfIhE42B8e
mWMHElPd4TsfQbDqg/fGNOp1/i8VAl6E9QjBNfGNNF2VkTfshg4RGvjgB3GKpoOa
xYHB/Jwo17chnVg5XNBVl6PguG5sNY9J+n0GvIjoO8DiMOfqdiUKzlP/RoqET9nO
MSRZIq5Ke7Niq2oikuxq/72DRi4oB2YymoIot48H8vJMQIRaCLwSzPosRHBGi9aT
/0pxyTXcSc5ZRnUT6b4pXkBBlv/VErnuOmbOzH5RqGqC5o05ehskVL0Z9n85PGkN
mqWTNbK8ybR0lzSWW9TLnP5SDAvyDTWoNv6by3/9ziHh5sMFNqgBHohKrqjGi+rF
wWQ80FsSVnGU7cr28pjl4O5c93n8ELi10I+FNbd30jbvPRsDiiKeqAXwYRsUPB5F
lzhgghuD1GgllayMxC6CE9uytyljn8ilMMAlcgpfBEvLUHnaDp4m81+2cFJtI8Vc
KHuf9NcJpjXmh/6Rr7HtGS/xoSHDQpIJFYhq6dG661XIYJZBf9Y1usLQ3/+HL+de
6q9RLgteOMl82oN/+2+TGhHowXFaSHYoW83E0hd2qrE6T4fRD7JE5Wbqjr4xttEj
s5EOabPcswxSR4g9+qPmnySjVzkb3PYmpLuv/mayIM0eLGciOwJwTdyyemK8S7ek
NFtFtkqZgpU344eM2mUXMtyw1Kni306ny2f1vh2BT8g7sVGjxZuFBwcaz/YC+aio
dz0ZXiXn7t4RMzivU+0kIL1WLcrq1oxd5eAvwk1AMnTPd8U90AQ3AG2jxyQJaxP+
tkFWWX+JaLCYNXtyw/NlvOVu3k3Q+t6qd+A2b7vbArwlX9H0yyd8Q2Yh+zEBRaJ6
Q1jM/jE9ADeEB9B9Fg91x05K5ui+XEcAxZR5JyGhaWeREpKOylrpLG77ZALz+IJM
u/yQYjRpcmg/Up+3FO8fV3PABPldkDsdd+YDYXf7XOFrcM8UwLCsq2pfcPvaFMYV
P+SHyVcfjUQavPw9mT9uxe0pFkkgWkcfeuzK4rIQ/VREbcI/z+wUmH6P6qlv3PqC
VoGjZG2ugjwCsg8jRWsqMZy+c9ATQUmulIDuWB0BYFyVSYDc4VKPaPq67mODG0rc
sWrYRpUkIKvU2yl95fum/DZ2hUjlPOiPI5hJOW96NOZ7jPJ0J2JhLMf71KphOraU
L+YKGUgxfsgBKqFhvSPX1Kd/k9tRTTsqFZlIzZooPHqhNsvz88bM+jznq64oWJwS
feG/K1mWh7iu8O7EefyACbT85aHBZ7rgZExGpYOnFDxsT+m6XduXxdvBQMU6kKUo
pJiuU9lhWJA3L2mMc0E2D/3NvffjS5ndcO/eFca9hf75ButgqIgj5rWlBGKUJ8ws
87mkjiKmo/KAKKv+40vkwjS+REfa/a3haV1EyJ3MwEHINaXP8ddDQNC+MHmLGScK
eA4RiW086N9dANLAV9WVTw3lVyhUZUkVRLTWBpul7/QaMERQjQlBmcyEgOOsAcBN
lgOdZHhtQgomIs4GS/eGVI07bsrV/o1rR9unov/9sGcjhS5vBcRlpK0q/D5IrNyi
jik7Qpk0dIQJB5uwxGNJsgbV9nzKADNhn1f81IeOnNAoiOlZKYwVa0So2GiWLz3f
bFZiBV1Ern/sieX8T+IUr8PC9MnYvvUjeR/z5NyZ42+HXZLRBVeI8op2C6ap8dfS
JSKhIu5BBD78TCHnQN2XEs+fYsBsl4F6ywG0BS4kUoJPY9fqAz/+XEmILNFXzzwh
jeFgCIc6zifNw5fCXaCwZcX4yV3PBk7SJuhBQUoVSdhJi0NoANdYQRXJRTr4a1vJ
njzkB73MeLso2EboprUJ+frQy2L0yjyL+39w3h8OH1Wf/J73WEbD8LN06mm/iTFI
pLoFyyPxniAV2GBNk2pgOY8z58C9r6Lu98Y8end17XrATRUSvGw3Ty+00djR+XYx
8zSmgsXxJ+YJpMcPNxumEgHLFSVdp74+ENFubPKDTXF3ZKFOfuj1t+Z+0pVzwBW0
h9sfs2IasbjE9ZH44FX1gTG2xvvQS+WA0tw4A0IlQPm9Q4YywMf0lIhzbXK/rPkT
uvw1aSXAxAmdjG9n5efJzK0fqaEZO78ZkChRNZyUV25bAcRIhjbTjHRNHTZfjHWs
LPuwcdEoh/BM9rWdXswijXMEoQKxRsm5cXQn9n96MfqCD5R0SeFOPKz2YHljUjvj
R3TJfaIJ716DLaQ8Vq+DvWBKwvTLk5K//AlixGCwSnG0N0TLRiG9sh18hnd/NvWG
sOk/S42oP2BaHeYkd3vmZAy1pz2reJL3YCa72niG/kEtWZSIf1AMPvMB25JOsNJ5
6lPp+5/Gj99EPRn/3oka23AoDwq9XfzDgplbSccNz+AWHFW+C5EYiKN1oae7w4fh
Stco39xejOzPzbl7ad+FVNh9FJEOJpgpcmcK7ty8qQYw03gR1N9TbVaK51Cq8OXP
J/S64PMRqStLQMXGV6UukpyGSHCiPSHdOX0xDsQXwjpyArZCUJNZzxwK5ws9Coxy
94kEb8yIJZ2S4oV1IiOCgni0zuSw5932B1K/MhJOSnNsYLu4ad6OjCn6KqMMtayc
5ariajXSdHzxRTUeb1gvfqrAL00l1hWpbYK4szg77YlpVYUXgMEzhMUnD/o0Q54Q
Z7Pcd3XXuxUB1ESZCdbTwav+VofSPzI7TZBu9nJeaNgcX48zkCkZARM0WFo9kXin
iyj/WRcCg0gwo8obxVV+Fi9TuSHR2MgP/qDp545g9NANYJNr96ISh9m803u1hVA3
lpXH/PlDJ6ibmeh+hjEkyU62Bt18cSTlBLzzigVrshKKDYhLtI8q3KuaL4olV7pp
JUcv9b2EfGU2RfDYHa8wLTqwfk4wB8aRlYIXspdw7czoeZZpqbyWqXkN360alXHU
IGMRg1g2qU4T9CDqjp/Zf5FEm9isouaEHLToIvFiVLjVllJdaZrH+SOAgazW0Oeb
O5wR7CInv+xZ97V0PuDP1+6098GylpI4Ademd4Ab1ZxtijfRaaqpD4315gH0z0dO
PSyQpZcRuAJwtB3IgQhY8/QQ4fgfXr9NOjn7tnbswFU+sxPZRqGmY+Uve3Nu5Cpl
OuEuQNHO7MwP3s5jpogb8NQdazx75p1KM2x1pNKUA43JL9/XC/3APqHM3zQjRvRF
RU1NOzdPt/VrbxrZ8izqnOIfU2NE0RMmIC98UFJi+Xym6gHcS0dvUUPVJcKONGfF
y6VsWY20FLPjojgry+WRRS/HcIvJENBob9bmbOLuYQpHl5DNq9HnmdVRb1IchvLZ
oaZF45LVNDh4Bn0HT2bdkBEtjb0lhdKhcwBktT9wWTzPnv01WCr2UD43JZLjZtNg
A7Xy65adO2mNoanYJjj3FH6VxiHSfPCqBPMtU4UZj/8S311qL5P2cZTljTaWscAa
ipOmu6MwwXW4kTULPRZniIzaOEJxhU/RepJQsZQBFC5h9xjaGfbV0kpuMNKTyRpM
l8hCVIDBy3ac/VI8/bQ7+UCQSA8Crp2IqDwD4yf4gssE5ZeAYQHkSKhsUnlAO6cX
plsTKw6S92kJZeH37/j42FjBOGbgMwFhNzRIY6Zhk25CjZGPClNgF+OiZ5tVuZeC
xdWJ3+oBbKp8wE/rRtBjHIN71Puw+fIyOXxj+8LY6Ul3wTL5SRBVjEIuLlLYU6EV
q0kpJcRvJufphhtyI+rZgfYuQOaabn3z5F+BkqM7cpwmXe6+5GdGa44iRq/g61Zn
K5azXRPSOY1xxOs2S+hYC0nqgfjkkfpjz0qnn0ek0YQhSVZQ6+5BgbRS3QWrLUaA
RMLcWpkTiYztv9IVXJuT8Mv5OxBxrhpnjmLuiTZTkw0ywc0vaNYu9eNyJ3Nb9ZPS
USPWEDaUyyBVLF89VZGaHqlOLjHa4sj8Gssp0mmweSzpaLwSZsHtknHRBN8lMGKV
Q006ObnafjSyi+JTl+QRtQm1X31oedGgHAtELw6sBBfMiqP/xMlHv9C2dMXz2P6t
7e8Ov06K4lHUSY/FE98hCdt9+e0P0+VyMIi+Qle2dEqTcBeO9A+e4/JW/l71ljeu
9gYRuF8HyLL0j1kKZkY7h6UA/T1KXQ2dBaZzZUepjqCNJKm5aUBSSR6dO9L6vkVS
2zpLa5buZDBZvfZYE8V/yHHgIPF+yQjwhefLl5urC+tHkX8QKi+VDvPoOnfQIpqP
r1429Pvn+zOCVNJ3/N3bc/In8HmV604YybhJE9wzJw62bc7l7I70T/HZjTmrS341
MEtowekAssqrsKBfymCvCJTZByIQ82VbWYDYJq6Ooh6fY4kA3j/VV2uwVjOx6uOR
DfFaa9dWtSHYaVHBkRGFCQR+js2APw1fqfK1iD8IANF+xTPmAOoRtEFQzf/8oy3a
jHfd9onwCEBLOrDTEWSpN9lOWCRDeCafrrQ+2cw/0jv+9VpHZkgnRipYtHuvdU7M
6oq0lnB1r7RUN6biQEJMhwvM7uIRgBifD7f7CFRYCls4grmGO9O5rT40DSU+LUlR
3i2zESL8NE1zQPiYB9fqLjjwgon4QLEBAtgCFXPZB55Jww5IBxnrFha7Lt/HWoUv
6r31hy1MVNqnH0p9gUV8+ZpXJO7BkBmmNVhChEklRX7yqGpTl4yMGrFm/nfpp9S2
cOfAfoqabEBFhgsEVQ+pU6Sk7PZVM436R424hI1PCH3ROV463gC/pKni3SGpiDDc
JeizuaQOiWbtxLbAhAVHfTx8aRVukv2Q65JatXyFChhFnvY7av/Ile22ZKr2WcuM
VgpmXySej6m9D2YbOsI8AKMF7WnslB/VsFXqsqFq7A3aJHCJnDIYEnoSR9q0Meby
3Cmm8rZbqPESNjVdieMbGr2fFAp31Io5GbKjl6FvTL639VULqkLp7PijjC5nvsuS
hSmsDT7cB6DwJ93j9mByuvg1ni/epMBIyaoqKz9mS+h1PgvHciFijOI2aqyRFIOs
gJoK5o0tjIkuJbDEERwy+e0ZsU2qWsZcFxb8Pp+ukjIsfLKTtQ+6/fXxQNxaOT0i
dbJ/m/qGd4eu0bMy5WTiMdWoS93gXcGUaWgRqVNorwOY2FcVpOuNc7Jh+HsF4MEs
yvJSaToR6TCQX2O0pWGqIIuXVi3NVSWoh2s/Uq+aCIocVVA5GeD0aAw/CCBZ9Pvn
1wttK9mFfjs1kqvKaitSgGO5rMcLfBxjAK34HNSAz3sVj8q/WhQ0BNYi62elORmU
fMVj87htxVEJClfwviJnhx1PpSS4yHYlxkh3PCTziYa3YiVhV8D4QTx3T4+SePZz
GjYSF2GDCl7oeWvStcw1H/OELzE5NTMl5RIVBKtb9sV9cysvSKn3QMOAtTgjrlVP
NsfGd0nyBDJUwpuamZEyDo8oHn7j2eoGYhgf9WVCLuWaa+GqKNgnI1aqVYj520ZP
j9cbSVnFNDwzEneJ1/HGnn6a1YMmSAvBAyPehBDkJn2yLdErpzTD5qFcGpUJGpaL
km4nrJvFiDy4nBEy/FgTOahFXc9uW4rDJk+tZgePMOFMAG/ewXhkzI650ki3j2Nt
4fPuzguxzqN3fFIHPVUCnMVtP7ly44R/3pteAOwXvdJiF7M2ObDss/+CoVrUfpZM
i+d/HphagyweA2uhJWwWaX2kKPFRd3HUrT9m5yBKdVh53tnU3+jNLBU7s1qiGmQ/
KPLoDTGbjlFruHdy8Pn1tWc/R9KheXWtZYSI/mzn5cTI/5LuHb7jupQPaUeBn+Yq
EgBofupU9b6PHjNJ2DN8itNz/zskapnMUkXaJwDRGnKxY4M5+N+yFKQUVqfkF3xz
vEs4Ksno1YNXW2ARSrmPN0qcRLnkc8DkmA33tPXu/hrZgNUKDY/aEJE0S6y1SJ8a
qVPLIIFz4xzEgD9/TXacMSujCVzstbtoc3HsROYn9fE2drC70a3ctS7TPm3MH+mx
MUXIX3Pr+zen9lwMaDnjJiqJZjUDt1KSV17DYSMvodmrMwSLIgn8iHb6ag3CWIvu
A6fpK0x5DMarYHrFuFYsydfYY/MPsTs0fbyo2nVPI480wkEKTcMAtLIw+CoQeZ6I
cJodINpRiKiBv34R0Bq+CWE/vJWQWkqdRBq5C0W87FsfRKa9U0xJqqaQxmf3JgTC
9BETYWsJ3qx8z0gsPxCMk7ko5HiWKc8buE6fWZadmVcKrvO22whYNoFzp8CD6W9o
uJeGpKvskeJN1d5U7hytFsfTo4Pg0SxCWU80i1ifaZfT0uQFADzG3maASaBNr7lJ
JPQT9oeVii+1m6oc53FSaamd68b4K+ypxH85yomkIsXHcTcTQAX1qDsD0ue9i+my
K6UiPpJGwOfDc6wgoj5FEmqd+W0S9tmjD3NVhwTDNMmP3P/vnz4eytgVmA+OLi8h
B33IXGLPnpSEJr0ga8+DYLu/D57aeqWvBwwXry2Km8L59/sWvqV00p9U2AAsDX2r
c1MLQ8b9SC0r+cbGr2WbJwnN+UYzSbW5b2HO3otusqztyuPsPaB0BM1ayqaNWNVv
0F53rA7EBJARiOgjKk5Mesb/qe7M6NVJQCmyaa9pmGj+kFwP7SDHtYZvuPQftv6k
0FKspXYbs+Pgr2AcOEbyCw/3p3EWiw7VXsr5IUcQV0wH/DjDKxsZTCMatKfVAZlq
nAtn64xLRxrnnd1e2PSiaBSpP8KKxnwJ3cyEPLwRvQfluKxy/weG53uw+9TsAZTl
ghpWHXdSJwWWABIdP1SYfhWlkTJcdVpXMT1ZbKo30DtHsjEKbM3D2nMboDRj4phF
Ob3VRfvsvQ5TZikQKFBlK8ppagYmui2X7pSI3PTLN1EHW00mV0SEs8jUcdNsWjoT
9RJwa80Ecy9AHPnHIY9PawZbanJHRNVIqyqDMJ3VnDfhAX5XalyRFyUBBNz4ge3q
XG2eQvkJvazrUwa6ZpyAJ6JHU7zyQWpSLTGBKVXTcZ/zakk0HBpAsBOFY8T+AD35
WEjFuXF5U5MQyg/KW00TbrY6xFG/gfu64rzGyeBTP0fIFD/jiA7Nw0l1M/Awvkgc
G9t2EDjkZ5FQCc3rCFgFemF3cIdI7jDNsaMdNdn59xJXiJ2lVsa2PApfhEU2VpR+
kpJSKg5tMu2CfYUemdFy0TKEkqIkOkRVPI69euu8ST2Nq67VuRtOt9bAkBWFLmPX
B0kzK+0llEXz3fw1YHzMqp5LaIzJ9/qCookNQgxiw3en8cBkSdz7R7hhXvZYcEPh
cSD58WyqC8iFrjYlQxBY7Z0OSCXTXBsrYUc9gm+LplKErlvfLrMc9EKghyexyVCg
EICW4xc78lg+xNvT9IhmWAnkQbbfrXCoyzJfwu1SETk4M0cCic4Ekn8X2UWb4XVG
tKPPQjFr/3307maVdoDcGpfkZfk9DMVZ5RSykwXlzOdFuEYZvCs/aaS8wkMfaMNk
CSmpPoD1Xn97jOkb9GARBxdGsLxP9vbXSA0CMlxxzvSfhqkI27kHYGJn8ArU7G9m
iBIBuoT0k2Ht0btrku8VgAjV7e6lF+dbXoF3W2JhAB0wWy9c9EuSRrHI00ldSa18
o/+Nqs2fPj0em2TGjTOcQqfiPnpLoq4Z8F52G4vX0LzP7G0YLJlkfqpuYeFfbryE
HPo93PBoP8y+aDykdqSzFLVM2Vsk2nVmBzJcqI7zQEud/tyvLQ8mpcdBiOnjXLbx
V0eeTjlaJnP+WOQxTt2WHYhz2d8OzWxQ8gtatNwPGe4OGuXUNlIvDT3kGAYwEVlH
V8c2G/utPSH1BJ9Yl6WAIQueVtwtCmb22Dei9/2v8s5CyjmJY4yKSQSrf0zLqSBL
F9MV/+n5mknNGzEz/jlsDMrzm2ZqRj+uqaJ05E1MmE1O7FLrdVsanMmdGDWyCn/5
C+3y1aDdNfSsNcl9UlbURPWmquiZqNMov0hQ57Z5qRObPWzwocRp4+KfizWPph0J
V7nRAeviiAmJLVahycltUNikII5amffgsgu0KKdS6K8wt5pJe1lvICQc0xd3dMoP
zk0+9gcfVPbVkKx7rr+cIYCK2zcJjZP2BHZbXTbjs0tnp/XWccHv1KSew9yZALmJ
0j5SGWAbtH5D4+UMwT370FAgFsrp6s7sv+slAM0h06bcKS9YVwTixuFqZqK361mu
sn+HTY3Y4/U78G77kFzX0Yu3NfdPmzablq7Z+M/WaDEGiIdubZGx/D3bmbRdXoGX
sHtt87cJi3ZMxyBKgT4NWYqccpPN40JQEDsd5RRHMckiVWi6sLSTRNdIGmxk3AQb
W9N9/msxZyETdAnFA3GfB18wjxQGmHpefZYLsPzsNOvOXeHztIpjNv3DpGOFsusl
ltaDFusGjTUikLF0pDTTYV9Hs/Dn7asbrUIpEoph/c2nH72OgDW9jtqh8dQVfy/e
rGp8nTisFnJ3jeRyr0O1OiMpGrnDYOxJ826frWTWKYD6SuBnGgKjxRe7FXgHpm6p
fWEuO0v1E/t5JKWTw86fVcc6mRguUnA0OtWuJRH/Gj2U8dIpjEnIzySZYcIL/xjw
uQ/Q83iwGl88yr/EMxlJxQMwloclWEi8+UltkfcQfHe2K/LtF5ghXuIwk8b6FhyT
v3V6a+acFC0wiOVpvzXhfgCm7abgsaXuJJtHwW+6CipUezwj36nB6U5sEchbzBGg
HV4ooEZxJ22BIBCnuE/tUh7Ivw7zhbStaDaXZenBPXQaTiuz0k6l6oCypHkQQP99
R4e0KFquAFkKdjgLbtNBfdZGvCCEHsNbjrkO5nbiCY7E+0RTNIMTY9MVlXoYoVnu
f5Tqikbh9R3bHIVC2HPOJ41gvBJxDiLY1VqNF6HNpJi3QTkcxCPGgPmEfEu3JSrh
qc5jWWgUetNUAat8zciBemR/JLki4DfnbvEemzbh3bMA3NxKzPS1GPvUxRubVnCE
i6UWXKncfUsNQe9bC3mnfFUGlHkQSwIO+KXKjGBZaYUPENGJGgyRZsW2864B+Ts5
EDw1QhymRxF9XbvItGuvC/rG7yMscAyVlO/Zt3+orYQ3PI1B0xdcEh64rdawoxka
RE/1d+dnYzYr2TLRBLXWnrEnkNe6UQdgDAH7GMnusep969c3t8Ve1pcECdqhYW5Q
IcxPNB6YtY/tO+fTCBdtKJ9LjIng8sxM31Hnt4d/4F/AsCMJbfu3OX+8W7kVR8Kk
+0kVIAc1HTofsp7kaUvF46jKTz8FIw3CeFXx9DHs47zlUpCNrxRGvg4CU8Dru4Nu
SdE/eH+SauR4gINfxH1LHuzkLpkB4jtEoQVSNF9P0ADmFDSOMhxCPTq184FPSyxQ
WyBAyMqwvXuGUhM9XamUbbAUOhnQ9Yjeep0MmUgfwKpVEB16CCfrqpRjHIhIhZhf
+OxZdpUvefuVmME4zS9U1g5z0Yt/3vLpJi4o7stOHg9vXh6XaTEeyzZZXG2IUlIO
H1KTCpTYvH6ya83xX8ySvC1lkOXpGOaMaBbT2oL/x2xHpQ+N9FEOjvY9wlCR7H24
6dZhetPcDn+dk8oi+l6mcWE8ZLffGLZVOP2tN3QbMWu4wOM7eJo+CgfqYykWWKZH
B9zc+B7iQ2acsHK0yhfHtTDTo3QX8mD8FgAPcO+JLeB4eyUMo9eBNa1FteIb5h5d
wZ3xb7bc0crZaOaQDzqVntOxsOJ8SYrU6yEr3AeKoXq7T+3muro3OuzG9rubdmO7
A+TZ5nULbvbBqyTv8HxpOpyuhXnXTQWOc220/1jFf4lWWM+O655K7ONQSYS5xoty
p8Ud3K0ay6GSF/0gnb4g/932Lm+APbCURD/qPTxWLLPao6KznaEjuU2N/OFiXm6y
e49cUw2TMXxTDImLm62fKkLfmAl+GpRnnFvof2mPIWi1qj/TNBcfOBxFwThv7uA6
kFLdLho3RBtx+XNNEUCI94EmztiCD7gIek+pQcUM5vksooI5fx47uVVVfzBIX8bY
6gT8ku4wAi1bX4+TfV4XxzmPhjUP5UNR2Oychd4JJXmc5B+ngXAC9rPPtn8bD/+J
c9faCW+xI2Wk/5Ve1Qtrn0pQE2fuQ+JlvhmRtFSNNSXzVYYSSvOkcuzqPiGss5ZE
DCH7Fiyofrc6qFM3VtjfOAXW/uIbHnafY+uyWA0bJZ3zVsQfFBsJQFgIdnclCKpC
T30oyWx/NNJGy/hoG9pxDJq3RUPEH8tKNNitU0e4SFdzIajHlzW+68m0XTiuc8En
H7iFjHaS7q3T/x5Lf6qvTci2OHXcP7JkWHoAqIOUU6qU3VWywQtKCzagI0IcppAl
ITaLI1fPi+Y7BD7COQZiXVavCNzbBwvLCrEpwgP0dd3FBRIhaZ3EV44PHdKrQIPl
+hNGALi7HRqc4iMw/YcHcLpYXi6eUAvyni1k4nXfymWD1Of/Z7B10GMITsAP4+wm
87gZ8MHQIyBHA97sSOVF72dU4UFdXAzXm5xgii2BSiZ6jQfsM5uGJI7O5scncpox
RimaI2VBLbDY8TfosTQe0W1Ne8By5UPFwMoy7xK6nP+83xCvZ3KdQ4PfNfYWGoFI
It4ONpFGuguX/1YDL4m/9QHFWszK+c2WwXgja05uoqj/l9X0Hb1HGT4HPFYzDs2k
45q2xgKb5YnvctX8FD7FHf97+u1kmxioABPDDRXXRNLEcM7m3G4Ch0/9d2Rj6/K4
2xMQ/akp0WeetLv5bABwxD7g94CtqelDhI/wIZii/T3/NlkMW9YWENaEykADbk50
owwLjJ3XjQLO1pZygXn1f+ym12x1vzQMrDz3aL+6BpN1UAYRGqon/hF2dj4mo8nX
D2jI3nRJph3QxJ3+oQQw+gBL5YgYEJTn3Sv6P4s1kdvTVmLey4gl6F7y7r7R8ohu
9bDhk2FNjMpfjOfdB9LLipfljM76pxSbBY29gMUF4RgKnzLd9/cMf/Mu3kkjKh/v
aqBv4w1qAJPznJ/LpxHdx9uaPv/sHk1b19/bCSwZaaIHvjoSJeSPl+V5qsZpA76I
vmHHMRIRu2fCucBkehP4W2eGo/As9p2pR3SO7IUP5Zw5oKy7SGe2UvKKAHLRHMQw
CfRN0gtH7VgXgPqD3s9CULtinJMIYT27VaC4H33xzG3tQxlX0U2ukKcUHqd5K1Ba
xbH2ORiXz92vn4eK312AvfYNxAT3X8/W+igT43yBnMcg4Y2mby+gJRFPvN0Lqccw
WgBgRg3mECRF0ezdY6uY7UZ9+wsg/SD3S+LmMPMyeRmzfTuES7lhHas/nFcXtMgx
C0Ae7xpt1eX3h/o8JTf/rnREYmwL3/FulZuWegZo/bFNNL/wV7fesHfNQ8SFd5Hi
8Uvu/FXUs00TeIzyoddbMP7F2tFMFzkGHy5O1K4ASpou90vOSQG6kGhYEh4TElA1
FsHOF26JSOkmzTi2gF6FGaWdoJPopU0c9v/gzTk7fHSsYeRRPkI6LODysUoDWs5Z
X742OsUK7aDkDq0CodhNzWSaH0K7xSnWvwjdkHRvo134IQmo/aXCJG4tz75lZpCi
iZP/mpx23spNhHnOY2y9b9VfmH98tzpdmQwB0WYJVjW9cXh1+gzO6G+N4m2hia7Q
cF7Z0oKrBFpZ4VmTPAMUpN8xHB5VlZHGZ1BNGaTzEDCPmVueJWol4DDfol8ok9uN
JHCyYgrn8GJddVoBI+8j+ArfhkiwjqpZsFwmd9sl4ENfg/lMNZoN5W+qb0u/Lcpu
Wc5nTE/vZh1b3yNOkgDIyYcD82BPbM9ObEuV9ry6+u1r5jH6FKMjPC41W/3xAOVq
CVigR+uG+YrQ4T4rdBKA8qfnVEjeXzLsDHhtqWV0j5l0n8Pp7HE+GjyP9Ji/dPVj
WJzd7XyKLB1myJ3G+1lUIQQoixbn0tZw8Qd/8cRzaDxatb+QkokBjaSpT4RzqapO
Rg/5GHARmLn5yDlzYNV+FI3vTMm7PgzSpHQbH/TPhtVkdE8hvjUDnuXJy+2owfBE
cijwdRbBar1GoOn3XczrL4xInM91VjpkVEXKEt8mVFl/NWmweI6mxz4BUMZrEa/v
pzKKjvuZHyb8XJO+qouYRGWkCgep9bciNNzWixuCqAGxFbZFcHIhBECd7B7gGRRt
gh9yc9ULdy3b5i6kNvk6iyzwJW9+PSD5HQyJ4yFDDLXfXefWDPLXKEDxvxHAieEo
2tna+C8qCNy+5gNcKTB0OzB964LcXSMr2pvaam60NTNTxzrUs++35Eq9D+NHS9Te
8FurNdE33kq6ABE56jt3tSzDUC8Wx94C6HXBfqOH/2KaCNZ05hrX2wHFSIZsjRUZ
6U0HBa2sy/7RfvSRF/5jAJPn/edMhF8pIYg1dibWdW1s75QPRdBahU+U8BE3nK3x
8Rj4tYbn9ZfLkLi0Kowd32V4N+GBNfoumEOXLhdBtXj3UoYJRs6JazaSDhAjTGra
zbRZe9Z4hZ6D2ejRKMeDZ293sxOSq/HsoImxQO0k0oLNcQmKx4tkmFdJ2d1d5qh1
7vvFwWCSM1sh8Q1SvYXVet6/Ir2cRxtFeKMzVNgzdNL7v7seohXMbFbw2Om1I8HP
uF/IOXZwc60KgcuibPo9WERo3qB0C++kRaC8Z8bum5MG7gAgPCNZ4fhGSGAhUYzX
J5HZvGBYog37hrNxyyNWPb1/QT9ypthlqyL0jWEGzxz1HrWqhXn1z805mdXF/xeI
6iDNL1FZWm2tYTOO/mErX16tUnVD7ay8uBVL9SzVT1voXoRz8JMwl6TPu5rdZuaS
eAFLav8MrvlCNp9F6Uc51hAewpiEQEuUpBjOASkzW+FFBnxa7a9ee/P2WCJxcRRN
YHRx5/fX5T/XST1EpRfCOEERwloTskG4wDrFt3Ywj/19P4uT43eWIuYfucb9G04a
uzeJwyIY+LS7m4wVNMFjwjuZKZ0bwvkAPNelcDLR9O1ySQlie17IeayWb7XTaTEW
RpfGWNwtGaMPjiQW6YtM+02Iu8USA1GUkPL0u92UxzibVf/koyur+RBIWSVwjkOb
jmxbjZG4iQApIUUekOuDeSJLh1Luvr9zapB4lickUlTxKNiQ72Rop7PHv9ueTRuC
3+PVuJdEvElOupuzzRemGr6o2sOVWj9sjQOYM5Cxx30VwqP67aK67mCKGhTCQUii
USz2GDI7uH26VUocgXb+WEjA2fc5FSeK5RntRRkHSRGmF1Z2j806Kb1llcej0VTI
1E1ExMS4nKDcL32cFGHfJXiRuBYpDmIXCnYFU2P0QN2bdqcHxS0J91lW38ixUgSS
yrQJ6J8mC7Fr0lqH3iDRxGTfjaElZermm94GltytVM7l6lctFOcPFJsDIe1e1vd0
Mid/q9x9FfJypxfJqyCgAxbHmGZ9RZ0GwFBQNhbY0lrePYKJcbxsWBjsatpeMpAQ
bZRINFKoTR0VGM8GjXJfHicv5mE8lebvtC5ESfi5ClsboGB/se0qceB4g3u0oIy7
igwh/PRG4c8wxcaDCSJTaj79tqAHsDy922CtjMwRSAIysN+vOw/JFugqXpz2TnGY
0HRZoRv1X2jdj+nqvci/Gt+WJVoixsil1xVFkh8zVteV6qptPv4xPN7WyuLTMsgS
PI3mPIFmfHLyVXo5qbGeVBqlC8y7od4M4u1t9BZBhiBs1c3Y2SnhsWwJQ1u93K03
DGmR8x3b8tPgBAyGYyYdbAeaRuOuh8Z0rhIOGEB8yuNCYH149zTingAyY4iqhOxd
ROoWJMeGLbzyoMAj41o9p1w/5ALUkcDNls5uDqXwfRuPi+pBqn1fG7rE+kNJoBMt
MmoyCZ8gHZmQ8mPhF2XehXK5/qIOjyiTwnHBvJQX3x/A3ExxNG9Tlvz8m7zhjRAZ
/taZz8rhuURxdAgeyxef3KnaXDFP276QpmosWD8h6cF20qZ9DTGfgHPpTzCaBa5N
M8i3VQX3VECK/kmGfwSetT4BMQdmtsRrqknMxk/5Beg83tHVDbGxKtQu/lEqOmaX
OEOOCmkJzKJY/AfsU6BrHJABEzmOdcerF/6zYhSm2Wk2cLxbWKcrTGjCkJj0HC5N
576vsKnoNsrCfmh2nhBfxaFhrVPQo+DHjkA1zSpARX1kw10cfCZiQfyXvllGXv+n
2wzRnThzd/BPfzb7QYbLzftKNNExdcfa+erAXgPjppYwBK0kBsZ3lz3O36OYp9e/
4hR735pCTel+P9J/xOt7Bv6PxN1j4aXwx2qwABhIVGubvO7Xi2u9Yc/hwlV47QDQ
AU2PWzC2YRLpIP5mwJHxAks5auRe6PkDhh4dw2WbvLNEG4+AuD5+rhQ44yha+UeI
kDLTHmotLjel8xm0+F3NdvXEIWVVjzjU4W0DQoPv7nWjiInpPhNqd1VdkuZXEtBq
MzQiAalrDOIu9BO2ATco1yPnyaelWph2FX3m4k9+VpfuAUtjiNKO8m7tFDdzTy0T
RGRejJ9tsHRqWEIkLcLIOkrDFPkOuvwCqlbHeFjUtxU5eg6Ffl8c9XcFAnvKDgyU
TNB2JkxRi9k6v99omyjMrK971k/6qwdPhB4Eb9g8iNqRCFPWjB26tW2vjUpTlwaY
libA6v9mEi8yBXMoKyQUYJlX0o0oSrfwaC/R9bOuj4aEVqmlm7delCWGH0EYRSha
MjaPMysHDTAzCEjKrt+nrzeuVd9wtuiOnsfQPUufAbotqqjZTQZKZfZUosocx8tp
BC9rGepvShxZhodY6OkI4UsItfhSYtKw/CV+eaILm5Z0tnNp5Tq8t0v2WgalCkAX
lC9ndcqgFV0gwL3EsPpdsTkKlSx4TbhhF88BvzLt8aydXKP3UqQ4D7sUEtTEhN11
GxqVGEdY00okIo+hwADNV4qDVmiGggeFpBSHwPkO5thwUNf6ns5j0ccKZ6Ha4dsv
Usduc2NvaA0xvrDb0UKyB6LC/1nJX6e6GgEA7JQ4MbVYJKek98YQ6wv31UWVqovZ
phfnwQLM/oZau5vpsYEw39ktfb6+4h1m1DRVXDhjuNxn5QbDFRxIt9AJ0ActtywG
nth8KzSbz5G/sfDQIRwdDfik0semHgGRNMTyGZYab+Ne9Mp7ixwmGocHbqqlSeN+
qpFt3HJYuCzhi9+UPtkPRn1UcMtf8NOGbaCZ49Fj3qVIKz7ST/zGvsEdyn1TNDie
ojilZQtz8ZMQ7u3lXZmyiuSOQx3W/dTQi6nzQqV0Cd7pdYJz8ZpE7bkIY7jKqZ6Z
g6Fgi4H3PVqmr2njj+lY3khc9zTSb6BVHVEmf3LdPuH88p10f8vG7Tq2dOFcwVw3
npwjMQroTGVCmxTRZ6v1o1J08yEAM7JhhHmCHi+MW40KTDt3w5Pld58DmjkwpQPN
y/hesVqeKsQqprqJE9V+uBg5cK7nljNH/XOsTpvm7EonddqMxNkiV1bYHviumjoP
roVfSjqqWqdYral4948aUHK+5RJ6ucmIwuIp64wnK+PwUNwvFgz+2c2kUtQiSee3
ArTv2W1JAp0v/G9xzk7Za990+zY7EwWJV2MHt+mJc6jZBRbSzu1UMI4x2eYeWjpx
gRjiOcAeUCLFHWd7dtrus84Dp0NLSybO2gt26Upf7wMy7hSRvPLgWW/Wp2nx43Xt
67LBohy0dhtLUr5wqc+BKYO495qb+sL2vz76569wO/P0TSlu3vjNpKyVvZMaXdWw
ldTYmrFUBgy6GZK3d/mVJEcFMlLIflos7tElwq3a54yUqbu1OfOKXueNRhjz8X9/
z2YxrknAfmvpAkAr4LcUjU2Jl2dZlo/L7VOcS7aseWf6XvggW6FNCq5NG8Y2Pfz+
dqOgwg1amx3x224iKSL6cVZ3QDcPsXsQvTdmbolS5ymtxk8ZcRd5WWvQAOiEYsTD
kzGVAhRJHOeADRTkRuPxi1a6uHtV5QLML5IOsP68DglZBB8/CKwZcurknB4IXLy2
Q+ueZ+EWQNr+yyX8/7qrS1IWjQYhxiTCF6CtNHqzrFIPjd50dVigyEUKLGEQgTar
ueMDUI2zK0bVDDF+NMBanO/Yzth/D2J5Sx7m9gVVdAZdF29VEenNbBahHnhpnJX3
Tah47Rh2MYAizP1UJKn5nfCu2Qp9g9JWwBum2WUhJ+oWLeSN3sRD9pOY+mCdeIhA
TCn92DOUeAGas+yRjt695fDwQ689+SKeaTvLvbPYZpUc6oGv+vDHlAW4E9OAIUUk
v+8/DCpSz/+qFV4Z4Oi3sj62SVp5TSVjsDG+IJkF8CuLEocxwR6aZuNC/yT6B0YG
bRF0JlDyrXuOcqX3HPwFMAd/iy+q9xFfZ3FvgPLlJt1LaKWmviSYn4AAW6BhUV4T
4b5LCIbMA/ggmmt4whBiqqK8W90C2BgVlSRley6HTAJbZ4lBPNCaS4ADu0TvcMba
mn6FNIWSUkDbVCoj2KyvfUPjtD3VUazxuDCZ1G/E0VvvQmwhsCgidPp5zu7n5h9u
QDtPA8CC3F3ExZx/o+3RszRBCtyDTvxQCTSZ+rO7TwY0L4CGf4lVw3NEBrc8Yrid
FHXEODXS/Vg5zX3S0qQugP4UgHxvtA4HWycc5ZrB7KEuYOoy4+UHzTjj7HNhedoz
BrBTACXdbipE4bznvF1AOxcBOiQJ/bo5fGi1+uxKZ5WZX9chSNv6r8sg/mmZjUNl
ZciBZOdmcVvi+Wi2/QMtU2z3QeRUB8vhwpAoTf/A05BWqoO76PCiNWuxdwEK1KVo
0KqH8APy4m7msmwggQqAQkyNCxl6eOHtCX7FyryCwj9hbpzvLH17VGeCj67MCjxY
8iaTLqWOaBsxvZJwiZx4PHNZLCndBOWz8Xi/0pez1XiYpGacm450rer6ZkXf4sBy
60h2uJ/KYduhFTpXzqvn9pA2NiiGEFbD60O+8XMPMyhyCEHC1Ej7nu2OotACxJdS
WmWWyzUZGAujdBOeVtHYRocqjhg9mJ3Z1Gm7DOLV5JqusmkZlP5xhWnv8u1/20BH
ZmByglDndpMgGLf7//1Pd5PBSy6EicudbZbQm2ckttte5NoZlY2ViFkNHrEHoK6k
NA+YWG2uS65TRRgwXro6hjA/OHaUlFGDX6l/OBzNnSMDHKuOMISSmmhrTeE2P9kC
lZfCVynds14jYUMiGILt/jK4PWtWn96OArfRxVfgW4kb7eeU/f6ayvIILEj0zDHL
aOSwnim624K96MT3SduBLKS8JETpF/v2h96M1WuMr2KRaD3zC4MYZ8byw3ODzyZa
U9uJzL4jQRIxq/aGsufouG6Gbf43wkqcrj89zUobm64Yr6O8w+cRqb6MvdzzvaC+
PnyDr4kUeIaCNvs055oAkT2e0bGDyPRPPhoz/b0kIxq8uOBL7vxQBPSt4Xg199UF
czyo7wQTfqePimLMt2qAIrugbW7hhoBxmLp6BrZLfL9Hw71z6iOZem01KB78JUgd
ZoU/GIQmrKhtjKYzB4FZ8mIhyN415lyy/KX4vA1VrgFB61fkuwwZqU+bloGfWGks
oA3g4OJ5k4LcHeYpkY9yiipXlHKQE4k9UvUTz86OENXkHJNJt4dDjmI2P1NOHbwa
6+sD48PkgDVlWxrxOqLk/+8XKRAGDsQdz2EqX5xlYDMbGDlO/mS23u++6XOnfnMV
ZwHWIbqLstr0NOSxboH2gAEbawglZQUZs2NHyRmdjhcVqtfjGOMpjxQ/3IIJEO0u
47nQJiaLFwINZRc8DTTEG81gJ20OU/ZT2c+pvJfVOR1/LqMzRCNztQK2hfbF+DIg
j63cox3e3sOMV7xaWWXh9G1cSTBAS9NCVr+JOsNjnd9/uhkP2TWlesjGY+WV+XK9
ClVhdzKIpjyh5hDx65HctJoasjUhULGfMoNVCAzWDd898G2TF4Bro9bID0Qh0xuo
h+k4B/ThYKs4kCDCpwotwOblV9diWSBXDtXTMxfRDInGTELRcToNWtDSjPz6DzMG
6gT6ZePjkUUd2rRSGaoUi/igKfRjE7DKDShtIbw6ZdfR6DBPCVXtw5nKq16f+z2S
1UBBIfxPWSXja6cZ6sM2vcfhPyMlY01JzWjN+YsmQH9eVz9mCJryVvVi9RrezJS7
tzeHI8HE8fKSK+mYLuhDaYnehaWf4l+nXNPmOTMk03frIHHLa3QCPvMF9VmTpALC
L1Je4YTL5IvD1ssZyubGzh+W/+8+UA7sdVHHrmCpHTObd7+/eDScYg+pLYr0Cq9T
AEmQbN+vCUMDKjL2uwssZj25K5bizdA+YPpHWCwLmfpYh3I2eY9BP2YB1/3PIXHI
oOGo2rgaEawCwWmGPJ6hdybGQNGjMypZanDp6q7GU7TKLciqzevISYwdepw7YkYa
1RL8AcZJHfJ4DSTAvqx8nyVfHYXt8NyC8mr3jYn1eLwWzdsayHyyaT37cvG09fQG
ZVFKfpH9JBvAVrpaDaqHNY0V/D9uBR5x8t7STWdbTApJLAwSDJY3zc7w2v9GAfBg
2N2/BgyHQpRMkXU3hqXAAQlPn2i/d73zVlxZRvjaOeWXoEn2sW3vZ3JCYCJbf7Bv
XUDxtJfjMEaJfRNjwSYJpHASaRVe+1/8Om1TNnPmCnhMG24IXPU56AHkbbzI4v5p
cGmMa+jxcJQeFFOmZ4E9b5+J5Wo/PlU2d5UmfQCQNGrEgnv3ECY52ihIRdy7j/mc
WG6jhu/M23qD+Bm4ezYamY15Asqi19/dwA0N/jYmj56CPA2q25CzpN2feT+goXPU
rcv9S8RL1YwtbCi5bH62XYX+Fws1vxB0rky9KHxf3PdRq6iQAMLaJeWIbfYv9xnK
NP9uRrQiMVMgFEAPSjZKTjZQo2Ndw7+71Um2ILDO3PNAf/IcGRfFJemkfFsUqbsX
LNWxvwrVPYQowhFDKpY02563W+yS4EEidviEG6x3AIJl8NwKn3f4+5KlOaKALwsc
IzmJTmGFKAv9Pc7BNPtk1DR3lIZY+YrHwTKf83kfACTSwYMu+0SrFvxdo+cV8t03
J2qZtFv8eW4P0dAUd0Cs51CwQwNPJC2F58fqmBIxJRgwUzLxKoqpuEfUxbB2RMy4
jpFDULosUMfGWZ+SYpOi0CoZ9YKwFwQX/6Lo952naqAot/2GAG7yr/5SVMgd0H5E
yEvUtDwSPr2nVjGwkO1lw3nlDCNX6+diLN+CUNnCSorsghgTs+MaM0iDdRRi4Fdl
gOG+gxMqVoSLuUz+KW22fPupy/xFQH4YdfQr0WTffG+hpGKLRRICs0XftTrqN3B8
rOQVMY9B61CmRqYaQC6PrI/g6UXgnt8pK9j9hX2V1HlgOSI9l8zoOBs2YwJgGYLz
Rr0s2iJOOb9KunmYvqpdct9bDduH1NZmxgAx5PCJ7QRmLTWda9DWkf+ehe65QeZs
0EQ6H24r2BfxLMCt1BM+fYi6jbxLqzyhPj0Q7hlaihmxa/EkIInc3qNhRcJmP4eG
u/dwlbOC9WPhQYM+ArGuejuL3O2pzwEQJWMzDQOOcPEgZ1+SI6emkGBXDwpY20NO
IfsHdJZZdDkgVO70YTAmpoMZNaBnIO5/WatiVxxsnbdRIlo9m8x9GUs3RuRYA2m8
3GOBNXCHtUW/2Am+dhffloCsbofvGP+ocxv6Q3AxN8hx8Z6kOT1beOo1svuwoghN
9RjVEJoloNkbh48fRVRJWwasl1jMQ1PZZiBROgnEEinZfaD2XZUqnDxvYLlOfRPd
dcnlnuKAWszRlbZKejOBWq9LCq1a9q+Yq71XdRPOD0O6hXJ0R730lecJvV54m0GP
V2ZaDxawfrwcN35i71YsSeZE5S0EPq8DIWDJKw23DYmv/UdSyF/L+LxvNmtR8Lpd
1iRe4rmSf/EVb6iixzpoq/ieThYP+s5s/WTNONZ6ts+HmlGT1jigcSgN5duO+9Wp
pp4Fb0r4DPx1MkPyBsMEBhkjVNc16keRclvWgLxaAZXWRV+e/c907+xOO07B2klY
t0VUVWp3U/ZoxlxOQRoYVVPmXrSMJ3iYYjJmYzhREDqngMmBABNH2iEHcmzt846L
HhTyJLytYkzVcLoLfbXX6Jxck33qUo/Iy6XEteUdagJG/MqR5ZWU6csJBB40tU4E
y9O34u0vDeKBaJWzG7fqCQBC2IvvFVaIi2BdmDRRR8JCvcWhfVrJWCoB+b/rXczM
A5j5mb4JAp0jPlAtpcS0y9eqwBan/M/LRI0BihRv5zx1XIz41oux4V4ZO5PD2rD9
JL3iuJylu6kpIeW3+USsKWtcMFWDfL8mzFm8e/M6ePp69IcqGAHjBSNLuNNP3/dy
RmkOBe/bzMy5OUwkdfivE3uGR48u32efoTHp/YTYEcXRPMpsVf36q4715ki30h/A
XWI77MY0oKExjVl3r9IVYfIgMOticyi1Rs7Q3Yl9VY2TLEIC2CIDzYsr5UJgh2xt
ymcUvM+6ntOt0u0BQOgVMX4s+zmYiSdsAKkfeY0Wsa3BYmO+tejPQxJPzBmjdBz5
HK91lyXUFcys4xCL1zgLbaltyB/yo739OO2LT2f/jyFwtWeO+eqgkh8NWZQDOoHn
BRp+9XndwTv8SZzS0skjuybNpUPpR7SZCBPW94LXCE2eugfPbFtDCFnmjganNHqr
B0Cp21GH+nHi4vjWyxiERnFEkOSUysMgWl0g+WQ33BJHGT4kZSPadj5C+e4R3DxS
Jte56h4qTtsmCIlcLLNXi4bESZDW2dP1YFfpGFs5l6klmaqjrSTbQiAPywutNI7w
JNLJhpe5MBy43iMTHnxgqfuODP6EJxC+pSV/+x3mjMytRTsVXmDfxIf07OyZ/VXf
HzWjo8a9twNy9Z1WEt8TQ1dcsblcHYq/hcYEvMwK/Lb2L4Uz5H96OSvl4XnZmnYd
6KVNFoUogk3w8HV5bZIf89jnKIr+t/wStfAqTyB9OdO7ajcArteZcWKkXk62aR2N
zz+QWRk6VEJs7XkzPGvUQBCXslR6pHQwTB4sS7Kj4wQUcs4NrTLzKys+JLI5M1AL
FqCMX7+SdIzHt426F3PRM+TnEzoCld1IqSwWwBrsw0rZ74IUu4irhsPzAKpElEAz
r0A8vlri1MGQYl27painSuGZ9mT4bqS1VCV1iLwqWFA5WG8+GIeDGtJuKAk18n9L
IEES/15w4ALRPjqRzaWtTEKKcbwLMBqlwDLq5e5YD8UPjnAPnOI1aJpAzgEVptV6
NKdsk7UsO8u3/W8MuTzECyzAMbyQp70tt6+fUKM4a4ZLThyhVLDvVvXdyD2+dn34
X0Ze5e+A8GLEk2eiecUg92Q7oZFh/PEiWEg1Btr9+cb8Q7UeQ00Y95jHeU7aiS9a
CPxqZMyxvVTyubuTITXgVaaklXCUyfTcroxD4jMo7LqRydmDbt73hQzcY4qaFWBM
XtlwjwC8MR9UbV/XM1N0VhIzNSzreFDGT9gsN9Zx5BbUhRGbop04l1R9rHRHoebr
niCSloAxb+NzBRMPTX/SxRZa3ddPnQVIDAw6dvlHmOAsmbGSX6VE+4fUjsu/upcj
ZHfHBvgvzMSU0Kqm8BwO7YHisB9Z0ls6D8GX6g8JTqLdCYumC1dxooVcPp8KUO4Q
yzgFYuNctmRro7sN3f8vuq+KuHVvZBlJkoNckKxcYainzHPiUGPKpvXaiO+aOCyg
PP+F0i6iaCbgd8RqhDxkuCeL0BOLm01u9M4VSFDzt1/l2bgd4jvqZlwuWTPFJfo+
612+J2odwdMnzHwbxFPXEzHHyBceukGCufcNMFT46p0YbJBupiowwzBGKuWtgxaw
EHEN19a+RKMpvrqCJzEwnNRvApMexI3mM8MLyOKTnetSo4yZdX7tVAnI8DBDdxmt
7u6LLUas1/+Tz3BYLjvOFq0nA5UW8dNP+1tmE3Ac8NAcPTC4Ny8u/azpIPip+8SL
yD4bjN6zeVj6X3ah/pnZ0tjJJDAJfLTu0N72jiN2ITMVqT+GKcVHvBhyoK2d/CHN
mi4DCUNm49PTwSp+P7y907wErxCwFvknjmE25NIeb2yX8vAOJp1PjtEySthldk6c
Xw6lDb2TpmKP4oUab9wVEI85TvNdqri4dKyjPeT5jmLiVYra+HNUUzIQyuDBA+Hm
28tkDmpwxy8WeJFvmcMl8b/11+IgRuKZcrFMHUrvYFxA4eKmfa2+Ivloos//edOb
sq/4EvQLuRExspSYkM6aUbYdhtdIsjML4BnDyLfcB4sh0V+ikFNeOeR1Dzjtezg1
82XSJnXjvfO5bUg7gI12WFzNCsgwfZPBWfSmpvcGexitKZ7lNx8tszRBLw52xyQ7
eQBREai/KVh1yVtU7+pL5rfl8mPuNVvzaY4IMCTCELKZX2Oh/JhVIFq8lpXC3HJD
86IYd4c0q1pbsQAz47IuG5u31fB9oe7dQPAlUp2nYLJKkMvEkSHoT5jQ0cotdd7u
nDdgIL75kCiDz7K9ENpmgnLd7Rm54kztwxp4ELLYveg2Tn74d6ao1jgZ4mIUmUpE
ST/GY7CQyOnZhaXYbutugKkNvyBzmS5aHzw85K3P0luSd4sQRBA1CNQOY4U82GJY
dYPdBx2J93wFYjRgwnsadS9JHODBXJfXgCrPe1zDzcuQCSYZrnE3AYV+yuNDy7eU
uahy+djNtPMNdttieGRy719QfsVptVYppWkx4JW0I27VBGISgGkzNjeNTtRl1oxf
Xcv01ir00vXNJuv1UgAAgbLaGGB+6WGFKN2bp+Qcke4+06nCJDduDoCHa4WH8P0R
a6j8LN3tgnVzVGn6eLClqHaEByfQGlNmZ/inCqz+jdpy7rq4X8j9InEqHFWYeCh4
LRu6f2oqlF8hbiapMG+uO1slChLi5IVF9Dun+okhsA+1mrYCp+aosUSGb4d0a80d
bL1kGsuQaaKDheLZfZEHx85Gaf32lTD/lIkfOd2fsQjbKj5bq7L93HlFIXNWbTVP
c7zgNr29I0Bw0wWxczgkX6PNAWVZgeP03jeYkp6HKodyxbfN7fuSf45YPrcK69Uq
CZgpXwXgJqEjPCX+arlpdmDaBDVRnmXV+7KxSbd6p0pykkAt/3Ab2NfJw/Fx1rsM
Jk5QzlIBC4sQ55wflRiDXxpKWlCsXadCWorKiRXGM5EBRlXmUyXT+haCiANChPLD
qGc1RRJ3An9TDvtEaqWu8E1O6IjE7lo/HMxas8CoDb3A/GHukWTOP8OL8UyIA2pu
qlHZHL6Pk0eTYWuUsRIbMze+M+IPneplrn1KNCdX8UidkveZ14w7lRkdEKD0dpP8
yqKLuxLrncim3V/Xt82nK7BsWZ3Zcp+/sIacI0NdVLU9MnJxRbUmy/DhYevofGGh
GFP19Jn34nAAXQv1HnvDEWXEPyb+Jsl4Tukr/JBPG0DSTeIz2e5OIxYb0+SpAXKi
XXTtI2KQGD1t5SidUf0TYc0PD895dwSNrbu7RRzzC6/yp+7+QAGBVW66w+q41TRk
t9U60THoAbsp86Avi0XaiaFQ1MO0uFnyhIjFyAgcLFFslYf7DFJg3d0+dZpddVL7
5eok1xac/Nm3FPuVMzIm/XnVUvFpdWCO4oj0rlon5e2coBVGpzRHMZ+gQ4eNawmj
29VZpmAySdusHdrPHy+dIOFeWee/ZKvDelkOSd1xKuDMeZvC2G6u5o5zkUnIp5fB
072bQyC2+cnIf/wy4lfkk7iduAp0cweb2nQZlWwd3LSdSQpJipd3AX+0hiRcVZwB
20X8qRYZv9U6m0BaBkE6ACTvtzjaGDTsxYbAUDiKSpk3g/St2O2AQpUQfkV+AWqg
H1Jbk1iqPdlCGpzryKrm49GqbUslvjf0IQnOgEkcUI0DbT7eMlxWg0mBwx7AplOq
xZt9vNFvWMPSSGXWsrav0xfkqCpWjsM/DGukvgtTtdDevSS+b+wLr3BsldNiZGUC
FYPV4gUtYgxNsAkrDmYVooUnGD8Nb/jOz84x0xyfBpwaLIZ4N/Kb2XlYYWDIkXo5
ZBpFJDlInaPvSdW+7xEZ6xJ0WgCUpJGeOzP8JUUINMTWwUy0Vbj8r14GCipdjvfi
kuwSMXShk82DEN3gtga0322aZcl2zx72Xulo/aD7KjvGOO885vkTt0s0OkbAOTxS
Kpb5VtEjbt7J3CxUBmxasmc8fBgPElistw+jRaiuWefUTTBBxrvK6rD5YOZRlJ4B
ZF+lWxRZ3jxzO3Yp5NJk1qn/4sRCL39mzVlwWHmkiDLQbDzoGclhmh9O7XnJ4oZr
KuMEIu0MbjmqwthDbqB3h3PQet7vxBmYtO1ZCPVXT7cqyV063f3rsaMY33+8Dz2W
rnfZS56xAdrGE14NX3trEKeWJqty/AH8WFMYrfPDrp6lFfVFmHTdA22auOgCXFuv
Y8ZbqB4RPjZcpT6d40xEuJjqKqlC1+vn4PcSLYSe2MsJotSP35e2i8BR+Z3b2PIu
5RKFeapIyklFY1ATTbG8n0v105ATQB+JieeS7aDHl2hohQW+SFitbfSEI1UAArJP
/MscbcZ7C6rxWdlB4ZBkG4bOqKqUIk0Xb1U/jNQTSnEZZX0i88/1o2RrqoHje+IQ
SWEOY4YT6PnyZIcUvMtW+dRUYqhhCZqtUb1M66tqOEmhwh1nQiaKd0EDoNSuLowC
2An4z55lp/XAg2ldPygyhI8E19VtTvm8hEmpGMrl4F7Pzrhioj3FXL6BoFsql71J
mLR+YKpL85phO7onJPmA1ILYni25jE9E+A5JTRyY4W8u83TBm6zFbWwS826WsRs6
0X6EVr1Llp9prJFeI7iIsQ1E2auWEOx0LWIcYxfNBKhxsRwrRVOO7S8fcDlZYHCl
7Dzm+aTVroi//uUo9oLNg80OulUPk5Yus+ZjK4U8YWcACfATO5xH0wCPCRyE7YJE
SjrgNll1EcoCAd97dEhX6EshR80L/wUgPKgHRcVhQUpIjez5NHc1kTa/C4Hk6EbX
t4eyiuUWessmloAEyMGiGDpiPMh3/A4EdQiKKHXHIxZvz1+hFi+ZkKfV7o+J2DkQ
AWJ/9YxeIN11lcWSIAxF3/gF7QKbO5/f0IYh82TbP7nX4D/eBnzYcCCeXLryvPTS
M0fnXUSCShmKRw/J20/OKTLTQ+wpmNa8K7DVYeP6D6mR4Xzh2iDLKPkVFcEgKTB3
fB4/WIL0e+lmdyK+9i46Hhr4W0MpiPDpytrW2qccQjDZ029qZCc+bE7uv6yF5Dyr
onEHljt6UjHywot6kILsj5U5TiOo/maMmlmo21NfVg5vCH7rKICU/wh1XDHmRlju
waGuZV9ZVRksXs6nEeVECASBIg6BKar9VCcnoENx+RbVKtUF35ymVsqEU1+08oF3
8lM/0XKF5qHNYYZhi+gikYR5YPBDwI0D8IYmMG409Me0te1F6FDNT4DieO3o8tEK
Rox1B5g0MSsLcrAFgoZ1G7m41WgYRb4bc2ntv2n48A/9KiKF5/jaLqXBIOVhEw8Z
wHUv3Yyddk2sR2JNqjTSDt5sBM3PTqqsH6JB0PnLSnD4cp5Mg22z72BRRU2jCobI
krD964KmNegVb+Sr0xoqHxprM6ukhC8CqVhudWGBoVXFKnAERNaCc3i0hWvEcKka
qqNqeekhcWBFZi2xLRDy1SU61YsxfuRemkE0zeDcZWDVkrDbs91CaU3NvSOYjtLK
XCFb/C9AnK+Ys8LpgkbPiq+M3O2tIQv1tN19pXz4205tahxE5nn7UdZYGSZdxA/y
8azNTKXzX3bbsXGVtnWPc2gWFTG88yUgZENeTW8qkeoc7T3aR07N4VjODIJmOv6o
Ht0rchNatP/NzHYFoc+3N9diqiraheJJKbDIagf43XgnKD/sfKMG5pOkM/m4DmKh
fpPo4OhJ5mBsa5OjJtGlOEaxROBcFA/QmzCjC4bTc4jbBUxBcGfP2zM4AQnknDDm
KFFxL+INyRQtGIYLDHK/xLZQYXFPNV5nOsXMipkyf2OGs/HQtgLAsSR6CkilZ24V
kdVrZa/b/Te29k9XO/2v8Iz6qAJdMGz4s7Z/y3vs5SrDTA4fMeI4g506dZmerzC9
saD7yqpnfVDD3D3blZD8FJ1MNZkiLmomJAAFi8JnFEPlIx8k87wBotGX8as/Mc0u
i15cVDVAX0hly9nmoUmPEWGBXGVcn8lTBwkzNqmkhSokGYNFJOgJ+JS0lF2BPkk5
hg5b9sPnKwaIH06pTs2xpGOdNiefuW/zze532zW8gjVVnkdN5oce/i1Cb7V3q4yq
rRWwHnZ5hoQHcs7hmGx//2aD/5yi7kobkOIjMonXQ8/qh/F0FuUNRIHkQAQKtcox
AZW9HeNpwiTBk6RJ59CmHQnrdhq+9k5HYON275WaFtXmdPb7SmQ5nO+2vuZLNMMi
iz0NTNg+rCDpHrvsOcXOcqYmU78thQ/M1XgXI8htuY3MRmDOFpEp26+Gaavt/0My
zNfZPxXb6FLWVVmKNnmzXxVZmctKvx8Yzvpg8EkQQVrH/LkGmJaorwXQfHzpTIXo
S/QUVCtywIjriIP+/E1XwnX19Mp+RXWKCUQd1wTg2iQVMtX+xUunXMJMD0CrZwHe
IzexWAGpcuqWbTRO6XUKiU+BkBu4ZQaVqRcTWvvIzw6FX8UyEPdCIiViGOhyKqmy
6rXbcl4uy7XIdCFpQf7ATAc1Etp4kAoj3K2e5dQy3mEtxiqrdBpswmkIy/yp6IZr
Nd12FsD/cW+Za+FbbVkv9/awo1tlWulFfid/J2EBMmn+f9QVko6IqXRZ8gsTI/bT
wxnIJRs+XMxkp3qGBpqJRd7/wzA2D5/wsNWX4cBalG4epSU5QiYlwsYnts61UWPl
t3iMn8mshusls/Ca6X2HRnkmqMrr8pOTvReApFDwXGWhYDJeyHjDI4ZgMYbLGS2G
T1OQ4aeq5TQ8Pq9Fhs9nDVDwET0wE4ylK+MyimGh0Y0TGXUeZZhr74aBvz5cUdbE
3Znou/BtHil/TGqVK+KkJtvSVg6XGYl8/1og33BDUFPcVUFJ++TfXKY/ad/Ivmyc
HIaJ7ojRx/40H2mW9f2fOTKi5SZGLnzzxOjvjQpejz/Skh5sa+MjF/JGCKUn3WZs
8MPJOwWNYauezqf3o7kyHBX+OHPxSDtEY/Xfg+0QNJLZm+soL+HOY34EwV2Tp5jh
4wkVOqm7Sii/JZJeNrn9WCVvPIkj9ofHt4f0SaLyu5HONNyQLTxIuRbJx0nAjA3L
pp97AUAtlGKYLTEZycjmmllaLIGRL7KGn5/EkhKqHsqj4KJMUjDMWjPREq79dL+S
gQKPOVNfMn7gUyT23z8+EK18Zss/o3CSKX7413RyhxlimtO3i+V5JSZ3TvuvCnBl
Bx+y0LBVE2Slk181oGIWC3oglY24Di1PdP9zzmzK5irUGDNw6YlOkURVazBkGKW+
gWDvoJBnajeb/Sdx5WD5LAIpGJ3gKnos4lkG70A96ZRdK7jOuaebxQfL4tc4DRn8
mlbr1Dm0JgHeDuf0hTNPtuwyXChs3osG+PEADHJvMIUGvdqhrqFgenrlyLrOA4Eb
lH0mQ7p6k0ANaYaoYyFUS1IutNDoi1VBZwNN2I5KOjkdyROCE1ozdx7V/XMnBnxx
ww6cTBDcgKZRfElrAvXLs5L6mShFbgItmvOcStxBgdhb3kaydiW0vsKdEUGgSgNP
dKMzjTpmEbhJG+YE4e/EluyN2Qm6xUvyqB9culAUonhE2vIH/LdS5qGwepucCOHa
QKCcNiuuBmI0isx4wH82IxnUAgyLr9Y2b1cB85p7AROhlvVSVSAZ4b1eocFfWdj8
7Z76f4yrNvlXQTUN/qx20iMXgO6jqAOFA+3Is+owa818ffdJYLaeJf2HyFfPj9g+
mUI933WO09yhBwAZk+yY9tqwEyNqCt95XXgunh00ykXayjUBc78xJqJkf3+3cXdv
zRTOBk+FtsIkLp0/IMDYKBYT3Wq4VeykY8tI+KCG8rsdmVrhtTdONvcsfbtFxmGW
hhiVJqIBaiK3dj0YdO7nSGJpqui98kFdqrjygm393agDmPXtwu6oJ2UHVN5oY7O7
s6l1eVNG/FL9FQUWr2jVkqBFg/lEPO+pKj9i9vWpIXmAKy/VXasgmSd6/lavcOnV
9PDveF9E9JywhBjwwnlwqF2otmLqC7Hlc8gnlKgexVPfeQt3sgMaWR5FF7Pp5DBZ
Ij0YPOx2N3Ykt98IivG9s/ujCbTHzRbWmpJJf3s8jU210MSJROraAYlINvW3eGOy
YKxH9dB9kx0lyrjj0kFLZ9U//iru/5y7iDPKGLOGBBsfMTRu51dimUNfMCKNWYNE
am/Tbveg1o0BSUdCR+y5fvbp86I4kKmbBWpfvxr2JAruNs16veXL2tqfuFaKLNiq
qWk2kjTvx27r1uWymTWi/16EZcaijq7eM1mA/Ixz+lfttyTFY4cJu1V1ZoOXOXZS
T2BMycCt5ZT/aP9TpUBBO3OZiaa5ztiDrFq8LBUbeAKrKbhwCmkVmwCDnFszyIxi
pnnXT9YxSX9RmTa8DwQEE5dK85ukUy7zwvKrpHYj5kJkAvkKouDFFZ82KoD3rwjq
MXUSiqomPtfBUlhXZ8Vi1hpw05HNEaW3aowxS+xS8n30bBxTn8bTua42dspzCEq3
dP0zhScz/2ujUAwCDmPcfGDFYvfyLLp26J2MYKm4Q0LqIXclRhbJ7YTgbydApq3r
Rf7Typ2G9IlCiKnkGn4Y6Lwm8R4eSIHIRYUs7EGZfPLrJfybiSqbRnKx4aeZNrI2
4rfUB5ycNwsd7M7vWIfVmsMW/7ddWJHqtJofY7I/Nz4vlzReYG1fBFcOKS5Qr3oz
p7QtBjZoymZV7aks9WgYyGtiWVxVGCnnlnrfGQX9InUQjgAdpv4d2i5QHF9zp+Bm
tpsabR1lBHgM6HV5dvA/AQ3roZolm7R8NSyxVH6ZRCdmtNX/WbM1qJBTzU4m1F7Z
tEHssokqkDFl8UXcLD5DQSBg2YJ2gzdjv0aQXmg3Ntqw2kMU2XG84anoTaqCAK8G
l0D4yoHoabaoUrzPOoQP9BpVs2RurUB3/J5qXc52TxL70KfvQsl3rqM4mQzzfUwL
O/ZmiwAzkmzv6IKQ02OC6YQGZpufIq/0szBwaSnqFvyNEEuOoBlntaKLaEjm9nY/
I1hCZcTq2ciVgkQxOh3/sLfGdI2U01i+KGITba1fcjoUWnTaVm0YSxhtYXybmzCF
6gQ5IFDQlPrS3rTFj7/8LDBz6JkRC0aD/Nr+6WYKoJ4NSspEGbsGgOvYNdQd6sfg
c0KzV0KF8lBptXwysz+ez73skMKVJC9YwgqhAw+fHgZ4hWT8mnirgsXMW0m4UnUg
QY7l/WUCqs1PSSR4NcjmJmZ68zyfubNDt4Og8KiQGxPI+P+9K2RHHRp6dZAQ+7q8
uR2OQgdJGBO0ZtSO9BkibdwYDT1esB6E3rnlTGI65pxMpb41i9iprVHEMKFsHlej
BvYf8R64zNBlddz68TM08O4zPQq2J+pZy2JrV3q02w1Cg8mtDcwP012A3PeEjv+J
p1vhtT0J8ltAp/RsLgpJu9txkM43lQlEmuIncq1P7UJ/1VtK5n8irwAB+FjbNURZ
UHm5tgYqEFg14NpLKIoZF08OWTEBkKEdCRTvpOvbGX7K9NBVFLJ0oSDIhdZdME4S
WpB63tc+UaAb+iYGPMRVrlRYH6UV9CdWikmwyYuD6O0sW9Pc3Ycpnt0dGmz+Bi8W
xfp8MgEn4v/fxi0VKw7FDbqK3o+MHQcWBj1CbW6zEGrGhIoDn3NR+QuJEKoBQ0sf
ruHYM2DkXXVaBiLQnpVj4ut153C3ZirGLCk3T5O1ZKO5u3fvKpNjxmeDZEcfUX6/
+aufpbhmsWuCLfQDofVl9I9PypTlkUauvt87EEWc4QjdoCYaXClEIbfa5mYJX0QG
NQYpyhDmNT75wP54BgUx3B8igVK0V4oj5EPQ/eyfqF2nOdvAUTBOMC4ssBIf4OYx
uHvTtPLGxQLaydQdywDfFVu+6i4+Kib6B0LXw0A5Z72N/o4jc2T9Aom2cNadLZGz
iYkJgU19SewgMD8Ijpnzwdkc3OYQ6DmxOxndkC84pt0qV5LjKkVyd6AGgFBIDrZc
O2G7axdimLMc/jxy89/Y01NfsI6yjxp0AyCIYGqy9CTkM5NqA9qNSqsqFUDfYkMj
hlbrgcF4qYADQ8E00NU+nqjwVyddY/MtdF2rDBGYbNjZ1PBJumihK4XBglK64Uq2
OkUMd+nmvTVBCG6MkTKAlov/jmGvU2SqXoM0Ip7+XPwAzJA1tn8ca6+dOU+a8XIp
hqgNtcP2ZKS+anHVxYEm6boa7xmtVHOqmjcHgJf/UReqX2C+2xQRM4WOopBJatRG
uu55nRMppSjGzbDzkIK2ftkPYnpsmKdJ9SPbmp6pu4Vc4hRdB+Z99ymwnKJV5skH
u0II2+tL+nfIq6HdhYJ1U4cUEesuivD5SMnppEOwGqFDf6tJCvJJx0175yrnW83v
8GxzKIyGMP6UfTmyFSG61g8C5tOYYDzyzfaZr/9+xoOX+tcyzFnJICd/fjuQ+owf
8hegXGTY6WNZUdL/hjyhth1FzUak0HjQZF67GN5qYb3wRp5LYOy/+lAU7Q9NEUKL
hy1dt/f27S5a7hzdvbqrynAfYz6OgUC8kLBfYLL0iHiSy2Lc800WL+wy4rDSs4dT
gkF3vUqEItUcvb5Nv9LkW6SrJ5LngLON2iiffqj+aKWY/+eIt7azuRUxWWeqRCMZ
Unu7PyRy2Ohj+WD5I0dmOk/g343vL8Ccne/MCacDMetUhPtkR6qfpF1jGLACjhhB
4QcwCAkVojFEDZSWQk62D7n5wquPaaIQfA8NwhS+iHj3n+cOCtmDLjdtJ4Ex05Oq
4BHTONN8DBMhcJGrnriPBF5Di3Z8tMG3hW33ZxLIDM2buZdQfZadu16g3Jkn67Dk
YAHV+RCMOGQ4qz7Plrdt4BZtPfFylecqtzNSeypXa+1cpwAIKqk/F0JcVzvxrcNf
ohmP6PuHNSZtGAyA6lxkYWcqBaMsXRkzupj9xvFUIyn59pspJjN6mSpDXOI7lxEs
lBInHyCRetW3CUT/YC42RI8abYDK67zvyq2fc00CZfxy1nkx8FHhBWbkF2A+91yx
+P13M20Vu2bgPJ6XCHP1cUtOMsA5B4Njy7OoUGOVoz2q2UaqwDTG4GPc73oCjJZ7
Jmkowo4zM3pM3XBdSDoGGMuB0pt3Lb9NNIvYYmjwYd+V4qhy/6DNtYKipjVBANR+
vhjPe17USi8/73o2cLqDLE6cfjzap5cTGcGi8uOEdubxQ3eUPwzuNk72VNxuc3oZ
spNelSZFU6G93mi19a+GEkdURU2Fye2ANcwm3Z6TK6hRypGhXh4U8sT8C3IQpQaf
srHQJo4oh+CmT4wJemAGskL7ZmP7Ss8T46cyj0qb5RwheExPVr9B0K2QNaHmGrYN
WWXL2YzQO1Labfkf0oDyiZuHoCpmp0cddCrOgDPeS/LVe0afVzgJ2q8U8TfG5au+
ydxMqXGmfuMCrFfLio0y0xuuoZ0U0C7IG6ux8Bqu9F1GGeMIOifzKm/BSmXloDAC
ZWL3Hg6MeiyvoyyYCyyG894x/KbMW3N5EyW51uN16uvgrs2IzTY+C8ckPcOkioi2
iE7tqN/+LPw0XJ+TK2jPG4lRCs7W1NYxw2XbrN+eD+sHb8pGTjNlJ1O7EIQuPsSm
fHXa+Xu+bpwe7Dj83k/OAZEQnZtlFlihg3JQ8CMkPX+GpdHqgDIxSgpmyehdaSCg
oeVF3bVk2JRdBGlLhtOhvO6vHbxDQpw08THj9Zqa1uEVbeWne/ojh9exL2b5OsF5
sU2hhN9XMIocoBJg25VP9RU+uAL62iXDSS7GNk0dhtJyiyArpiA585zyNwLQ7oYO
2TYP9fxeEoBQdddw8chCqiOzFelfcTllBM8JLGD2UVxJzCCt540buWC4K3+B1aih
9sadW6uivfZoc8wR5ocPst46ndIzNVdiqnLxqGAK2ltwT/lNYReTkd7P2RbkSNiZ
42QBBG6gUsSt41/nCj0pjHpETvDmxFSVV/XYDIpaEo3aI36rHK8cc8r5IP9yOlQ1
DNiHhT+T+WjlhNibe87cT7amwdIGc/kk+QnSAaSBSAuXYZm2b1SleRrHBM703R1R
kUsHwfmMiZAqqHjCIzUUkX7W5m6euPkXw6xePyjYcVnDR7mTkymgIqK5dRFj4rUD
iLUNSaCxsSmhTb948fblQWS/3Sl/KvdefzPkcOHspPDCmIU6EEeVDqCtMq836UhJ
cGIGsa4o147D+oYFOP+OH3t8BnaGpUaorEERUU9dLDKuLCpGvrRXbzA7yuNYVNEU
WQ/9u36W7yolB52mPDivq8MgXQhfMpgSKrUqimvtseS8D2zzVs0db7zhXZPE1Agc
cNCxW/bDUbO+9XudfON21bHwX5NDSQNA2AJEMbdc/BUMiAqAkKXS4TEfj2/M4DtB
ZVvz9YzCCIaJ6omQK+FwzSXZlcmnK0kRerOTatlRv3vqHex6l8MeBkzUi0RuHjrV
NQKd654zUYBhx3eWTW+W4RfnCoa4me6qU7YBHtvdkI/E5FuCoqQavU2ATCvNyNPr
JzxQu56oOFsvvCfDhOCWamv8T5AnHWliapFO2hLbzXl0j8SC5Lu7RUZUtbJBLhgp
whzc3M6KiAnzLUmMbDGHtDZgmqW0SyUi2FfbyV9Hooe0pj8Gd4clxeV75lmVj1FK
4dKk9ZzjT8VAHJmGaUAx3344dNzA4km443coXdq3xk8jpQEAnEFd/T/uNvaznLKv
oIRtgF/3VhBwFvShjkDVZPwl5u2lo4+fX8AVJ2R8mw0nUrb0pLM3owSve+Ndpd94
g3UQMw0QDZedYdLeGudVqbmrnJNBB2A6IayROGjAIVU3Sw7o0hQo0CudFmkuoAo6
NvTxT8ILLyscwBTn6L5M4CKv7dv3Ijxfah65FwCiXJV6elIvptIcHhr752GO2XiG
U28c59YXfeFaKWmHsvkBL58totrv+CCahdhgKCuLICsy1OzLx122dS8LW6ku6ob4
BpjoGMfpsEX6KJKCkt85r4vHRXrasTDXdBLQM5rbJRe0hTVNPQcQCasZ10iiYnUu
JeT1BuMmF7WYMi4d7fb2+eLmv8EuNxmvAEUPCiAGdtabLSfMNyN8yFbNb3pK3Ti6
VsUCQ3KUXpbVfUv6UauLFvEIYJoUTu8p5u9USKkPn/Nn0r2JcCr7vwf+3pEZIVvO
xglePk+7TsCyjFFTlyye8w2iyaz4OdCEJZvXWpok0JjjE5zBqVMGL/mzd5e/i0AX
+krdMbwPUWkB0vbj4DvyHIfLEZvBhY+L5X3yvwGJoGjYiK+8+SyFplKzZLD8cxJZ
3dpgcKoHnhhQuUCZoXa94x7FMhTdRwTiXL9uiOykDcGvWojzr80LpfZ7bq2UIoX9
D8Jc+l+rTfxXOM6ObGVwpAd5DTcTCzdXvidYJphCIFstYEh7dRVYqkHltTt954QS
2ilzIS+pLLgTw9jwUmr0dlsHEP1qfOkuRpRRyujXuq/+zZ70Rk3eEO1xFBg1HzoV
4xEsWMC/vdvfVVgRPDBNfv4sei0Ym5QiZP6qtnIrOwejEeEDD40Z1wATUimPS1IS
9I/G50xy4quAkobE+YU76OFg2OwxPXIWq6QeyrI7gS06/UNnQGZkzBwEyfYD448a
biFHJ3W57pV/CRqJ4kIOqC9It1VKSQ7XJk0U82J+99kYo2gs5c1zxOTgxgyT2h5G
2V69pB9gnaNdMIaL4ZmVLJ5Bc0bOdO9ol58/Tug67pb+qF/T4EskhfFFgxVkq/ow
zMZQ1zRx/T7oz2DGjhIpRdyZWvK9Smvq6hTHOj+lmBco4RDPF5/nEPgOqLgbIk43
EWbzk1R+QcEX8dZMRkIeW4RWY4HaIivzoW9yMPHwFfmc+YwuAOQKXbJJladIHJ31
OqbCTY4E90Gvv2kQnFRn7t6CP7nZIcb5CmCHcy6kwKre+pqY2p620LDyU6lN328M
XDenpOhV7S9xLeqtV7eVHXkyKv0Fn9fuu7Y21jGpplu1eOUWYY0InQf4UelwNSaw
y7anqtxjCLxkWHmqj5QUNDVMSnX5yXjXX083KBt4rwpaFg0KjpXueWYX/xlG6Vxj
ghbLOdU4EJ8bkf8U81K2bkWcyTV4HHFa2zmRRG84BkBqwWcyXKhQrNphNDeJ2EM6
MlRTl9WkHlwg8RyHUdTXZCmGClX6241ZMJE27bQSSCV1yubvEDAsSXaHUD5+ppTm
ZuCpkEbS+cs8G4IgX2SDIdjTv9k2k7R1AxS4ryel18Bp91JfY4t85Y2YdfEv/QWg
TiYWi/bK30ISXx/uPc2DPS/ZAgBqzb2/bOXoWmfvoFB7dNUqlO79A6gt5HwfcW1/
XabEMNYezQ8dnBlkomFi/Km0kojuPM1xP1+tGcn8iNwF2RLSqJGOkI77hpAjORy+
8tuOoe9wsn7M7FqGO9zkThyDJ8R5YT7aVaPRIVQhB2Jej9vvy3pCvwAv1mFHH5bY
EjDznAavVGeCRWBuRQ8SZU5xFxToU4IW93nSevd4pyIulLm4jLBnD1TbVrCCsXy3
RlFusJw8+8MoQxdWhb6aMZOFlPj1FNxTtOtRMZxNYoXT47PysbDosapivsuwjvob
p6Snn8QeOfBqsPHCFEQyzum0Uh2M4iSDBKa/D4Om4Z7O7bd0/EipV4lBET1bsZgR
UygKgSKMdg4XUmFcjMD2AR7apx6NNlriTQXUHDeVt+j0HNLd8M3hoHLHDoi3dGvN
aFmcUFia1KMXGRC9mFgvx/nPZk0rCjZBmL9bINt3ajZ1R71kbB9kdij4dC/16QgR
uES90GICgabL6Ncc95NmfFyMmfh2IbC57hbYxTNXFCpFrd8FCgfiyigit4ReHp04
nhwwiSgXFXxGo8WumMAGGmoz6L9tXB5tkptbnVLvRFDfouhuLGlZftnERQBgvS47
UjyqkVT45QHliXa7t4EFYQr495CjKsguAoIm09JhDtRfMH6sGiS0txFbXGVO+e15
NbnsGTKDQp9HsnlsEOMCNVg0IkAd6UFmNEzova4jCB+edpr5VEQ5jUQwqTGuZfrc
LvAlb/cvxrGaJgAt9R2OTtshCC3TFwWj0GWLEZHFU9sUtb92grFeXpwqt41jav5Q
6IdfvvpJIimK6AWHPFcYaLwaCm5mUZV72CE0utix5klsFD7YKAGHhavdEA/UyI85
qpz8uCZA1/Jv1esJmDJfYSPrBH6L1zM1RqezoORdQqpxvSj0FrvCYuCgshDgTBKI
EhNTDp//z4WLJiH2vLIGTGC/wURZiSxPH7HfyDD2bAHnWzmRGSxvMvl7ae+xXBY1
00LPZD7rLrJBYzo4UM/FgdoSMyQ2pbibL4jp7PG1Ogxr06aZE3jzYF57IkDq3x8W
g6ZNKWCKR7jn5RfgLFBSdGdp9pfuO22j+67p0eZdZs+cnj0MI3VMlW1Y7r19KxuF
GemzCfiNHEr3fsCNWt8IHn8MUXNqp5YmZw2dJvrs9lLCE843md+gCMFQAXMS2FhV
80PduJuNzTPQ8fiCDmkbdW5VBLj9q/cgG/CdYNA5cQpH8TmXyfr+dX3ShmfnehJO
bUmD0teW2DfmWrONOpi846aq4lNOgG1Q9nJBr6HtGkY1ODjrr6Rd4VTxyTCzzsvf
rxvYGhvnyJpWNYACyRX6eImmwVbI3dUxupl9/i8Q+OctGMmL4/Rf87mi+GNMcrnf
bVu6ReAy0ZRMxt+d0b6TvFWZqSP7oGgIcX9VLFF/j8WLMY5z1r1wOesegfr2Zr7g
cz0DxFQeByhXmNiJKRn9wNCrmChJc2e4Nup+uRQXM6uNMMc1dr2c47OdCqFMCf5f
3GB2mXBgsIXp/7JT4AHTrhP1wipuSb3ycOiVWaL7R6Cuq32ooLCaCnNGbD9Q7XXk
1KhjO6zbkSKLUZHMLzB0D1js5o/eCPIdUmcnjiDiNvVQRh5Qwgj+vFXiXCrFmrmI
VYDjzNmivNXBqYXisELRLz3Xak0ftI7ZCqWHfVE3K0tMshzosJxEoftl8/ZDKTWV
V3/MyTP32DEHwe1OlR90tgAoXGoEQ3SKRO5qKtGlolZU3BABThIa6ImNXqNzSc7l
LKiQTvkll5Vy3nFC9cqEeJ3+EQan1JYNRotVbWnMDkQk3JFSI2OMocuqmosCLhY5
mhu6nSwhUKqezRyUvMsaSU9jQ5YgJ275k/XNrIGfwyujuCsfkxZPmeT4RqBgwTRI
Q4UgCxDflzKQSFmCpFHtcsXgnx2f6N4Mtwr075hLVoRXdeN+BhB9DKiFtJGxDTfO
utuLlUorIxUZySvDPLEjJhSId/I9wzYPHXpvAsyGkSP1q8EeA6JbQRJ/XpEPCXhC
9YZ7Q7nZz/XdUCqZtaiHZGynZ2pPwZHG55bzPwLaZtqLfLzhQ5Covz9/3Wzt3FD4
oQ8qkdBm7KF0FZ/RFUAxft6zGK+NQE+GPtjVKgQMyFdPWQtZzYx9W2PQF/8VSkzI
PNNBjUjImDYgDTAl8wZw3QpGFGB0YZhkj4aHDcfF+y3A6BHvMoxdhCb+WQLZWHXL
GhCKCRy9rB8vbeOzQ90Vdyuirf536jPCOVmuoQkgJaaYtO85cuAQR6MMybnQIYx2
cjH9VNIrUACGqgmloKDfs7Bcm3CYAChsFxfvq3uVJFGKv6iDuUABjSYIFyqn8amd
hfOjLGd63UuYE1UuYyL6WZkFLo+HTt9DowkamwrmEqg1wb9hMFpL+miymmrr/lXR
HnlVFICHFMjWJg6YhVwN3ioh97Y07Tjhh4TG8kx795Ym+F6ROTJa4wuTG7W7pyuV
yNZ7NVpLlLwzKAI7nqDVeyWwLfMsjQrTIygzCds7cjaGSW/IZNtkzdIivuYMad3W
3XTlzFUgLRxI3j56rlAPrICpmAqCdYcxbrc9y8fS+0JV9IS6E0SmEzRIoNn5vvLE
`protect END_PROTECTED
