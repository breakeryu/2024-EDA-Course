`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZTsCCl+ILMtMuceuXmThW//Blu09/0iWMTRPiXAl/d1SYxpHJ2GTkBen7AqyXsL
jkxZOgoJCerUdD36oHHh/Q8V78RILmRA4MIS1l8hVRs2nM0Wb7Af9/wCYg80ShUY
cxA7sVcp9ybwFmTc3PcU14ZmAyreYIjBCs/Ij3q4V+Xq3JOw6dPvuynbf+q1qyb/
FkRMocBpu0gYSuPk+10FA0yKeOIJ4YcxnYjoQGPGJGOvCVdoM0ED/vOPjUcetWgN
8B4qQsPaNsrYFGKB/wX9FgTDZCijDb28RC4Yh1pyTSxvHfcoywU3DhvyIVDx9YA+
Wcbgi9ZHFpiSbTCgNdPlOId6xmAjW4ja6ygF8sIIPsvjIdwMLUU7ICJfPbJ0Xx4t
BlCXcB2YJuyF7f2M1MoGXnp74rIm8XObdnfYMa4nJIyzWG+mXm+vEv5D8nSRMRCo
i1wEgqZsod3Yhfp1hizov84H2gh5xrNhNBV3BjP2hJaHvzfqbo2tdtUzUSag8KnY
9P3jY4AY9O5W07mhElwZtIoosjy6GHroSIRgZyfJXWCvsaQnj0xPYVq/bMfcqX51
qiwcpibJahbmc7ip+UqvLEFWmX72b36uYl+lwPurijA=
`protect END_PROTECTED
