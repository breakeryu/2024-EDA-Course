`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5CsSbNTCiYxOULrC1juwCaMDomSTB38rZcFsQ4iY9qcRAiSfTslcgsEkWOVOp4j
t1CUrBCtNYEpRMzDQcqOGUKZ1gESx9I/K5D0bpi4n49YufusxFEOxQeDOnul0mKh
84Hd67HYsFCbTB7kI6DUtTfhASXNcBaDCHu7RABSQEXSHvnmS+eSa5V2YtV8r9De
cHLBfwNpTduiYXniJv2R9FoLJEBVcM1nsu4eKT2PJU8kK1bYcMggVUF7yHkefo9l
XS2y2e//bZHOxoGmYgW75Q5atLMPCji+k++MJXWaJnfbOzOfJ88sZbk89I2Epn0D
wGBuZEYan6XHP9bPbDvYu3WhXwJiLJDd5U3Xi7pUkdmc3fClql7XbdYwNJSkBRj2
MY+W+wSuACk5pZekOkFLfYwZIaH6T207SNVL01c/z3+jr0H4jW4EQQTshcwNzHMe
iNZ+TOsuQhybCIPQ/0TbXLCkk30IDBKOBnITiyno5Sy70wvTa6Pp1zAqjs1zfQS0
VEKC4AMDmdQluBtF7xpuIep5if9Tq/EtnVeEd+UvGdAit3L/FzShE2I0TslDb+qU
bSpZ4h5Ayuzb0xtsxxHDBWDfhq+9Hq7gJ2qcdZbFbkdIh2OU3Z8Mhy93CPqSk6jm
Vxo2vBWG5uadyrt/lV1Lyg9ZKZX1sHPmYvXhOZN9egpSkT3qUuID2sDCzxCNfytD
RcWtVk2e+PO5on5uHXPxrFTnbLUSbtmq/LQOp5vC7iAg+BrnXfoJ4QbGp0+2qk+8
RgIt7DLhDyRPnxHtcxMyrqz4PeG1DxP4CZNNJaiGVD/ZRgYuFJxeySgi6kBWKqyr
Y1UXSbbeIVTbPGbtkmseEXRLCoV+V1du+de2t+HH+Oejy/BtnMDgLF8e3S0oEyT7
Ab7XIdFB9YG9dGCA/kZ2POa7PXYUn24UN7uJMVWI4zsxmLlEjXYiM6XSZkg9Dy6U
2Fp4wwU2dxDP0CTNdYiZ2ygJZBpH+i9CT1HHjF25IdW7gtSDzOn3lk/2kabDGkVJ
5TgZQNcg47mEB+dHxA3Rntj3HZAIc4xBTDTf3yPeQ3iZjVc1H9hBqwUS5rDFm1hI
djq7HAgqigT8e72lK4hwGCeVTFPLQ37DMAUwI0c4iTEwY2KvYETPK2+x4xIKQQ+g
VVenKUNqth6MEL8zMkJgHj4SNX+RE/bZbGyhKLULbxVWK/V/xPr7ZSVcEuMuLHx4
aS7cqV/t66BeuLlTikTz5tyu4hUiRMqFS7bmfje/K/qjYphOvGpueU3fP2mDK5CT
Hk4J5JwEI4AET9fiHsN5WQyAACCrxx38te2QtTjYbTYxw0jPJUe6jRXGBuO7hb5m
okgMItQ0BXcFsnOLY6U77yQZRP71PE4ZfVLz7Ha1hd2TDu1XFzFsX0cFnhhOjciv
X9WVzlqmP3prvCbMCAxTXzT5Y2UF9rYeLMDY/jJpjDJr3VAKp2jOOD1MLbCE4g69
JiJZ5sBj8XyY4kDoC25XBgnEggkpL1aftG9dmommn8CASmtec5OyFyO78IXpJESf
2zAJAb8dP7L4J0h3VgsVoVFzUOzrqnNMCbsjugo0dbsXn6QxtJzxkFLsx7/77HUC
UFbJ2xlZlVQCRvyBsNPe+UaAnA01+pZica0t7LFsJKV9OzIDTkGCI9WPplpgMMEW
/9ghWir+kHtgbI6pYRtPZcb5DkCL/uxbV9oiBegiXy2olqkiqyQVkPMobvNgfzWL
xCeLtgkQYtRia6qIBsSE7vaX3gWHR9ImplLekHQ8RZnv71nE+vwbf1IuiX14L4kq
/2EwZm0D1CPFDeDWtRdM5lU6mfHwPTLBiMO1IMxNoWEBgOqp0rfh4qhn0bk3wJST
eimXRFBuqe0nA+iSCm/8q7Xq6d0WdB7C43yAAOK1mcJBNGIrJwPIbKks+jiTPIte
sXbeg1OHbW/9V/299UpC/fHnYlbtmoonEtfBJm/GzUPeucD65LqTWhPNaqYVn/kZ
ZWW8XA+x9/ll7LCo9EsKV2q1NS74/QEMYmutrZNyAjRW7LaBgKyqSzt+0sBbW6My
Lkj8VA1iqIMynyIxqAK5bcJWYfL1d+9JGbibCFtVihe8zPYXf1t4xNaq2E/6fizD
R3mHFGdReTeqywIYYZHPA9kaorl734dNpIZpcOlAO5gQTokkbp84ZHgjTywOPe4M
/oZTtQitGFEWNr4JEnavyJLSMg4hLAD4Z9Q7xIAEy2DVc/6PhtcUSD/6OBDA2VNr
ftsmDFHT0nojhuR58qxI+IVxzoKr+RpDHe591fHtLhYmQ7/f5UtTDDBwhEJ4jF+d
LHvPKRpzjUrFUIkOrkMtyOHtl5A1pxshRqbw64Xh+pM3F+yIevHNf2GgdDPaArHQ
ZHedIVivizATA+LzB1BBuuhWi4xnyRwABj/i7ZIh0AhcAZ03Kwp8g7p8EV1QvDnz
Znqm0rnMKXJHzl3woeP0i/xDrOI8f1YkNBZkW7pA64fiHu8CBb7ii8uWeGjJIRUl
UOWonbwqNt+IFFVuqqmVUdFXkH6pRJAiyQS5o3xCOhuE+N4OQgHRZpj3tVhH9Trk
I/DZikGwicnIiNJJmcLcj1unPyZ/I3O6EixrSuHRwskkPvSWIhPc3CtQxVpKjNPB
cnQOkKdB5wFBd3cKX7l9ZVt5GgirWU49PjTNKiP9AClBAaLN7cAimuSZgc/xocBn
wzOUKeHKmSWbQBTwF4PAQYs3/hF2Skl7mF6C2l+Y4PnkbjrpwWKCWnCBN3s4ZxWY
Zr37cbjg7jTBRRcqwpwdxddF6/+1+KNZwH1dSrGe1FoxJRbCj2dAYPYG6dkgAW5j
BXm9hV9FrhK4wQd6GZgJPpF5eJwFalrZeCykWtatY7aLYqyXI0VhGLbkD2Q1Mcgh
0F0Q6quvu/LxZj86NwIeGKJ1GXfLMJEMwEffbPdWcQRspAd9m3EEwaVmlopdTEoa
EmIKgprQYjUa/Dbh2NkF42raQ5pL2INhNSzbSLYD2PJXwym63Hk8NJP9TQiT0iUB
WiDYLDTtFNx0TAsjPaebQt2usCrhoCu8VjYw2wZyI9xgTULhZYhOfhesME6P4QMX
gtScl51Jf40oY7+MtVClK+OSrgZSlgPl8EsQ23KvC48lV1g1te5lszJKb2TBNJZz
qs5aEaghSLaeYVSLATBWXkpr6MQEPNsxVLlygWYIYN1gKuLyMsyoviBE5QBgE1pl
iFWnkMoifWDXxixiNd36EA7Nf/YRRcEEcFqqw9bJoSwSlorwydF8/nI90gaMFXaF
uFl2y00zQt9g9oFByWw881+rdt/tNGSSPHr7in1CNlcdXFRtoDRbdlv0EA6PHhw4
xOipKk7fUJNH+PX1FaNSV6eNAdEKGyQbid+LavfTUOiJ6eLtqSazai1TyD1MPf46
ezMv4h0y2jld8n0ok5vXKqRFtW+pGjMJIEowJ/yHSqMBeS3YrPciNs1IIuDJqsFc
Ce8dK5RFTt+FE+lEcdEB4kFUk5Kbh/v8QW5GPvwM9cb2I8G1Em6lODNdKEpWY+Jj
e7tiHL4tV1wIAlJi84rT5uWaRLLSevdV58yw4X7dObbBIazXrHoR7fSjr/AWTk74
/Xjk4h1QYr0WgmJGBhsXUIrIVYW+9LX4snuxSYhpfyknG0WQXEQizZJ+OY0wRDE0
7VAP/AolrPlBRycYyFmLcZ6rQP3M2H8/ciH6bS7nlrTf6LeQc+8/ckrMUxyrXrmG
pCChZPboWMBfcDMkANIy/oZqt2ZTQlMsuHqOuebjy5cuHSE5KO0XbUYvg1evJJId
p1z2Geg0L+0WBnAWWkxJ4Dd61Jb3esgTv9oLeGLlbpBr9CLlKGkHpNJ6yHZ0PTWD
dO13VnXIEeUIV4V/ZnCW2b2czcrC5X7JRXRt5fkqFdeUVSL+Jmu1upA1cIHZSrqm
IWaZRBEHKC7SYdm5gi9zNNaeSqaqEPJnJu8/h14mlsgiFswpXmGO5+yTYMSFKyGQ
CrBPNUMcOScNN7qZ96UsC05HUA40sdjLG4D/HWMzwrhLLu5p+nooQBYGXT3jRKCV
7V8LnsXw5xDCGSbu/PZ80zesC7SZ9otPsgxImJF6/aEJaXh+kAi7s9SNgUUhDDok
aIdGlEWx4mlYlYu//JpscDCH/TobD3aaCfXSLzqZpwqb5o2MBr1kNtZ57JoN/2Vw
ShChgQR+TbvM6bD1PaCUbBUl/iJuoEt/1xVWBYN5txJEwafmu5YtEouoNJfo3EUK
cD937gpsMKnpy3Tn04gVbfI+sA+jbEjPi8vEBVrRGg2yYvn6QZFYoT6zcmVb9yBx
/ksPX/wAerA6dyrkxXQ1z8aJGlmQ0C2gbOBaBZ3NXv5uRjsfkzH8neZGMJnLKXdx
FeJ3DR9THMUk7wPWHh977eJ5OBMnZyGgR3aQflG3NeucS9KWNwqiRu2o//WSEAPK
Q+ov3KNprAGt7gRRaxKdM2U7IKI398zSO2qtDKeWt5j2ClDk8R+StmaTK8yZ5p6F
jTW33I4ZogLCgunc0Ntk2iZoF7c0FB2rie2ngbmPQIE+HBBad1TyhGOazbIOPYrJ
QduyPS31LJpMfMakn4sGo2lOIkm2GEXLHk0PiFTRB0WGhob4hdAc76FznsJr1xWz
hyJ7W4KGdrg6pEwnStvgXkz8BgAbDJTGo76BlVG4UgdPbUJcAStVUzllmprKKnxV
RjYEBbmsxpPVPex96I9u7m4FJm8zBLye55gyez4lVKw1Rtkcj6H1ac3RuptQHr9m
0Gk8zMDe4hqPH4ZYCBEtuX6kZnv4NKVvzS6Zn7uxcn7nKMoIF3fuXjVaD+cyGoig
TmDLBel++jEgYJRxwL1xHmVIzBiSzNV/nvMbhTusPBvzEUtzP9ok9QtgujMuhQg5
gW2QW8mcr19yNzFWqN9oIN3OaFHyMSwUuQtit4T4NBNAYoJBAlP6sfs77rENOp8L
1+xYTEUv/hzzc6pa/71zo32Emk7siwOyvv3YfLTsK1ZBuS6++e5+DhV1ZZeOZxUN
1dOH1yJS5ZouLbr1ne1kRwHgzgsPhi90vYOwRc+ahGdJR+AN3/nDhxWFahX0m8xn
EzzzGH1PG54/RWDCqf2L3HSZkSym+LrBRvvA0mFG8ZjP8pZok921FkK7ZbZZtqEd
HRTCjYOFEIKqAUWkppfjqTKd3qQAjZddYnaPEIP7HlFaUTUm1T8ktLObMnihGzqZ
f23NMUv1YMdbKPUhuUay9Ua77eOdGDKcoE8HnaT1DUcSuuKZbfxpgALZ0lT8A2OX
qWs+xW1KLtZhxEAO9oHB4gJ9aJcBGqdX1DYm/IUxdkV+gpqFjHF3RAHupcJaD5m2
/PMBlo5/w0AbzG8wB+FXe3eL9GlVC1sNRhwIxo3yJw7C6a3cu/Q67HAG/5vDJ6CO
Y+abd5/9Ir3tU9DaGztlbJOq8eAw7ghCq+g7dpXS/60bD1tMagFDn2bgImPX0lTm
nEUAe1Y9z6UHD/DTKULokq9i+xllNQIZbjt15yt+yyVqwdL9OGbOYU0Uk3dmj3xy
YefTLdsQyNNlQ8bZmsyQZlRvmcJ5HvKfLCzSu+jM8g6y7xtOUlOuZcOinP8LKCWP
1sOl0vAU0CxCOT4f0UczbxCfNIeOsGO/2PmqEm3q2atx9vxslkRoqznQKJd2+JLF
6TyGZo1moxlE4gR3WPCup8QLkkIFXQLusVKaX8skMAkoWedjSY5JNuoKUmFz7WAf
RAJ+HhL7cUWMG690rR9+pIvomiBqC2W8Ss4ddKzK/OYTAy3Yqmho4KhUgWUqikCg
efR0mDia+VoQFymB4BnF7jQU5dalm5Z39l7ZZv2fHkOzjRKjXUJe6Ekv6vxEOIg1
DAlpUjQaGlAw/IcydQnE0yz/Ephdqb5Jf0MCcDJhGS77Q8oUYWoil2YUSPQW6PJl
dgzZ1hCI9efE3/+m9JU9mNtzSHSKjDFoZ3PENkXO9xAVMln/UAlvQ+hor5SXBYx0
PvJVJqLeU43D+8BoEt3CpQ1NgNNRhigmRG47kXje1Ctg3JJebgPg/hz+Z291zBDW
Vf//rP0U5Ywf3mTX4fNVGz62NTBryIrWWTqWyeVdFcN1yZEJfAV+6IgJXmiO7Roc
SGeDUuR0ud0J7fOs0Ljo9HjRlFvLvnlC0J3Y4Dr0bNlBCTWyyadSCFxC7l6v32pI
Ihn6oIXipZaOYn+cFASkn7QY4UpTdpbYVdf0Ae70wqfrNY4PFL63zoD2dBofIjzn
uYTDw6fvWfBNtTjYJTp5wZNQODEQub8Bny/KIW4JGrqcWXwmhrA0xQ7o2YIB26u/
Xgn3iM36I6tmoPx9+8ihPVzN9Gmw1ok++RWVqYC9l1B3Cb8OeY7coGjQZcd0BKAf
2nue1sfUmKcf/Cic35bMZZ88xRjgDX9EDrgtONlra0Z0Jx5XHRHhTvyAScc84moG
xaol9moAVyaUoB69J/HYnhf18+8CxfwKPcmO/lMFzTOMSpHR3yoOJ3x9bcWkYMKi
bXuQzUQdc/8SvtXfRmEiB/IjYebCqNwnEhyCO93xrqbuqsZxw3b5Bg8uwPrYWX69
x7Z9SZfJYHjLfH2rCHzg8NZ2CHJjW3PpOhhoE/a2egdciuM/T8K2N0a/APWozExU
eIYSUkDKckBdB1uMas3BVfliFb/9UhbeKHG41Lbr0q7C1WCaCP7tBzn1gaFOGUby
vPfEIN7flpsp9fjbWnq/kRbDRYlp3DHbWFIKT0wJ2V+Ei2rBNsKPk6DGUvx9PxrT
Hg8K7Ku7W1VPwXQPmfuKxB355swGe9qVWjpxMYfXjTY78FGr6WBj9+g1hRU7ybjB
d1axAi0TqE0t4irDex0rXlhmHi4spPxAhav6dmbhYxP3jdmktGxDajpg274OB4ei
jGL1N32d7RVjfDXO5Ur4wzUs/3v8/NDdlrSbNjbP+9KEa7SovvNmDMRO915q9lpf
/oQOUo8xUbHlbtOkdiRNtSf56qgZFHgcOhXFd7HybOEvGo3TH8w1Sc28WcqLXW3i
vuQNeIcGtAva17Nj0J/ADezNiHt38HugXPnPTnMvBb1aP/aas5E+Wt+vWAyIzoOC
QA6EOj416qxVYJ7fadcYXaQblWTW5PA6hiIz4KImJLr1KHI7m0wEsli1N9TjB3f4
/oxOxV8dxVz466NBpOhfZX2FI23u5c3OrCslYzeld7e3OREZhHHPE9jNFT7GMYZk
RVXNU/KGmZNwon+zU+v9colWidPSPq7mVvuaPQC710VY1w2q9VHHKJt1X/w7kwar
24VsThL1FR2Tj2yvX4hol9n4pj2LKEQ8AzCy96pS/JrkEvScu8tlrfW+dKYo+vks
OQ3Z+TclT+2qdAFq9CEURg==
`protect END_PROTECTED
