`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jK4PWNvAznYq81th/0n+5AeJT9VMX6YyUALZ/ZuCPLs65OgUVpj+msXjotOkp4HX
VeAgJ2QZpPamfa8fjR99Bl7KcDxBncf9jmxdrTk1G1THP6XjoEXAP/9N5opo5HhD
54l9rl0N93vjPVNApwAgGvOh5WW8pwUWiF+RDtnZlv7sYGHvoVDyoDrydyhLILJr
esGERSFSWwtBS+ONhaCHSPxk4jfQ7NgcPVH6Ru8/Hj61jXtwm1pree6BopZ0SO9V
OayqdmRmMCq3k4TYotaaAFahsB0/H/jW1EJb1b1+OC90GPWfuc5BiRAjy67QlU5N
5+3y929aMD3mxhcV/d/4VimRD9YrNJxkeQ8Gg81E657R80peKU8V/+7+t/vpKv1U
QQ1QxZoXEujUj9ywuEwWUxflmZuqB4q4k4xjy50MND8lZlctPnjKAXVr/t/6pqiE
+RAnTuMlEzHwlQw8ewDGPWQRfqOL4rGXBjffnmIJWrsQRve4KBt6zw1qVJCWMk10
5J+P5osuMndfLSuB3g4miyISCHWwBrzWZ4Sj7kBSM4lGs7Gh4w/sSaE4gscd2NO/
c6Ev87ZQJtQAKkeBQtTcYLv0xksSAjrGeClL4n1gZdF0Mo+4LnT4q4EbRUDm+9Sv
dwvZFsE0yfP1rpTM3nJDo9s6ZDGQL4oq70Lj2hjLKaQNvl5smZukEcfQPKYYgSxc
H44Txvivmb5s75Z3TNeMsL1OayCbbHW6pc7441LPIwFbpxZaKOVVYwbJf1QUlMEk
JvTZ47D06yl0WArN101IDEJqvvIHPebmtYE40FM0KxTTYqWTQoCEFh686R5G2ZP5
7jZSrjVKJDTW+x1eN6YjS9KKnJCDTP5u0ytXZYR29Knznm4U2CDk5RI9ZVdxGQkW
3MkuzrqgCe9Bd5capyTz5nJVGDAF93437GTJXbVywtKf/jiAA13hkAW5eROX8BW7
9dAWmG6/q+d1LapTdjpZF/c6DC+iBMqCHcB5fUic7PYZoGdQhGeB4VtKsuAKNxb2
51BrkA4zX8JXcb3l9XcrDRY6NDBmtqh1roay5ZHRYkPLCIwyuDPxugZv3SihODvn
jl+xaAjOOJDO08Fk6guRgTRt7beVVSoHHKlVEbktIApHvB0OZFxvbwieNc1bXyOM
w7awhe/wKZvBCi+RBjcOe2Z023ku8XmIxwXbypOWNR+FFUfpML3pos/4bEygTtzz
VCw2hy83JKkQRrqHN+XkcCzbW0Ct0o65jvTZAUHGbedPLivnZ5hTXHUaawbdydbb
9f/MKfw/hoD3PBeBptMmwX6QPafrdxw0+9Bc9ORHAyJ45h/Bv9dvzvCOuNmvvb6f
48pPcHaecC2uF2wb/opJIVpzpxbOLeYda07baj5qMAz0Jq8Bxn/mFCJKXtXflhqG
4z7WkbKb2qgRZ4jOwI9qbaOYmcdFKbRcms65DdSwC1HcJD9T0CXLoCJHNUOBv5fH
HjMCCyEPYFMOvGTENsQNI5CFRnNp5/y4xmprLh5byQOjvKQJgZjLU2s50rf67b0S
tSPC/C2tamdsOW5iBeIHwk0hFzuy2zCMfQkHyBVwJ7W3Aa2Mu2f/w2RixrKZxmlE
TkVvCh8WNr56r4ezxHVyTGHB8w++xWtP61EuK/mIOucBTtl/++vqNB1ZjBC165EI
AlrQ7JMj9qe1nHnvT8DZ6jzGXjcDyHkCTT05ZZ3Bn489zZXTB5xCYZ9bnO2DzqMy
T26KrZwNmt2UqMdTi/5MNUl+IyURfj823NImv/NiYz8gpuY/BxiMgT9pJ/yghZSO
ElM9tytwJe9fsYHR0GuNq/h4RrDcWaLuotJylxmIm4K66qEiMi3lXpQh6BfiISTw
NLUkDZpXeTscSJgXsWp784znTWHaC7eBsN5Yt7gzfKLnishRgTWDUK5mYmRLn9l/
++lLQ/RH2rrY0674DpE93FPYbu6K1/KNtuTANvqRpYZnnsEJSwyjEKzpI4C9Pt4V
pnLeVwRDyXDcsLTUAj6MYsTZ1xuEYBGXNrtLwySEtJ+uZPvJDa/tRu5w4f9u+PUo
842dOMRADzNmy4ixucdCCZCPwca2Jwbuso8TK6LtHVDQWFZM8sTBcPs/iU3Vr4Eg
8qcuqSOM1Dy/E0fhl4q3k8zVAxpNPtj6gc9eKQZn252INqW/dbOf3Y8j/8jkNZtb
Y86ou3XuBsTUYtUmbfNJNX8aQRNBVCTTkirYK/9Tr1Dfy3ML0vKzosUtIXEvOnS/
FtXPIolQcbhBR4OxKokh/O8NBbrQf0Ml++m3YUZAMvY9H9Gd7QqXw4lYawuC77FE
mqkttygQyIJMs4Hwg9eZ4l1fic96Whs8BVO+us87uj1NYnZGptHNir/F6YCs+caw
nHqbQDVsTIs1JUjssnlTe3upHFLHRFxn4XWBYcbwaZkUqDZH4puLBzYtsdrUS7R/
r5f2UNPaigmXuGq31t4AMGeEaRIrHoVFljyaBnpK9H5IqMLVvLwo3UnTtRu7qyW2
X5VpkMDvTOn3+beZI2T7VevR6eWZrbq+xIAj209djzgR+1SmetIYFExoTORLkMJm
AmtlxJX1G67dgaCZGpFxCPMN5sX6MCOIbg/iiOIOaLmdFnfJeMDYXZQDWE/JvzJI
ea9WcpPPwjQvcPCEQ/YXWEOJ90sf0gV1xwXfG5Dn3OuV8yRC/8d/X5o2KtGfh6c9
BYHhm1v05GMy3rLS2z+PAdamSJ5UCP4xU+hphUAf1U4gxMM8k3VymoFDcFZXRVNj
KnV8usRXkOGcdnEvsryhi0pCkcabOnrPm7t/tX8d6UsNGNmBJijF4AULTK7ajlbh
OodXJEduOaLHrWHYiMmi3o5SSKoqvFtEKOW57HUZRudkLOaTkMH1JqVZa2RX9Ge+
D5G5HpVkf2d3qkpkKzWRMaruDkqGDLNXyUq07kv43XTUVz9DOopuqsMrpKoZi7Ul
r4S8IfMWPh2apwxideDQQoEMOmDkfRljusWOfH6zLcz3wE8kS48AGNoyMarWbJ42
5PFXuaBTGfXpW7iIS7O4hfcuD9zLKlWqO1nw38khK4yyQZwfFx63HjzHYxoL/LmI
8FZqXnlFIqWkfn663UW6aERX6ItsWVLFBJyT9jxNWwBRwnrw2mQFOtkd85CqSSBn
1vGZ1sLRrFcmLbpInRUJXWEDvuhOIf0OadS4gMrfN/BUQ3q+uVUPjwZyTlOXPvMI
YQlccEWJQeTLpk+4HMc4iDPgFWCz/5UwI421gS40pyXY/zePHBVTh6WH0PJjtkMX
Mqat6ibJrFT0hVapZCWoe3Gs0wpM5b3umd4s6h1KJ3WuXVr8zusZVhn027L++7Zb
6n1cQGuRXgVAOcCJ1qmEWmf/oCCU7SPkoP09ibCNQAQcWy1VJtydUfXFAf1+nsN0
lIwDHnb8JTwDHhdPhbXV50a0o6FwMyWFhBgfcsqqXuKGt9R3m2dg4orEzuyvWcW4
tq791Z6sBRZLvPg0O9YNum4xnKdrbw+ugTRkmBEk1Zi1pxgYh5mup6NNw3Qpu0Jb
H+h4BVvPOvptfQVlMmdJWHrBkrEpJxCriEdpKkL3Z+dWavenX6Fy4cFGEo3C3zwY
EeYEeP3Lt9T4uU2fu1SewnLel0489eie8eXgznWqj3okihlXndKDUSuhZ49wB+Z/
WOWVdRu44YSeP9OjvZ9nz0WmjxuPm+G8+x8bXZoOqnYiIbWq7yQVaO2LMDylLP/q
AnHuFIbMvbMKwJYvNBUGlGRYe91Sfux1U+Wr2whmPg4xFpw1i3WP2lr99rylI4FP
QUuAxrfF+Ifaez5f/p3UMDssaYPRXX8hnQoY3mCyAU+i077+h7z93iDsugT+U5Hj
yP6rortdm05mxH8ecFUAGwc8ane7r+4iT4L90PjiYjeiQ2tmw5/gipSq8E9jRHix
XDQw90GTzGCCJ8zx0xI/TgAs0zJCrHX9F2DvYvfDefnmY7jZ01bYmF2pXhhLrTCr
WgQFAmVtVSUm4rRyGpvrKmFytGfnyOpbU6aoSLXdoL3212CHuTDrmzcg8bFA4r3u
7l1wF5BevMp0j4v0xJmSdR6rJ9aVdLw7NpcCFpDngmB0/HNPJL6A6y6NHww2TKJH
BXf5qnfGvhKHNkvWKER0lRTZ6Blv0b1iGJeS0AMpMD9lCbRbRik3ByeQ94vmsFkv
fkRKE0FoZGvAJ0nABRSY+7rqQ9Kle3HhXi2TtACSb4xq0HZxhhZZoLgeLacqUCu2
sjcU5bBYWpIKMzIqQYMSMy3ydmLOzltKc0o+xcV6D5wjY7/7Zoa0GmV6DZRMZIGz
z7Iv/yeShjpkS42ZkoeUod8cpzBTsREmnwkQYoj494Mixv3j6SetYXsay4KWXPqP
DSBNYBXQ1pv+uX+qT6O+u3X994WXsgS6CoBvbTiGX05QUJnW5iVCQxwnjpkhxddG
2M5Zrs48mGWAQ6zfQMY1FXgLw3iBYbGEcdb2bU+ijdewnAyDW5qW0p81PuqGRYwe
ro/q6TeFD/SmoZbnpF3lKJJgvsIuKYsnXg8RtMCJnAk3uP7F6FuUxBV+3FznAWOU
0grDtQFZVgL/dUP7l+xHvDKoKKLYoH0e0cLqSi7uv2X3WYbdCwuKHGofpDgV263j
j/FbDPwWYTFHb8GVdJLFSqnSI2cdCPX+fFWYWkWKKaSrcSF6vHRSZORyc1wt/B1x
gH2awlECrAJ78tHFsnlFUbkcsz1GOMWIq9mfTklz2RzRfl7wem1BzsN12GoDX89S
V4leY8nsBUefbq5IUwg1E31GS302+87kcHTWe57mluaNsZeaqWhRyCKP+kVoOC4l
7RmY+BVsXRuPF2ubkk22wvmBGpKfsBJ9W/Z4GHBTQBPsceKk3u9RatgZGAHi1V3z
RL9nDsrMKEQfGDLz4jnE4KHLZLCB6grjiHPqfcabquZGTQrF46tweYEePG5k6/+r
iJUMu46pT454FIIrgzD7kPzi0lvYAdhMne03MKsBrWiUTzQjBKrsbDnJ82TvpIcF
OufbKzdUtqhiopfqsyUiHgN4yWB9HSh4xSW4LmVV1TvezAz6nr6HSUvq/Ui/Bgyo
PdWFeRlw1Vr2ZCxnXllqKgQBVfXftUvfwMuduX9hWcdFiIW1H/toEu7CQszq8Uut
BhY8IP/g/WyE13b8fMfbSWc05yel7vaY6AM1r+1bbrntDRQ6RU32PMo5g6YmRJt4
YRRCw2yzjXihIE+Ckh9fq6cVHSI2S+4mO2cjmxDjZeNiXD8sORv8aYEr+ZLk/m1F
RiZykWYJPRDugzd0liAo57A1mMdQzFr+59z76Vp8Yo3DkE++xqVCV5RX4svZUbjC
3YoFrB4S9kZjlm+8dbWitWafOY7iSypRBS0+mtqs4x3SUZkth+joPkJWsYWHyqaR
VVCKiX/A54dt25xe92PDZ0vG0FYjTepKamEl2STfoQlXJep+/ywtHiJkaOWKO9tw
hAjez1X2CX3V70qnWy2tolMsQ7UfHhBWt2hieHm0av7Z9s0ceL0J4DoVUwfuAybA
oOQXLqmxT9p5rStXPfTXA3TbJAOLoFc9SAFwA2xWWWmLBaEDfCsCChjVi9XrwAYA
uWEZx4/o8O21wYmBNkSzI9FCE0dc1ou1T9tEzJkdvi6MS1f6nLSxEfXRzNKjU70L
kKTdTZ4bzMRcigg9bE5djpytMjU8/sKHwtaH2rkbVBLfWthkgHCUcIQrzYFuXHoT
99TvPQGQ96ctz/cSPMm4b9VrDZUuilq0+F6J7AJwrvKHJVlLvQ/UwSi8puzpY04Z
MXrSITyQ0BepQ0o0BkrHBJqK/+E0TqIWJ7mkxTKXbnSvyM5hihnE7xkrv+/ytSPe
YMfvBNe9jqkKhRCJ9iIdd2m3PgO83gU/Uo3e4YBRmrnblASheFP3tl16K2aAHPSD
ouQuBV5s4wLFBpHB4hCK6ICWyPkcYtyAMvRtZlSXpkC9R2FB0DlNR6ERXjgd/2lG
tgLa1aEviEK7cU7Z3eRWeD/qhXmbEnFBRYOCRnASBgw153UHxvR70bazDl+G5c54
lYym6cDXI3kIl/91AoZ5MLGBiQAzv1pzjUZNUgcvzQ0ftw73sjC17OGWgxTmDjbc
oU1F8susyP0UXgf+MD+csiWOs/v4rTu+eVxyKzXHXzX+2PAdMK7tkC/V27BMG6sl
Dhbdg7ilA6EIUIzOeYJxSnnGfQvsGyG/+mjxhb0HvWkeGSBcQATwvOQzWTEJVaL6
5V326KupNG/Wc6BC5WeL+VS2WPBS4JuvN/5Vh2xF+6RR6G0LKKwoWETwOiMkHBFA
/Uyb4xBuakNR6rcDsFX1WMGsCwgFcJBwZ2zJnUwVLv8LK/moi00lNeF2NebsjCNt
BlhCwTkDS7aUEgF3jpkVcuQrrrHHVBk3cxiBau7B1akynSXmCV1z/eV9kiDfOFfn
t8ab04mFbL/064Zb6xjN0E4pQOqt2Auic/QWp8IuCfK6pNxgrMdBwQtDQ3HhhCi8
tYP3oL0zDjCXStfsbWijRXOZ6ouM7ppqwL6Ykvdjmi0fb5VG8LLS+hWJ9OX603Oz
nqtpdgxlHUUaoKFc60f5cRNZ20QJH9cUkrbJSbJd0vTFDh7ETymbwQ2mqd4q5hA4
bj8tpshRM6Arj0gGbAQIurfxU6+VK8/LzvOvGEpdInZUwbcKRCA4k4jspA3wCUB2
TZC2gNTeAFx9ZgalAXvUWasTU4OeBWob82IH4it8TydqZD9TrVYOUCmUv7xnbR5E
cxdeXFHKIxy7UW4yR7wz3CaLMZMoArx7XgAt35dEyAM/FcQnQcE7ofGvJLfLCx+F
lm66drxfvbGi1FQ38kQ7Pqpejhzw85Cn1Y+thvcNPRRrwsJQaARKCHzKR3DrDF6d
bQx9giMCoS8nintTQAZBBTsaKIdtwSkTN/rSbW5z2UWZFV7YS6AaDoAFkb9EIaMk
6quugOozgickENWZR0Z5r1vfLH7aGYp3doMDlsR/+2zxyYppoH4lmb9tsdey0e3b
QLk5zSMtd1ZEFVLkVv+WwISGIaCeEhU4MZHl/qUGQui52NtcxXaS0lpSc9wJRY5+
mx5afSDLZZ76jGArdVrxIiSF8nhZUebj3Q56pkUwCi/3GnJLYtS4U6Li7R136o4z
kspgLsV0CRCELCNsJvvmH8Ma3mpHNiCj7piHjhszWHg0NmQMf9JYOjp071iAFhE8
gc86t6/xHQ0cwCg9B0P2uyTns53SyPXtK4yWu9H7Yv0pouhuaq8TpFJgaIjByQiI
kjailkeMBvzW9EPL3UvdzChDmiht1pEmYDB+GnwTxubMvppM/b0TFsKJMbqABl0N
GtFAvJw3tfPxjk20xlU1d+T6nXGAh9OHpy1TkEqxXiuV2o72OhvRd+pzZZvAMHV0
b8Ym3jgvPObi/5h8HCAdbhvse4Cv508dS3CxRJCI+t202ZT4KNEGuJ9CT0jJ9Nhn
x7OQ8J6QVijtpKlPhlc+APEoJgv1wWEraGtIKdRcctjY++/Hjt09TTMRrkK5oBPH
eTSuRW5fsqVZMegkUjwhuYLIdlh7bUmU6glkiotWst4QmTH/v//AhE1cRgcLzqKF
0Yz5IKu0wDbeVxx2DEiKERW9W6f5We5p+KkPoP6QVK48thQT5Ag5txwnaH8bQmwW
/5ma/j/p0rJA1u+QKirGmb2uwc+id3ZRS04/IeKGDALXtR2+Hlc+jPI/keRCUOG7
C9Cr0NIfJZ3MktJOXh/+3ONie+91EaZMduvls9w06z7iJpnwlL4loCshjLFUzszj
d26nLjtg27FeQbl2GRi1VeQcx0wf6H1Ryk0hBjEYmX5p9qJgCaSCX2AE5iPznngO
gnr6uEV9aVwyWDUhoiBC+oeRPUyCMoBkt5yf6SADg9X+RiwnkqsTOrOwdLwTbBgV
s9IWRRdVw/D+0/bHnkjPWqJnUzKEYtOr0xqIbmcI8JWKydBSQuACP5T6MVo5lB2Q
nshU1367df/zE6E45oS9hFXEjr4aEKAB0C8aLdN/Rfsq7biBSiGnb19rAf01AIXw
ieUnj+TmS1YY6qSCK57zqPqacKER56GYl6MJbMF+EF/fvbtDzjIPR313poAvx1sE
WlZGhEu/84K7zqanmhrrnJWLKbI23LDvWZXeUWyhYUVr+egl09g4653PzoU7xXYd
+7vQfXzMUeBBoBoSbiI6SLZwvkgdlns7uMJTCX43sEM+euXAdwN8so2shddVQ+kq
fT4ip/YK7uUEy2IwpgUval6rEVp1dTlpZDABrT/FWbPnmKf0+ce+OhbAgMIkp95E
1xmWOOAoMazkNIqihjNTDlaH5X9waLaMiySqpwb1BP7yxOHBe0iRaaFgJIpYp3yn
CvOjmlgb+ZA9/8XRhEzP/23uQxZa2kaKxauNd5XxUkVFafXE5qnYf09SWRt3AGX1
Gp7oXp1xnwPOHIEZ4+D5rm3gayHwCWhlXtTRml9mlv6CpdbgPvG9K3pW+M8XQ5co
Yg1yEMrY7A5ZF6gcjX6RfapilN9TenI1/U8N1PnyDmExKSiwB0ZNIp6eIMyUtgLU
s4iS/aAEMpEbUuDiumv4gk4ImTPhLEhrq1izNK3WIjHGnTIHetgIVofAg1s648gF
g1CiCRZ+m7oP4c5DanBsuyGsTMaS3X0OiAZZmI59IMQSusF1cK9rx0oJ52otZXFn
Qij8ZzHF1ASJ1rLQ/cdTnXtqddCiP+0F0MQPZxhUo/Ihfhy4mN6Zyr2XjHiI7Uwb
x0dcbXmp4l+vixXJIlaNgRpDi3CspprYNLsqqwx+bbqTexzNfa0dyQWL8yWC89Ow
uTKUZJNgGCn3a3L85gZx0Nun2uS02G9lip/FJSr7VxWIHiy69vpd32IsJxn6hmNC
tCWtEWCxpTVQO+CMoVtq+m8k9YdDGUI/MGwuaZyDRJ5AHZjFyb0dYDwfmAgYGKv9
lY1KmOmMbiql1SNiMsqiuVVSj2zkEW6x77wxTBB9CNw9TjYmbI+nAI4wY1XsF9Oi
5lqsy6um0s11LFknTunoRJdy/aO2kXEgAZt7FC6acyDeOiiDRWXEnnhVSxug6jgZ
Lc293joMd3xzJRVJvGMNXjBIZiYP3gwb/X92ksLhChHdFV/P5cY4U7CwSiTusXCj
pE5SNzabMmWbBknKOsWfevwIlY5Xs+pguO77KyHdVnZS779vL7EvHwaRs50Yv6sh
IOxV75GLtq3bZH2fyZmlrHuG3636iKnnqrOtaYkuf5vbeii/B7IwxTJ40wpAwwAf
cvlLTetkNpf3QiZlYEbSgYMny4/hT7d1+qmIqsaf+d9ccZwd+DQSIYnSYOZShl1e
1poln+m8DBCoX5XAxqMpWczDjpOo2dhXmHlZp5xoEexCgwGeremwkdniDQHjsbOx
7oQfOmdyGaXMnsUPUoojOEmxqzeJ5IxaFFIowu6pYWmj3o7nwrtyLNsZuWcE90TM
qigkkHVIeHDPM2W3hl1Lpts197kEop9y5AdkFg1Mm6DGOYySawCR7hw6bXCvQ7bz
pKh+oQ0Edtbo9C/sCNcnMEx2cQ5cropkTFBIZjbEYvSqKEkryesQSQekd2Sfnlu9
iylof5x1r4ePfyEQ5hWre+eQJcFBIWp6Bv0DvBCqbiHRFVu2SU5zPKImHiHBQ9sy
NqkXfHy+mgxlzeVI+n6VqD/mv8OUgapp60Y8awBetXyej07QZ6wZ5/BuMdI00y+s
MiLmijDmwl5DxzdYkNDRcnWYxvfa6U3icz/9uObIDgUOlVT3PnQDeHSe9AkbClEH
RccJaB7tNEEdmmDbhheUn3oik+T1ng3mTul3lohe35dowaAUbPuquh7aPkC94hHZ
97b+BAbvRY4P6UThdHiYB17b5Im6kxElElEgfNM6SrU3sdZvWL/nyGZVPNzJAhUN
OtgtOpj4EY3dq2AB2BGSo8g4EADYlIp60PJyMZLKZvt26az1t2pXb1Y/meQX1i4x
AW5rlIEBwMD4JnGiOkzebBWgA8jlEKRvaE/tdNQ7OOKrn0EfNfxcKGReIgz2sYlj
spymzlh5nV7ZaApZQY3k8K/ls+JjNo8Nj/k6Py3+1ezKHO7V/ShAFGi8uibSjEng
MCalIlMZqVn3msl3//lOPZRrnKN2E/JJ5WGhAMkvNEbzNXNE/pSpuYbsQdvpKKh+
lFYWOYr3K+aEQZ2DiNo6ZQ1z5uMxo3Nq9QbQLM8Vfv1L9W6wYOPU1GN4ugG8Du3T
WWsHLLd2YRWlz6/6VAYzxRgaUMaaN1hxWf8yuGHpgWKHVTevwECqzXlskXEtvwzb
uv6vkVbI93d/79lWDVSsbk9ejY72R6H81OzatJyycAWLvzspoNHC8PIphs8VHppG
hO6T78qGOQeoMa4YRPEruB053BEk7GCyNYwc9q08T1wsNL2iUnmC6fMPWRgLTT10
LrS3y0yX5k0mBNoUjWheyfaYW0qok2WJkV1XHC/mNTc58CrJMEAafCCkyap6U+14
2RAWur+9I24M+LC6lIhxuDTyoDkTrlPrnHNHsO5bstbnhhsXfIDW6+XfjyP6KmlA
yYl8BfY8zusrQv6UVxG82tSosBgA8nFB3iDxFFz8xKP6M+PnUTjHqq2k5jKpHdmO
YNbSbLiCLCKSUCyAEEtbDZARCmEhu8bZtm1lNaBpVbSwvOaBTZ/Xn5pcpOmaCWOV
I8RJ5YzpAxHkqI1jfYuR9+oZpv1/OMaMo+HuiCIxyJmr9KYM6BjIjMpuqMatOHja
q/Px9KkE2phJEvqWsY4skBabFTnQLfWZBIE3dLk9YgDY8Hh7mbvyjHtrD9pj7TOD
wtygCnwUgw1kTnIy42x9DMBL92lMfNMWXlfW+GpgxizsrVWSEwNYkLAt1AvoVNkf
DWvWf57f1c/9WazvcYzWxbBcpDmPdBsVr/5syN6Fak44aR7+CKSpq84hIw44aBxE
qcR9qCEwcSu0GVEbdBDyIyR8UF0G/+EZsH7pvKAQNfg5TR8iQL6vc/8UjMfESJzs
T7xf/W0DmKkcdPxC1glwbhkh+9H+ZiNRE4qN/27BlaU4Fo2LRG/gmpjZ6wrKsyOq
S1W29LRyzg6vV5WO8+TGGSQFc+arIWj/lFabgxi9xu2iPqHYfCEZtJkSvLkc8J98
no/A313TPPUfFVTohzLKegmGbo/wdatepHIlzSEeJaKZUE24pcBkP4qS/ENS5Law
fPPXbgQgfNtbNP2cgFODYYygUBh0H+g3Ms+wf/3st0ULK/b8lsMBTLpbny4YuAaT
+amX7wu1RVZ2Y6PnK+VJCSoAtU1q58X1stg0SL4kvjyFU2iU0jc28L1UPfvanfUq
Iz0JThWgZU8Wp2E+grUA/+xMihUiiOodtyZU+8jaWhhv5ANqzQoe7hdOWiSlTOMb
S7UTXKyc3Xy1cXhDIGMJYpSCc4qj5UZ5CPySb/QLrI+nDRqWqIekG1oN3H6d8ovm
AwoaibyxC3X601y6dxeeG5SH18642Qs0htRpQRroJvTkQVq7mz3vTuG3/gxQyCHo
8yI9dxvpiW4e/PzsTL49Z6O61/TSL1dz2gRJonKYm6rtLWLKHK4XY+7iYEJNwPlP
LMT0j2HHGbZt87oXkxyKQ7BdjuaNkA2MPiFvdfhQ9q7ic9ToTFOM8usF5EKC8bAM
lZSng3Z/mv9HJw0v141zcT+zBFcNLfwZzEuajf1XaPzOMUrcnyHYKwzTU0ZFGGI+
xfCLUwffsYZQ9Xe4HD0jO4g0exTm2lCxy5Xvm8qfThyy0HxIii71e7ZLAewuXr58
fzggXi5eR36uBckW9N+PoBmV18yP9OxDcePCW8voaXCuaxMfaYw8kyBJ0pNIflCQ
ajA/nylvSuXXESwWBkoMB2267+OK0ZZ2j7zyqcdZazww8j2a7ZBwpCR1KDJgZcmf
LeiKeAkp2kWT/wYQqnB0TloKYlTtXt0ghfAYhngvNikCs8EfJ5raF2D8MPuvCDr0
EJIx0am3T6FN1YEtRbA9IxDq4eRxRXPDYSgE4nidlz1Cd9beMB0rQ9c34lZxAIpx
hJKkKTAlIwcStGfFNn4Cd/eVc4D1wYTDCdoKJ7K2dGFWejOfxt6420vPYipE7SJx
Ud0nS1iaWyj0948CG6xRTWkOSPowUlBR+DfayAVW/wYuZdDrv4yqHKa8rp+43AWD
HsZeCEvcP2kRZD1IvHVHD4z7p8rJaAskaEOwrGWHCwPrkc5+0jcvbgJVMUNNkUYM
WN48kI7jYQ9rSf5fhqQtdFs6tGY/c4vdKgH5g2SXVvzpKYOB+eXUbbOCGHyYe1KE
KSI9fdIqBMfICPc8zS59W/TV38JeDvgm4It2VxErK6T3Fwec5mvEfEsLgPyJX+HI
SY91q2FNJGYB49y2dSz7zKEM6kqdzh3A3MsHuAMw0QnxUqrQtAwXJr+QrDgOg153
9YkJ+i12JNulBEKRk7mWe2a2NQsJmx3nhe9I31qI+XsHePoufO8YookOjlZymz+0
aNy6lV8qQkdZ6KguZbV662IeKoaxXEmRo1G9vDQHTB3ez5f5AjR5B3gMzgxXdBob
xMCgu8cW9A/r0j8YeFs9NxluDr17MhNfxLjCdzrTcIi4FSFZIIwrjlI6LrYYgw/4
5nstfM9ttsWZXIsaUKBay8hT33DjAaWZA6TOBWMzF+JHvoYr9MTMXc1VtgqD8/1w
gGz9MTtwsCyHfPKsq/WstdDIleskOQXkubSDWOG65l5bo+tq3uUCTYj/nckXSEwo
R27yPHq3U4+CTi8fT1yg2jdKVni9jC+s5LKBFb/Ol4J9jX3oIYxEdbE+G8d4j9UK
6WV3uyo0VhgObzccIqo44Er82qmLuOd5hUwjZzC55Tqun43PJZQWtvnu3jsCh6Os
p+I0XxDjICp4WQIEnwQiqmELDXtpFUS/tMFn5M7gZU4a2zH3HOtmv4xTpp542v/J
Q0tolBwD0sHM//7VC0NrwNfqSUgd7GQRPhYcxJv9ZXL1I4zZupwM1Nkbbk651xkR
tVFkFCxSQZsY0NbEhfuId2yG+n8NBS7mj1/qf37lLjCwQNiKrCEkT0u/Twthtn0H
0cCAZ2aB086Da5XlLIXKfa3Zx43a/8DxHmBK83bTNAmAOgXH0TIeOo/KK6xgpV6B
QXhmHM7KddY6ubv4Um5TUl1lJR2+xIuw5uW94HHjBHqO3dAzvX/Mv5dZrQJC8Kh8
ZjzxLZrqFIltqb5tnIMjR9emP7s4nzPheTGPCrxiHVdlTMo6QFrWbJwttitgLKdJ
NuPAenKOfcFSfoXjp+PwaHtkFEtEOnbk2CV6KAs0MJ3/BklBh4AP98PU/dgFNiu+
rOFS5rLLI8eX2iW3gJ8uGiDHT9bT3F+7TKNPEWACJrLF5V8aGHs9nkI0QTzACifh
sjTNZg0IFN33jb8UpFnlAb8Q9s09EpYeHhHJktAL7TT1winjbx/xujOYrzj8KAdF
9em59NGug5zJ1OIJR+TGGGtheE1QxwGdP56DjF0y0LD/TG0ZGZcuq1E58jab6dHV
tPxZkmSaqXZraGviLfbZVzX3Ejkjd5XDRBsojixHrlIsoiQRLJ4+C3tVpOvUR61G
SMmdFt24gayFfWU1cJ5AQHEaCiOo+SUCZSPq849oGxLQNC5wSN8jtLEN1RoWZI9u
5FNPgmifFuvcY8BOntKzsohn8uhQzm4472ZTup9xSPhPWE9M/Ht9RjTkz/L2vddZ
naCwMfg+n4qDxUClif/sA+vTVjWiatyWnnFNaBviKXaNb3Npyw5p1AHNElDkLY++
3zlyKEI+9RFxRLNjFMgE4z9sp15N4AySMu/gXV7XoyYX0Ix+rSGmitaN08OF2F3/
E733YYNxTnAlmw4UzUPb93RWhBPdAd4cmZQekv1Bxg7QgdNxFKY3Pii8VgXLfhXm
aW/pyiO9c8jyYMesuwLfxTK6aMnUZkWXIzNxnXfhm+X6gzCbFgDu0UCRri01bnNf
y+YRrIfH3RambFftRKpeLPrHcs8hvTTroLtqx1pfKizboztWuby2Jd1LdmJ+KLmA
ZJNZDpSc9XpO0trCP2JoDs1q9Q9UVSUjokjrlLvRal67ztJSXlEWLvFrrGDm2zz1
tg2+SkpvU6vTpFohqRl/RHdYH4AxI70fMV9r78mlp8L3ftLmgnuz0Xl9hucOdkhJ
ejJP5dATPeIHOZaVxz96g0wBPEPHxYoFlRjKy55chOP2PxRRUGMySGxMec1kBES+
R7jI/Sjmx4q+63L3pN/eeWbhboWmaZ/RuvxR3+2nfRR6km/xG2MEhgY5a9zlTkpN
p4FQntTIsEE9EeZUKzOxsiPlBRsOQPcwmU8kcdAp/ZhTXBZ04PhbUhljh/ZLDy9c
UnPWoGyiNUDSQQZz9wcZh6TU/xyDxXeyUtvE6LgiJavCLIWyU68NR/drEnCbUu1M
vRTN1zSSVI27QjU+PdF0zXDlqmHesznLqzQuRRUL71Irzu9qHzqcV3KRbCzehS1b
kom6PUQ5sqN+Hn6Djsi/IIeOYZ4TUOErz2eJi49C4A3RdXjZ2FkBMe4Fwi9VLMVc
cVo+01K2gfVUxCT6lgY1on2vVDQ3y5FF14ImcBSEDgsufHLwkixWLFy6l5kfjXlQ
Q/PQgn3Z2PapDOrhEePQGafNtA0a4P4lnK+md6mHTdGRNeD5Xa5DGvOmT183DG7c
dkWURLtTRYLtqp1iX1nT+l7ppj4QbrowE/zYUmQYmIt6XXladhAqmMWRtHP4VKRm
9Jf973EvTJzcRgS9noy6MfEumjAwhLq27eQotGctwjtlp73t4KF7IrldK+j3LbZd
CtS5F1EcJF82CHBTHSxOGyA60kh+oUMuh1j45Jme2O3b8gIvKOBSMb0bywe2xHL3
0ElLP7spQV4unEauoxQpAzBzRU99c7m8XwvYRaJCDYK7yKwpzYPEn9zuOQt8CREI
g9SoTmwLQO0fIzu+QQl1cAWPvFXOvHQolPPrbwCoEnLpC9BSvmsb+ANU1u3y62z7
wEMrYJ1UNxRlM+LOBOW9MUTVmbCkRfDrnO3FPeE44OuMkBDhC9CywL1PoUEIAf5q
XkSvicW3Vkzzerc47Kox2U6UOppbkeNHIUrIPSV6dK8q7hlLotgzAP07jx2cOKf2
+MvRWVS0DIMU/XDCjoXM28GBrSv/HX3oIepRb+MDlYNGxtIeT4uKqIalYcrM8q9F
5YMsHy/99WV56P3U4hugelbRGGkDVDJIUVPOicW932LRkxQK89aot2QkQ9Z757uR
WYy5ueZ8q+PeItXqdhi9xyMZflbrE/BUGWXE7Eo6d14TJq3tOawGIZvDtG1OoNHz
yZHXq5MOSUKglsoi2/um8UU/1It0QRxflGtHBJyPry6bvmQa8vSWjeE9FpgMqUTY
saJ5YVywKdk+eX9/VajNNbNwB0WYnDZhNgi3RB/xGFjA9T1mHx7tkeZNHUqt9K6d
CJOyAMhdr0WqGuWAEiKf5s+UEGbmOG75HYhjn1r0eqxEg476sr1IRRLMgJSwjvrN
zfp9qMg+axpMRqDIlRnFP+xkRFwkM2FP/nlBFPkI0x8zmOJB9DgOOu4WqixJppTb
m38eg8YaV17tcM36M/IYhVPBJp5Pjgf4fVN6Z/JVhEva9CbZbcV/io2vIDIfpESt
RvhhA5CKJ5SPbddHbDyiYLB4e94N7cUX102/QRxeKILBzFlt6GPS0uXAt1kVsgI3
JpBVThz3Fg8dtQjh3RMTTrModsjAZF4XNOjWrjph9rS4zos+1wQlo3y01BWvmjul
yNdIp22czUNGWpHDnGQsXtW2r+xi3XpvCHPGKS7skboK5WzeXyI+/If1N4uoTmsO
KuoW4HBIuJHlVPBgBsr0xHse/dkc+TEkHyPP7MmrBfdHLTOm2NYgemcOQHQNVTuG
uHPOO0+wyyV9UJqsu6x4WpTggEVf+Gj5aXdUbK0Tzvcyp3i6C1Xc0AzgjNVW9i55
N1ZVPwb/ppgMtCddUx3LY9wPNO4/C3izkmD+g5wD8/z7cDKRhYCD/zlkzd+VwliG
jqdOpqVeGGvtmSKzu0cJiqGPygHwciTLkA3zQKrVGjGUVZLw+uWqAv1hkagqVVY/
SN5f0xF0jbvbbGRfxhEOwJz5f/p5V1DkidTn1Sym/AlXQJPNznE0xd/BoxjiUiGU
y68objrMeWpAl3Qmq5RApUTiouiRelngSBs+En2AD/eW53cJ0DZmyh0Ze5ZtaBBe
g4KSdx2PXjNoGHdFITuhei+YI1oeDzIRB1wETYsxdgvfgH0AvOXMXN9Ea66RKfrm
BS42UbF8VKme986btpr7YcNK+10+pnqeIgQjI5iCW6Cdaon57cU7p63kCoqv2H4u
f9fD+OsqCmLWdfVE4lLImXZFmry2UwZqeulqmhskDKpSAQAjSpEEzzDYpmZu8Os/
czRky4gdNdhlgVBn5f8EytD/ZaDrMd8lpXtV6HgEuLoUSlEfCqYYidl3geE2Tref
Abm0o5vHg3sZsgr8PtukIDGNW3rhpbSDQgawVZW0rHOot3x5ecG7UKsW18KAAy4s
ko0QItpdpJyVGq/yXAeMd/6IVxhaNqVZsOQiiEgWM0xhxUkdpV3hfu6UOChqYUDe
lADE6P0Lz/w2LnAEm/yw65HWldFGur048gOLUrxKUYJ0TJ+DYkbaxyqICjD+eJn6
LKwz6EmVyOKwvzs7qJiNtILWp+tbL4cvwUrcEFUZl7mzY+L4tUu3MjEQTQ/dqUyD
gVwoM6AccZUKXqexiuUqxMaJd/f01VuzYecKTacjmvzlp4J4uo+j/xMjoYBW907B
MSDQrxkK53ksbwFTHIcNjYMo3/HBsjkYFbRMArioRCq1oVUHIfio66jBmjgnXeLw
QzO/iIahKcN1nS3mMe7lKO+KjvDTlotZqYWpUuGxRf+891R7zMjoYFYnW8j0/Wee
RMd/YthNVvolIqPE+g21hr037jV67lOWCXQspKk5qnHNLW1SNqClk+G3kjDjColL
M+ojTzu0Q5Asga6LP3JnxVBMzhg4Kxh/UDbZy/ElkUMiwzGl4D0py3n6whQHRBpY
hyjpy3t3AoxBeOw0b6nyunOIr43HorLB4t0DTHmA4Bw5Tk4TYGCuwCR4XHn/a8Kf
NX8vXuHIIkWItFj4n2vXmEpD0GcMqMEK6v0YiVfUO5elcIvyBSTem6GZEAdjQptc
/egTDw26xEkylLn4W40/U6rcv6jaNbSiQgQS9tixQ/sxXTCmr5yPYfe93VcJhElV
yeeZQbz1Z/cO2RPD2/aSesXBI8LNnbG8JS5agy6d9KxyRW/47sdI/0cA+Rwk1bNF
YziTaOwlDoyjnuTWfFAtuJCbUe9T30m0609YKape4TlG+MMb9jaGmRCCVfJzQxuG
4NpxUB2kpP0cgL+7D8yFarKRAzZibPGHyUi65U3xU5KfBkWnl7LGsvMKupkOzY1K
pNixi33WczsbPbAPke3yht+TPM1YrsMgMJ4StIA8wp9Gtq0ub1VfhnP2BTYvt4Mb
H18fDNlu75Bx9ey7gN1JowD+5lTTSmP3+PP1s29QkDmoqxeimhyN+QnOScfqo5qI
V8WiR1AUAf1+D77Pm6u0Yh3faApl8UOPcJ9b6Y3brAZ6QWPCWpW9B/Zd6V9HO9Rx
oYhTi6Cc2mDQ2sd+hmxkU9KJKJ9zgHhTJXBPEOMclaGvvPzmUt3eDxs/yTKXylnB
9zq9vD1nvCYGo6PyKGu7Bbk3yB03pWp3uidTsYTEXeU0bdwSnot8+8N7Iqbdvhbc
kl+adCe67oZ16b4/G429rmVfSUNeNfwBSUM50qKxyT3BUEQGJuJeMNrcbYwqZkp1
wOemx/kiuyBz37Ba2+dSUzsImmON4E1hzOXrEtl8TOocztfqyD2dumdZcpvBG5Go
2QNXU4qXuJ2yE6L+d40sNR31S04YJPNG0HDl/p16lAx1f6YWrqBw1dsEweJLbDSo
cJ0Udayq3iomrm38A8QET0o9nY0CJP75+e5Tzusy98AR1KgiuhWzU+uKAYveNoGq
bw+9WbjgMVPIYITzPyjFo5kKwkgV9HQef6L5DoOa6aaPyOfNjI+dVc21Nnczbzht
BPgvW6pOC8paDfirT7RiruZghl7662xYIb0UcC8sXG4Mf+afMTkgqjyzUciwUPC1
v5P+n/9CDDqY/A0f6jdqoWjfUIN+CjsqtSQrRwyE6C8bUgSC/856etuGmXnQxtIN
/wLURnOCl27vffkLLPRdNuqscww1O6ba+MJQDEd5gZ93Dxq6R9vgndPOhe60zS5q
0vRsJo8Y2JnLt30rF7yWObdI0NGYYMjbj9sKLrO969H+6FC+D2cnTBb0uT5dYShY
sf5tyxh4T6ibKFjV4x/v/PXRLBQ1bHdBmTyRMtZA7lVZl/mWBT4z+RmFuN0WHgHp
fS9CxWR2SgSWIt1I/8ts029zBraaaK4gfb8t3Z5MH+11V/TZQHTVLMH8wUJTdDbN
TsqWAzsE2ulz0nal7ZFKXUCjJCry0RR0vx4w/8a6GO8maaoVARMqNkrrDfQ85ZGc
OuroeV901nme7qQxPYVY68nSqIE7Z+DrtPVF/vlRHlrmBTNO+ggmDAW6YcKPEqAF
xyk2HiLboW1K1t9nMJnZrPGz07/e943ZzyhoTQ/a7ocgqdDqr/25hwSiJ0cinT+y
YlK9phVywXx2eLjplVMN3TPIjGwGCbVUkIBcFQ3G+cPtEZ/vmrWZ1C7sbkiYBeh7
DGxPqufA6U4Zidd9G8U4TpeZdahkx1tcZOLm6Ab5Z4LYkWQ81A+l/l3M9ovNnJOk
X/BcUVoOndIZkYCk9MuvRbYwYzbPShLUdvX6TQn+VLFIIbEMyMX9Xoi3OID2RyST
zwfg2mwC5FU8gAHfm217RAnK8YVsCc6YPVrqsxtzYDq5DiFgUFdsTvRsTDx2bPvt
/6mm568O2IbGpSDHg/VzYC4uxyBPElOPrSOmvDVYiY8WYj2qsh2QlYUmmrYJ6KUU
WBEC5/Z0pChOtIutcqjnrg6tFfOwoZu+ieOwcS1Yovr6abqqacqBhhKEkALb9NwJ
dta19aFls/Zqf4b0X/DHXgDLfTo5iAtG46G0Q47KlcITJis9+ah6jLOKIZEU5HHQ
+4w5ET0nEQqzDJgB1m15aiDguihemjzGwvfZASLwbOwiIvWCAa8zbdMMogofq4vZ
Np+odwUVekV4oTl9EzvSLCrDPzZyu6TE3PhbJHYd4DmMdkwQu/3mk62e7JyN168J
Le7qTnOIBhbmN+Dbp7PoOBEmgbptaaBH6wnH0HLikmjrLuHmGMZu17TDJWBWN3C+
cxR2hspF89H0ocLqIn3aarBGp2X4f6LwrZFTJZ0SInOsKDZGeK86nBEU4/SRfger
ChmQ1wQojP3Yt7bzWGFO5JfaGpqv1z5nUZMjUdoCS5tGBSnByWyOuzzujlKplugo
J4yweRSm6weBConKUymohFvMXoQCZQzgJ1h2qahUW1PNfSNtSDG7WT6OANs2T8DA
jeO0zXtrUuMgm3XbDBknLCYYurNqir/mafqDXywDSrtl/62QmDC6nqWiDJxRP0mK
CnZX7dZ9QNJ/ELzxqeS2gnQM2pw4PNYfg2GBx0XHfga9oxQ+s5IbxnHZ1N3ihYRb
F+9MtYCrGrTaTP0hvVJ79QQrpkr9tX8ErNWW8CJAY60GaHm75j2GwNK0It9g8v7f
YPj+fgGmwe2YJ6feT1Wqfk7KFQcoinNALKcrlFA5vcGrZKLaSAadZuTIPbhRNWEs
54qKZb6cCR3P2SNzKNFK7CDj6IuSx3j/QLgCJ9VDOKFkx+D9FulgPJ8CC863HOwE
Z4STpwKYXQciDOJ1EwNDlLS2Cr2AQHlVT3+y0CEWKRt8UUP6fSGcv2n43jiIbKhl
CyoXplrKaghgorRDfsc2fqgd1DH/c98BEg/rfzIUY7f8GNfTgWvbbvBh/tGwmO6y
vraFK5IMpQnMp0JFH4MGuD7+e8lf7Lk5kjL1ppo8A58OdFkMYl7nQahJToICgME9
NfR47+mqPYXA/1UZDSd7v2t9G1I2AEKLpuno7NsIwlpqx0Mmxln5RqUoC0qZK/hV
moSq+XUslnpRVFkBq+p/aAFGyCfwoWLBfV75oAddMabW6ogRZi91DiogSEksrX8l
J/eI4A3XRMDZwACyqQ7pKGtuLbPiranCXDPQkVDKsCp9bIyuu0PP6dobPJRKQOrk
/gqTli67Fk+a1VAOMGV+/YaHkr/xnek5g+eh4WM6stNaW1buY3Jlksh5XZUHFAMC
Ht3ul4BZZ9GUnB0Iomzri9v1FEEneDf9TcMjX21MGf9m6FTWY3Fn59zn03+n1pU+
e2lk5ASDHjpBjxWyf0QKj8LHQisuAgKL6UeBvMBtt6j2YklaitfnzD7VX3GoVTkJ
k0GOxvky/eyQEvxoC8CBAt+UFBV+sz8I5dM17oq+a17z23REbx0FUvr1Rfo6Z93P
HWM9CE4WjlNTwYQAiWNQWBCYfxBVyPLtERkrVklLBvmv7/EvnZ577M0WWSp3OgAj
PFDHpzFSsDPbs3YH3sEr9qAXJfkCa+2Pc0IJKgdHbXd/efI6Xf4qU52FNJ45M06V
sCHKxj7R8yti5lQiTPlQx4pjuO3hLphDrkSywa1Ua6PYRn+cURxs6qu6nNj75bJZ
iL9627bv9tP76mfPjopRLUTJ0Ar31mNMS26CIbuEz5VVW8y/npZ0iIwIb7G8yoxg
SX78o89dO7C5Fr0llDycqVWNVNiBVZUMDU7uPWsKYR5kwoFGurGUa4cOuY6+zggg
5A/XP8HEjdspavntuU+FQxCzMv5hes2bceNH7vU7ppqNvgdqX1LbLxkgDsWp92q0
s23VEsI9deN9Ab7/g14YSRefE2hpCEUAqphWzIjP/2S0ZENc7+iNzh0wLpfkvgPv
3Xl6p8CtgCL9G//Az697QaGzFJKxUntI0o/3N4+zJ8dxJFZeOmYqeKgXBaa3kPil
iz8pXpl2EaysFGh0g5TKk8ODjikoxzL31ADueWskhfCpMIUK39YVP0xw+qp5lvBW
wdHDxsw9bzSZqwRr4X5AfGE4EtOd9+I/XALq69sJzdMONAcxTzJBJAofkbOaZbll
m9qgbnSJS7CYMd1pH16mMl5JrE1EzBeptyayVwKOCTEwe/hZcUQHrsTzfuRqa7IB
jwi5oAJL38cdfGsi/qyrBuiWa4jVKDuh3GK5eNjon/45BQ5sXBD+N9eK5WUNPJUz
6y1Hb2B0LBTWWVIkJQ65XSVr35sS3SBI52bvu5AOuWt5PwIjl70EEZJOqcxF/5bk
DnENpT8xwsFP7sINFq4EFMsAaUnSVZQI0235+N4JUmxzfYFbriCnU39XmOe2zlpi
ey8ZR/t21gZ4jiUzDkxP69rs0A4S7ccHHDnYwLE0oK44eUgTPr+R/NiHvt7EgkiN
5iUVRbxlCEZjFfRH7I9a+gUfNrc3/ZNTjLfPLq6M9TK3vpzEpr6sjLj0ds2R652f
pgM/Szb944L+ql+G0h5WJUHbmo5IlJNwYadXNo/xz7tGrTRGVJvexXKT9EUc7/vz
duAfzit9P6tHJl8HNmTTovKh3mPEosI/pL87Kheeve4kLhXtIEYxSl64d08AYZ7X
i6hgWJQXDER76xeI/zQJH3xQMRWol+OYs+nle6PzuiSJHKapOxwgLGOlHejETfrC
O6SenS+t3yYKscjhmiE5dN0C7e2zJ/Premy4ARCWSKwU9tuychpRfRYrlbf3y6Xy
X6+N1jhTSRF7BFuchN2LIJQK0+J/xmEqIeJhssNe174PV0Ff5d8Rw3Ou1bC5twqg
FFdKD8kIdlTTvI+58VW1pixs4CEN6YwzbMWdRPUPOn43byGbWHhhwpdc/R+AdZaV
e5nmd9BpzSWIgG10lxreUtJ4eYdyzF67/SzTQzV8Ucd3egvTurR+PaMpXGFby9F6
/2vSk9Zkd0wtCdtQX7JJQfDvXnm7eCy0jenAB3lVTvmy1APm7ziOtpsCykh/heYc
eU8PbtWXJRto1G8Xp+kgSIxbPKL63Wh4xE+QSEHgjntUaWDWIdv70S0Bxa3wYeSZ
fPMJ1qx7IeXGZOk8S27K+NO7ehzTpsWgPG0jw90Q9NQYtmxB/8dPJUCFZfPJrOaH
0fdRHs8Pn/NT3V0fYdyM2qdbXVVe7lVVCQ+R96uk4/3RgHYB1Jecu2gz7TSgjFj5
Xs+N6i7UpqQ2V9Zz/A0bxiMgDqUHsKT7YtC4hZcdoDrhNHNPltHXQsiurWekwzoq
dj/5ANTvZhG/sEu6OAFjZyX7odeJ4aZpARc3hnjc4IpxWK9n8yRveRo/pdDGq/hE
QNtNoj7Hp6UqhGzyw+6HQjyZyUUNVTLdkWBSXrxq0PJ4w0031FeDMUdcE++1rGfy
pMR3eFdBob7apMs/1dURO1KY92nXde8DGzgSUt/B+sJWf3owvITdAg5MZkBD0QL5
YQpYHPIpWM1agLJEmLrOM40mTL0QEW0kRkvn0NV9b3xuRfi1bdktw9qObcPkJyxj
FxAr1pQiUFwYGiSwxIY+cYGt3fJCHd8bdErrChYbebDnEmw2h5uaij+Z5trvz0YC
i+WJnPgblt7CDqVoPsX5hiK7RdrqHpI5i3bXu6PTQxMs1q8dbbQ//MAruRXXJScD
JXR+igVtfWnj96rxWG5btjb9PG2bv13J55R+9GWLoj2VIwmZesqfwRG5Kq6i+R9W
rCe9Mk/H26Ro4Mn6hohG45aVUIAASF8fIRhb9V6toz9+rK7U+suyClzj68N83+mM
a4Y11917imr+hn4HTf4cbFkXmBzgQfOf8dK95lswo3hI0E1UTdfKHrbnkbSIORuO
wDgWkrCqOBFeoUIZnaita3TltgRwFvbbqNGpDR+1YLHaX6FPJFthUNsUJgPBvMya
QP7UwdGzMQuxZRgu6S0UzdofhBfGmgo2J1hxXIXgmAa5RBURRowuwju7R9195M3H
WBJT9+PJIVKx1wyUPToCCWmfzLepjlyYbSfBfRSC/JFxDe6Zcs4hPJRsYkkIrSCf
Rcc41MlJxp7GXQ3hhAPE8wf0yTZ13eHIITUlOBvt2l7CjCXy5nusV3TROh1pzbD7
l4fjj64YYCB7f+iTwHZd5E+xKo/zYrKVBd+D/5eqV1HswB9G4l3oQHBLYi2R0owO
K6evjMspU75n01CpKOxZXxOf/OXhb5TkyPHeb/6GoTRYhjikmeeZcIgRzoV7pprw
9k/ASc37XhOQPQ9zM5izgJfjTJ8HZxOwOF+rJWDGfsFwl/SCEyIjlJElvufcwesj
Sxa36Te8ncTA1BWsjvWMi0SlI2UP06KbZqJ5nZWHqxsO5JivitVBUGYArNivo4f7
IgkzFPufzxkPvgS1PKpvfEHDFi2xz+0NnjglqP3lazIo0eOjGPqeuiWk242UZup8
2h79EdHx3pmpG38Wy0t+oGjt027hqeLQVQeQ8H2SPy65a3D90r5jYQ6M2dmvW9PH
m/f4OlC5jbu7EI1pheGdrbZ1WppSY2oGNeFHkCDfAGq0B7HkP0ohYs9/LRmDSssf
ckCcAuca8iAGV1M/UhnL9HbYCabVnpGStgcrohZGHedkUmC4nnhKQzQ88owJy/1D
dBIsL2JqedNNf9kIbeH7fYGMwmGKBrYIOvvEiHjsaVq5qTvZZaFXbl1uFOBJKXYE
diczZ9tD+k2cOshH4IEtkPW2Yybij/34rOr3o6nTbBYjJDiq9McM0Wbds2Fis+k4
IMXucdEZHrZPLw+Lv73FMjPaMq9c4JsmX4lQpyY+QgIJfxkxc2SgOTz7H53BOnGq
QUoZKqw/ukk8CmohW6GyRUnUsgfKcZdn+apZCLzgKyABBoJI5IDqEkuQG6VRx+Az
gnFurR6FY4X2D1aTbd8k359xGWYtEJotqibgbMOXvuD4GPcWS4QnJXSs/9xYj7lf
l4ThgLCnXx9Jjdzdd8bWGfa1wssvMfc2JH1Mh63jLlZiUfyxGMFQqhQ7PqwbIJTG
97cyIhhdoph/cGm2Sugk/3vH+vDt58+eE6TQTqlBBfNcIY9eG6z3ExmXpZ9ovL36
xRcmbsEAjH6XX/RlPYiDlENeciVvndLucP3EeM9ebyjiC7gpSTV52Q/JRmbK4QNr
h0AYVdpVtxMNXpVBB5opShTPtZ0vVyEKZMrtnTpLjJj+4apUvCwERgvFscJzpXmL
/OzU8PcILF34A39nBVS0b11MQClq0CJ74d4wUkPPHerptgvIU4VefdGLnaSj5rkv
qOaLqjSu2NSG+AwcTfyqOURT3iV43++xE6HiYUMKZw4TMCiuE1SG93DfTqO/Tknn
fmHdbBzw946vSO3JoeG2g63BW/tXKhUneMmWSJ2rQW27ZuJW6dVdFksXK0Xkf3w0
NtqssmH061ZBb1Q4vITklUI0mscznx5axjXUNVmyeR3DBe20hPT8kU7wiFwRsyS0
ucu9HIUDu682APAQBiOMRK6dVjRrLwQOOVs8aYJJo9mnZqSSJjVSw3r3R/GPRNZV
KLj80g/+3KXro1vrt0/3HsgeRRUFz9XjpjKy96DYhb1TbTxmYCSAcwwIxnnSDDn/
EWUNMhDqs6wqXhEXpcHt5bXBkueDxrf5blkoqrUSWU1ImIBys0xxOf8qpeuKdJfh
WWzoltklvrbnhD2uPsTI9qcwd82mnppj03hbsSJSMs1c9tLmSGCQkUQ/BPl8KfIi
WZ1V81sNLCY+8kgCs+w3eZWMdDr/L+EjlIfvQXuwcLqVynkfpqsWcuICZ7w7SwhB
vVqBbr8x0FqRly2Kp3dGMz7hdjiDhwJnevhqBVCzUBOsUU3EFisAVphKQdjYjyRa
svsGjEsuozW9M3PqZI0cAqCaNlJm5yomEfOZSVGkGE+XUPynSAoghym63Wv9Xjs3
APZWpaWy6i983tvJRZGbg1TLGxykUrSeZB6EpkOJbm7uONxcJjKnVlkGEHwsJxZz
o9fZQxNPKL5u44CfhFHFjBlRZK345e9qhvPX6SO+CkvuLsYhJ/0EJTWMZ/eiv24v
KI384ksW/67s+yTdNE3tVzYOdtOuPTbJm0mGRdWgcE100lH2wSVOLa8HF4F3Znol
wqzUB/270oPnyBle9OrbpDSlzlZDxgxkqTDPvuFUL5Sd8g16peqUxAkfL9orxhEs
I3xFX6LZ9bDPVw09ZLlJQwqTRbbPN26X5D901mv/om/R22BE4D89YyjTdNZRsWHS
JTJs9ZT6UFuFEcjoJRFqRFpHejSXONeQ8WnoGcV5HIJybUr40fdtsjJwyut4fd1L
ldHZ9wCxprwDcXMF2a/jTOJConOm87hW3U5LpXWAG7FqCNhgrQBzqZXmQS6v3vJW
ggMybyprVjzSP/F517s/39KiUtKoi68cjnzzy8fzsvbIHLykkizXdqfYvlJ/CaPX
SCLfl3FFmtHjbrzOF8mOGaSSjuUIx7+DF3KMC/kdTZWEZGvCnMbHj1ukbUBj/Wsh
3GecOGDNptH+gXqsDA8fMYhgowhGLlCVNOc385QjZ2XDlKUEtbWeZWoqTIgdy7Kg
zI7oH8GAjmTMHt5Jo09cOPOpR548g6xW0W8Bxh4TIWU8nBT5ApJlIb17RFv6ALnj
wOWEZ+3Zp3lB3Vu63OYOOZZ3HXzOEVe6GEtWcl0E6EKIiNYCzWNNiGbjxJ5exUSC
IGOG1u5+LjaALIf5T/DAWFMrYcPVEAxr5peDglX0FNzUJtCu+OtFSFNvZ/fbB2fw
W5O9rpE2JPoHbN76O2k3/7faWP8LD9KIYxr9iikpuchsuTWwIobdZLwd0bKQNELS
DOhwBNdz/AsZfhcLElY0f11HiR3wNN0qqxo2oer7Ycp+o9Jv+FUPfWQ/kdgoGCQG
E/5zAws6ZO10FcIR2bWIOK4EUnlvj31vWG4lCWbMWQFBCXPWglZ7UaphxVFT1zqw
+kWx/cAYINSxbfH429XkBKgsWc4BZkmaku849KtTlxUJNkR1H/GYmu35iSIAQcqo
y6BQ1D0j9okvJupgAlcfbkfLfXTl7FL+Q8/7PeEATgIRymgMpfL1H9pOxJLxmuIW
VjyRpRIldDX/QUJVkV99WDRG0RqR5vNCRZUPRQWylJuOZyn844aAGNTgtjoP1kUO
Xxyt2mCmXW/bEhcQwPw64Noz1YCQyUNdhoCIjOYzbkKif79DorncKAmeEl41kCTU
MibfVCo3ZpfZNaxh9wJpAloeCw4YS3YTTaK1fnELEojAgeGVR2rtvADb5MwxZ6zt
7YcLNHjvD0sc7c9iaKwSR4m3be3bSRysxdXaq071qR/OpL02MBWTEP4jBcOIk6UL
RHxkTcGeTzMLXrGdnfI3YsuOwgN2G6YQfdNu39gpPa5NYKHpTycouFDVscxeWSLL
E9T5rPSYRy3ruttXjTMy+Vz6N+1xOk22lyCkcmZmXWJ4I+L7NIEq/LtLf8F+/Aa+
3TAWur9flP/iqJEppYoqhre/VZdEfgAkGVqK06NDSOOo+LnA8mODMU66uSWiZ0/X
7rSXcyGGk/+t16e/HmxMpoxdoLW6GTzJfHdMNTz4jQxRr5jItzWDvh4GrnMDIbju
1uQ3OdLInLm9/Koo/+jFews2vd0KcBDct0X0YoP5Eom02Oqxb0cYR/Xvhai6x8iN
FheC2ZdaP1BCRtRqs4aR+JsE8TDbh7+Tc9NzEZDntnomv1c+kAe+TPqGJSkC59NS
MIiWMEqysAcY7DyjT2Vl3XZtn1r/2UUbrI6woFnrjcGn2VjLtqYt6NueCpgdHtTh
AoD4bcPccMTRQoAR5Fl39NQkl9aSYuEA6H3UDY6KffvfC3Rky20QJIBi9C8h6pF+
USorYnnp2jT0H2vW2If9qi5NPDaKhUnuDPboPvcIu1k/AoxVV3GdBpc3TuZs8g/j
MgCoPvTxFOebOUX0AUUQL50E0FBILY78PsPwCpAha/yjn7evibCuv9qHwFevc1Ej
6oCB/MkXJRsuF6ER/iVPyQNoFI+G+9vRe9JuRwEE5vqknHd9uu6UNB4rF62FYBn6
oQU+LWfYuYrBl/ws9PpPdwQHjoe/6YTZX7FCz2roQp3DsrCESdlSSkcd0S8rMsWm
HeFri6gneqG8oB8g0xy32HYkDGNvZCAegRhmzYHZ3Ut637xI0TS1L9tbM8UHlm+b
Z2WdTl1UJnSMfAUS8Thw/9/ZQWdUmP0PP/iWvovSgkcv2YWyoz/rJGGYXphKchP6
/h4TlP9bAmCgM1YiQTksY84wbACjTs4oatEBdlDgS84dV/0ncwM7k87SAw+Lk0Te
r4wCuh1XXFZ6Hf82QtSObXNjda/cE1uky2myee107UEQjQXiIUmxsIz+6a52g9JY
nrr0BDEXqPHthkqM9R9IgLB3SMgRAOfCusbqD/TsAOLiFiNIuJs1XXknTxboNUF/
5gX6si+Z4wMqKiMn7mKFq+VoSg3WD6YtLkGckWZ3Hy0M9v1bNu+CtSEgCxRMlWLw
OI4MM8pWbps9l1+k3G8eKFxnHSSC80vEMPWeHH1s/SsN1AlFg6Z1PBV3kl9QsXEb
fz+hz8gEqdxa0YDzCt0AYcYNiTDhzZr1Hb0AT6COMzghLQWxoMA//Nn/PIaFVow4
kAM3shU+WT3yBPnPGkz3RFJSyeHYpNDHPzzBsfa2NzP402gkpWbTy552Jlvwb9Db
6zB3bfGE97h49VMU+YUlcV7sUjLDi4PcFWi6jvSkN4Vl/MUZzDlYnoHEOTsyIuYc
wU2G9MiZF4XmTzi2iJh732W8pubxGOIjQPnNbLbrSxt+/m8vSKBnindU4EuSzk6E
NPiJxakaw+YRLHVTFuCXXxTcqR80Wfd5Kyaj1+B9zqK5aEnPi4busdD4LNkZ+6h4
VWPWRfXZ0LLpKzQAe7sYgMFyUe+zfvOjs44Zz1ly6p1EvGwRwGZiULggQLyyytO2
mX/8UH4i5hGwS2Tx9/QTFEylYFD/x2su0WUduA94XZGOE70uk7ZNW2qmDMfHtvOA
4e1zr90tp5itUJ92wHMJA2mM46513OYW2yFDfJjzZrew4uKwo/QBSWPu5ank9LVk
6TwmLlZFw1b5XGcUsk304dBy3Ft1bIE25LJZeVmV3qD4dJw71pHNVH8dZK7ZnVDw
T2+aVZ8877eKTh6O54+YV3GaABObssa5XUhG0PGcm5zYxULPRYLbGebTqCXX5QSf
s1TgH+SDB9QEs/oOb8dvk3j0ESjOLkvHSILc+QT9tRy+fRpsE5Dz5Okv9/gEhQy7
bTAmHDdiU6Nr9z+gp6mZK73/LfYZhmvy/OFa0i7WFQekpLaRS/t2eBbbDFj9B6K6
dl2A4x8Dap5rg2vYtl9RRbb9/n1/JMfeKZMrp62R4hL94fCBVYMjUD3nUW/6Q4eJ
sUeI/grYbo+Vx57WMHv0cW7khAHfzOWmxhgt2kWXE9h8qhC9OqJA/PA4YzG6BLNp
k8KHU1fHK2LksXMfr5FF8JVmJIcry/7ih4gJ/bi3w1zWsRjLiAcP5LNpxdU6HBn+
t7ay9qt5QyhRIeEPAhRJ6Z9ZcGbYCKGAqwUZbkkh17OvpUkdRgIyqhx3uwXyPZ+8
rf8AcKAq2mEFBR+xrpFfEMHvRyU64Uf3ZgcCKHi5wlC5b7Rm8qMqE3mbhvKS9rlj
XN2XXGgw0W46kD5goc1F2uIR6ScZzPMMRf9ArtvH15m0r33FPfWx40Sp1Vl2LV8E
HUtqP5ezMSRpwlumLyJ7KjxVSsAOzFok/QmMsVUcvxmNkDshagOXXU/Ad+hlc6hT
X60oVOXLze5p4ORqKpMK3NWjknhpMUgWR4FwMdAh7WQa7QDYa0lnExfeCNUka19n
W3e0uHk/Lff7Sa6hB62vk2VMT9yiCuXdR/vP5hu8aIr6sWdXaazsfNB092kPZdNm
Vww2nXvpR5PsHlToV5K3g4tRhp/txnjWDgkjwCSEe22QZEt/1M8XxiocJfrP8TUT
Vt/GO2bvA7U23lmgZC2cQFHdBmkRe0AiYldkFohb8PmAzg5NvskcH+PSmT0Ekzij
3wlalElrYjf9XuGqCbX2gdQCUlNtxoUJOrcQVQ9pNnBQHAVg0KGyRoRdXqebzsaH
SoGmoPL/Uu48wAu4ThT/QMwaYMmqAjszDgBHwXZcRj2ppzMSt98Zetl3VnM7rtZa
JEzQkMmqv0v0DEzj5IZhk+LidzxxZUw37BHzWZZdaS+r9G1J8dtJDKg1l+pTtJho
eYylB6uFbwC6/qCm5rq6ixAoC13grkXxpEqSTf8Yw+d2BvoQhJPM0pRwS3dAjycd
y5/rCvCZpbZWIMfiOu3MRoxz8CKYIK8EgY/rUQVonWEha4zYkrNRKyolQ5LZXkBc
T1Cns1XVEYlt4Oy2JfO0xtB8dsDBXhI52HeVH/mGIRvsobPlWXNYDI0XVcc2fJbj
hrYDOUfbIhvEL/OZ6CSdIvc2RbVQdTqVs37fDkqoa/3ebu+wqsK2o4LJqQzrQPcX
udQ7s3WrYynvDsy1rcPut108oTyd+4m4/9E5qvFx/Yx0WBjIhvYVD5m9BRbBvWZz
L0T5+R1w9uWW0gEs2IA267dTi/6tQcrcxwWglpGTfv80B5f5Nkj0ZBGH+Qlir3CF
FJxq6RUkbNUpeX8+j6yHv7dZJx2QbsMHvYVPeh+j1B38NW+eh0FC3DxtIrv9WkFp
xgBwIt0bmtA0Il7+Jc29f1R5RTcWSoDAQ6pPjf3TeszVU+eqf4+O89sgvzNfzw4z
OUYJW8z+dAPBrvUAkU+TRd9hZS+zVSLq5ZtAIzbOjnBbTNspiEe98/5790PtWYIs
lZjw3j7ewVUAIfrDTi+eBDskEVD54NZ4KSNcEaWFCxtrTEgmrbmrNPRODmqqetzQ
6IFGHSpvcRRZ+cHkT5liQxIQ7iN/DSJ5V2i4dKHJ7qYlI3yl/Q4mvYtbnOFDc7mD
PVSBbo7XjQRMqVHIx+icuMt0K0dBl4xnbitSNSHjeyx9UepfekKeRS7XHfk6th/E
i8lXD78uWsTWi84OxFAIhgZkOfQQajkRK0xj70aYpeKHA6G605XWRgUNDi/PMimN
XRlmNzosrrHc+6gnWQPd0S4TodX4T4gKVhO2CbtEFsJzTscoucUaU6vKP+VJrKuY
l7qWgpM1P4SidBoO5cMK1UsRM+98SPDFQdGWLYQvd5i0ExZQBGS2sAYCyy4WTM4E
FtQleM7zh5riVRayMi3skIW1ACb7ZW9Zaw5GDoHSKHOedF2L6K7l7eBgS9PYtiuJ
pPnW2AVOyuItO+v3I01NYVOQxu4EftuU2HgwhZvJg0Dz1/cleBADd+xjf5R1vQAg
HYLLPK2Y+iwZ+Oe3Vwe5EmemWH5xEtpEvV+p33vitszUDz/IQquzeigtUOEDRlZp
5nCrCpB11EmLdkF/8JG5DBpr4lZSyLOjLD7S6KONu84+1+je9929MmcRiKZbD56P
dEYTzEqsPyacTtEOTj49/hg+X1rCmxFMFaq2iYr8/ApLDpVE/wRMQhEcR751mM8J
qFsKIeyZMYKXAkew9zbB3LCRn55Z27GZJDf4F4/iFf+w2xhOBal/mKUM6lZPwniW
PBfOnoFtmiBQFGyLwh3OQ+w4KBVTVPzBbKSzVIfxhB0f/ZDwQiYKyq34gYL+E8gq
aREuRNdy3cVv4WZQenoOIE/N6kEj281F7+jE8jxxmW9czoHG9T9CWKFrsGVYZil5
ViYEstkvZ8nkQSXNQLf6AYU/IAE+QHnOy5q8tpC+DNK0n6C11+l9BORLt1uNWuMp
mOlCgGAku/oruO4bHgywGr9JlU4Cjc9FK4eCVs7bSScH51FKDstsbaMr8dJVFwr0
6/R7jGAmr8Le+8qblBWwsorMLcNeu2CSdwT3tEz54odHAlKLLmIoaTcUmL4OmFsb
fIgHs2XErK7DrjH6gLrGB3tJ/oBv1LXdyxYckEzwBSvH9vJJ6zwiaDVxTdHdE59K
DEdWA7dgjagjkso/FdyQuCEFYm3KLURbnl+fK4dX3U/j17iw5gQRQZs8kCvYCCT/
Af2JtRDJJ8K3Q+aAUJYEc52FmGM9uLzBCntxdwXLqzuYVNOzx7J1HYYF0PvBIHre
AF8zm6Mt/vJxt2WSTNvi+keQJYrqECWaJ2K7aLVkP87iCFZtkmeYbmqoGzvgQFsn
fZAt7JcHM+o/xIdsTjSdo3mUNpWfk1Y8CYzBJnJU5aj8fTCT1p3vOGLR//q4yGNO
39WLDcNP+Cy9OqAl1Zz9fYRAfm++n0jNJFrH5lrfgikqGh0I8K/NmejZeIknhgP0
0zTjPvCBckobKGRQpMtomj9liU/JaO9BeWDJuzfNwv6VsJwgBtJ0zZO9tbvnkdxh
Ia0Tr28kA7YROHbsA7Aphsgvc7cr3KYGTHxkiAMhEEbivOhgeOFtUQ6Zh/AVKbYw
6lVgmEjb397CSsyU7hGiIN859fMdjgEuG2tCQAqLbqmfR8DnMIyplWAyIfeujIZ6
F+ru3CARohcS/G8F1ZtT/sQ8l5MW+MFOT6abpSnWEGkT2Kx1AzHWq35KcyMI5dSI
3tJqabfM6hS39hVsXcE13/XhnmlFXdiDwJcjdsEEczRaP7AskuOCoeFQi+JiguRL
lc0wRfM3lbeApSWvvgN23pST/az2ApdWDEI7ooOdgtzVZcb4M10pkNavWsssZ5KS
CLY27w2sB2uPsptTpBzyusioBHXv6Qf/NrIn8Ib+q1t5O0MAW3lKQAXMZlYaS6QW
OQC5C26L6gKIDTgpn9mPRKQcThXE4UdyMzG333h+e2hTowU/43Uu2f17qHkFIhtE
Tmo87GzA0shY5T4XzD4h5TRvn68wMlzgpABVoGlRMqhyo64n5uRB8TqNw9lRvdot
BEYr8oeftK7M307Ca4UYk/xoyy2xdDeQGiJYXlciKFAmboLo2aUIsjc6jYLctI98
0cjCYCGXYpmkUvlnFuB60je9sXzLy3OVAX9xcmQ7RQm1xtrcUG1ilY064cpux1nZ
vfrde1bk2Y4MMXcHWN2fFKbt82qFBgHHe/0khzWbNSKAn+mmkC+A3oKX2I3Ko16y
njDfIj0INL/YCg88VQ2YZpIU3Kt/5prBSIPEIx3tMHWgswO19nCGjfajFE0t9dPp
dlDpRbD9qvFyKafoEt0FLqsWUjmkIYhnNsddKmVZB6Yp76ZAfvGis32I+v7GAzVv
9/CtZC+U1DdCUMpi6DKhm7CqJMuKqRtj8CdaPqSVuYut2Ru3Ewc4XR61l7L9UByF
apltVYlJqtx+rA2wo9uw1UlxBVOG1VSQ7zLtjw+VnEKsfGe+qGiyCmmPUMby851e
IaWspOrymy6kIkonQbYcPba+M0YVFWr0R0X7PD2TnRLTgfD6fEC1QF23LSX0SbT4
kqzLYsMQcEnDMFsSMW/IWmP+3aOrq9WLZkZVT32Ww9Kmc2UBHODmHpVfeD7Ptxd1
P8Q83xkB3CKodrPPyyIZAXYYUGITj2ABfHpRmC21r2K32lLXC74Q4LAc9f2mhWQu
Vk2WBjR6BRct4zrYYimJTvYhi1x92wtq9CyFXmbssX+N/9EWSKLdJJ+EEeVnE8D8
uS/L2ALFCwh9rWd8sSCGnVy0/Z+pRQ1Ue9xFXVRy0pPMThWa3FCd5h2Sj++bpLTq
N+opDzgZnMCfzIMpBEnTV9dfsq+fxCgJqB9qJosYMrgTWuKTSi0+qIYrjrTh/TBY
fN0GfLQ5cGNBH9XWoqi0zJN2PbCDIcjWznBwnvWk4YpZ50SEi9YE3SiKeqbid0cj
9BYrBNd8RMjT6ASecQBK+07vVHXls8pHjyuoaTT9GimsusZ0PbNaS+Vv7Wn1P2oK
hO2m73PD3FskgeKyQ+UbwCs7e0snyRnevv3gTgGLBFahMmPbFklV386AMKVpzNvm
3oDgZGopNTumo8hpWfaChif0GC2A0k0U9vvNzdBCtsFUQQq/7UB3YfuBncKQ2Ge1
cEopEymuwrz50meKUYaHdU7DaNoNBTWP/x0RF+7VSQ3WXsuA5imgwnVZn618m5XU
59xx7LJlx8Zpk8wBQybyiidu/dFJ8jy8Dq0mk3krOIhyKFk4VFhzftlogWJZSrFD
SmujbHnZ0cL1AlVDd4wiPoQZH9PUoBAdYt1SXrUdf50ips7e8h3CRWnu/xdoDDeO
ht3dwzLDxWIq4Lzu7jtnaWbi4YTDwtWv7YC7zF8ZsC7MR2gukULIUZZMRYJNtMJd
1HVclr8zECUD++TEEJlzEO9l7pNt3OuyNl1ggtCRHjZCVGd83+OWSaiF8Sfy7dp9
fGipNAiOH5lMoU4HZyVIu/zB3OaIxsxELSNJwm+R3uEO5ZnytqoTVUUJ+vWsz833
WWr83Rf2teFF9Mg4V+RvX99VWdJze4TOe9CGiijzvV884OhCjULbupL/F0R3xWlo
lYa/1fpsBCzV8To0NxhT0vnQPgEIqVbHzshyx8fxtRhponH4QCdYmDPIQj9S3zdu
jdiXemK5aTKBR8g6MWcD4gZr3lPGFZpWl14jyfBqu+TQ5LNLH/+QILlEA++pcqiz
Ad2DO7oLKObqc/PNtz0FTZg60JEWNR3YOGZUfL48YU61e/CyNiJsxy4bHDoBYz8g
dx3hj1B5IRoiiKK70LRM45GtAl/x6hwpyg4tbdNHMRHh6Ko7e65oP6BNaz+alCmB
2LUaJqW4VZcqE3Yrubo3RbC6Ei+Y1zlDsoxNOYhxjAtVrHArhFXruJ/DG9DpDbgA
djzYl2w6i5r2w3FgfgcfB8c2fsoJJPEiwSNmqVK0Oty3Q2k9moySTkuYoDRo5MUw
iu6DcksagLMu4ALmDDCvaXNJ1zu1yPq5n8HTxObMCL1qkR5pcxTQoHhdCZ9N47d/
zxCsZ/mHekL0bjzovccURywvBcQ42VWMFSvHWXCOKMr4tWsdgGwaZPyZoQ1J1YP+
bT76NqlpCWgLmCxQDes2OALHZ5Q9Y4BsczN1VDtG4+sB7zuQqt+OBwsPYEV6NGQb
9aGhvnVaFnxhMXGNrT27t6Xlu6LFofWLvoEStwQoXtj9pWTZrVUuLqfTdi9j/Jkb
8VFrnluJPAjlYU5O8nefIEPo3v1QPrk/PaBZ5ebnHFoPthYEV5IKLGnBSNcBmxeK
mNGlY+8DwijVnlj/FXGm91Z+0+Vf5cVNMmZoyhyZV0T1pcmnvRVKcXpbTySwTQYw
peb4T0llEsJ/1IgDeSSn+xtNfWra44nlYHP/YJ2/Qa7RZ0gCzpeimrrInAUaVJdE
ioiLwx6getGsd1ZOG4QTajf25JPwogmnvvouctKcW4Vnfk6KsqzmNQv1v5MYtre1
fRQlBbznYwIn4JHyo1SW+TVVV7ATdNyfiVJZkga91Eh3lXOrUduFQRtWQB+0bOif
S3tRzW+692dZVVhr4I9+SAjOG0ie7oWZg0K5QA1O7SxD0PWQA9lJgvrvGqwTMhfr
ti7RsUBTafOxFAuQCNiuZk9JHjbWlNsENe8UdGjzewqPrXmtYSzkFUdxMuz7w2CU
RM0k3FfWWkObLC8eAnQX3trj1TkXHKWBN6audiljucHn9vcBIN1oxgoCx4pLvsaW
zbtl1zN3wt5GjIbj15wGwZhUieyEJflFuZRGCWIbZuhIO/6DpcQkZHx2fJr02LUA
+5v+oVe/daUKCZOOF85BOtzU6G7bmSdhYdI/WMbx84G9LVGzrdkzPATDyAmOxh2H
SU8m21bXx+0dAEgS7XxWYPjcEAGiq2tyvGDFn/Pai1uFDYTL7ScFzVENbM+Wk0FX
CUdGGF4IcQA68zpRwnDFnbrqFjoQ6E8GAjZKDBQvAM9TuE/nycJa00+Mza/1mARC
89UxiSlxmyMw5oRGdWy85cMT2QDXpJTJOGaUTbyqmFFHI3fbRmHqbnrf/IpK9HiL
enLVdTz5vbXkoA+a0us2Np4QLmdMJvoLI+vOCxyJJLy255JJhI3stclajbNa3JU9
EEZI5P04uPrQ4bYBIkJsjAfQ89yAH4yK11YEjlh4jAB+B8ZHtUok/To8HgtrWL9i
k56QUa6Mv52h9Sr2U3eM7EjIosMS8xyRJcSa8l5UGsi0Ig79NL51cJ/Te+TMsj80
swP6BsFWgEBIaofDqDjKfDtA+a2YlbL5L+nnypbKwFmNbVvLwh0n6kPpO/AX4AWH
WwL1VEBy2iRO26DAjXIJdmo8q4vKd/U7gfDwQm8EpJcTiTO9O6OJ+d6VKOQIcqGG
KasUdpVrnhOKMwvCC+NZ54+x+fkhIRqtBYuZVwU3hPAQbb9oQCHmntf7M2koTzTt
f34XDzps7umoJdHkPstZJcDRgiaYGShmJqAO76HjP+frQ5ZC97wjGFovtxl9gPWG
JqUruF4l7rGzTkuZUpkTDGEZQWHafE9/oNv1h6a5rUGZ3p0CQdNJJaFN4egUa0qa
OL1K1aTCKZqaB8npv5LWOucjdzHRgZJioRXOUqfnkfiOwU8PrOtjo6WZOF6y0Icx
YY4pm8aWJsF9gWpikfZupo1PkYdC93iPrJqbmuxzPlQpFkCJ+Y6oOkmbeJTTRyZ0
6D7IDDrcDXP9xQ6olIy2dQD9gOQw3WsssIenPht2F88QZNqvcNRtuIwCEtCToLBZ
ca0ykyVir9GHTsW/zxfG3pRo9mgR/JNSgc2mGwAOfdMO1scvr4jZaV1mAezzXoMT
XTJkGCmCQ5/Vv6rNa+L8t+tB0e2tNd6QAolAbxhG5CZUZv/5eqSvl6/ifYVQImbA
qFPFTuQXEPGiy24Y+yonQN5xMFj9lacoFkI75k+Zb1Ugbj1vPRRvZolU+86xsFsE
73LKTk7FUd4WP986RNcl27MBTxID4nfgjwhhUFfCdyWUsbYjoUWbqCNZj58ISvbz
/sUZ53theyTZQOpcf6n+iO9HeGnkkWwWDBJ6Wv1YRdC1IzbGaggp6TeLdx9X7pEg
OOc01OJdl7qXp6zw8huHX0ADo+ZtXbl3o4dhIghH6Gc6MxPYXmzoQwt7uMRdUx3m
PRQcFTgTmbldONZbmQIWYFzS0Ux8TQ30AMiVB4SNPtE4LCzEd1RjX/grwcuGBlnv
tbTxB/ny49k+0f0/UK2S1WejStO4fFFx/NNBR+8og2q7hN/1rjW1HWi6uUIzlr0T
0E8rZMySzdMwUSAYNOvvSqRjjxChQ1cnW2sy+UQbCgEkc7NUGbPKQr8wPpH6hyqA
E3O5YeDZVjtpkOF0BVzawuEGE0aREIKA7gZUNiQp+24J/W30VOSTBx8eR9Iecyt/
aqaYvXirJBqjAB1bxNR+29/y2Dup5rnZioVddM2CO/W/RbkiC0ApCIR5yJY0djrc
k7wnWevsTnSWY/Gc09BwmgWMVyR1X7sPOQpfG1J0nFAUCihyLbOTDhMJGSDpC3Uy
9WSMzTFJtvnpoqMXAPaWg068Q+PXBCPscxtxwKfJGB4V/ALhyi+RuyTjpsnzm6gS
dYsyhYagBkHaZIV0Rk2/goKZW3i0lNNk2anwuE/kDg4nK305BFAMYIUFtr67f3/v
mjAVKmrWErSVPBCfQXThsybM853o2qhREnmMjB+I1LQ6nAZ9Exqv8bhZjC690Q2t
fCijlLbu5GHItUnWqqiHOzbADL/geGfn27rfE71b3voWX2WC5e3iuWGUR5ODd+Bg
vdJ/X41KD3BB4UVre9Rud4b4jND9aemzbc/qCdcGp+fqxEoWzE2QA84zMQos68GC
J1mbj1Bs74tFRaNSuorhagc8IfZWOBA8Jf3GOwP85pGqXXLbPqM6oCsN+Pg+LPY9
sYID2MCRLVB5taIVuyGKiiFUzq0PDmunZWGh2voUJ9a+motgs2dwzvS+1EwZhf9G
2UFWRl+p7z20pKREI1PoRNlZSnYKDUnewBkkjiWxlTSZvwlPvBLZmavSq9PF6hP9
H1ntAMYWinwMyn02gmL5Wh5DRti0YfiF6bMzZogxODY9kzH/GEPqvwBruhapaalN
bsirLqiQspBMPoAnBcaokQuCX/f7O70KCXQhImjZ1zEOf/5EJR8OmL2r7AbosTyY
flvYOpxBlrSHj8cLeB2/nl8VU9TdOfY666j8hlw4kZ8lYWmzEkYhNdZyv4aga5ul
NVf9AT3wCfBhQXChGILI6du1MoM18q6o4yTmCg1O9shiY24orH9PHX0T2+E885dC
T39KNEZjfa5YvQOAjUeKhEo2JKjZ2Li/HeEAjAM1li4q9t/inotVDUDhc0nG5TZi
ReqE87PJQDytfTuTT0XR6lyPQczuASHkWwYjO5mYiGfjhgjG5CfohLNjXS0nwUEs
swm1b0H5jZJvM/XL3Ms4pV2W0qJYolDHZ+BEV9qjXAgz2a/yetiu0nE/jkepvqPW
6lW3mWLMoT+RsGqEP05xMxaIAn5kA20ysJgLkfTf+V0K5SuduR4E7JmV7dktMlFM
VBg5OyQlcphigpr18q4aoDW2vD14zYnSVvzPHDLFel0RnPqI4AYxy0GrGAAEmn3Q
0Ig7suBVFHF2YMxWnYTcFMZj7z1HhA/8q6+S/R+f1pU7fZ2fpNCUAjIcTSWxM9ky
JPcBTtxWv54s9Llmtfso7BH0C5U5Vli6vStac56djbIFvNInIgPdde2PtcYYGVcs
0wnCDXXeoe9xI7J1TDtWLsT3yKvkNstXV9qNncSK6gHqTcYNUc/7zUs/PSIJXWt1
TfBW0RM59K3ybvReHv4dzNxpgx6YMMz3W3oAYLaacyw/B3kJ5FFDMXiDJL2gdyzU
cRc/vGQhNn6FAW4W6Pz6lpxr3rqaIUCgTEzh/uWpXplcms0KI9zouyeL0y56zO+m
jvAhcpzSiBsjotTtXIhuaTysQITbAZ5lIP2ss5vWy/rg7ARqMJx5D+CY+lAFS0yz
B6djekcyrigwylL8CCU5BSLsk4uahgeidzcG2KfoXthyRegMD3vonqaMUzUXXTKZ
sJl5zdAjxbJlqh+K7jBKJtvCCLjBet6rw/tA0g31jsENZRE/km0ZFK59pBcpI4Cw
+Gvn/Tx1Enx4uX3dykBFPIgqVgy9h547kdyR6Ewm4vibzWkS1kQP54/92GZBhDfA
Lb2ZIMIz5Fj9udD9liBGYJDrU2YCeNMlU7u2LD4kFnBAuWqFygyg2l7TMGjgXnKB
x9WAzt4GNKD0+p7LNNdjUY/MKCdnka2t+zcRNOC7bmLBiDdvN8qY+RTbZAccI016
uueqEwmINbBqmv/cvS2srEIpRyRsW0W+6P1HX+93+sjgcCGPq4LlTI26Xy4ym6K/
j7HYrRTQ3XMDYCMoMGNjlQbGA0RiyggIajWexl/pzzZUvKGoS5K/sueqpYUK9LVJ
78iJcTBB9onnIO1ydklNunds7+Haab0ewvvb2YCa+VK6jVDZ1Mqatc9r3l2/RKd1
J65ZkXaL75BO0KMNE1Z8md4Y2dYcAqxWFZ4SDWyjzIa2nhFUhQcTQsljfB272kEm
KRR63swAwqaUAi1nGjNrjfImUXsjBXZK4oDcH+RZ+CefdNhlCrony7DLxZ/fWkq5
Xa4MRdVyb39aRhHmUv+pZwsNutQU4WWFpBmxywiJxQ1p2v6jg1ynMKwrY8JparJE
vDv9B9KMGx+UNR9MyNWGRQVA8kseoBoEV8FDHm9gFWWH7P+Isv+snIdazRm/OmlW
3novbO1Y276v1XGqtwIX3Qb9AK5iw1Dci8NiAmVYHTVSwV/1ynVqSmuOQOUvrqHH
Nbt5IPIeMLPrf0Yswk1SliS4T+mnT2Xp9A2f+PVBkEYh6pdEmgJh7qGnTRsy9kOx
G/jmUlF5HcvdeIatDe+wMbu85g6Ceqv0ZcP2CYrmpDhUA/2QAzyOp8bWC+Wj86xy
TTwV1NLPcCra94iNhTowZ48h93La43nCNTGJfk3nrI6+9bdQdrIuACKs+vwLc1Kf
kTVhY0bNgqxvacCToUM8pT6nDyzDsEXFw7Xhir3p35LWjCURO5GMgIC0vgZorp0z
LnsakLrsmbEcZyZr6Kvu/fw+xEn3+iXJCopSRYnhwTznm+NcZKCaOaDwvkOb1Vkf
hUvkzCJjeFBea3hXrbRHyLBxnPNSB+zhUtKtrc9MyoMjH18jFgd6pB1VRxuSC4tW
CfFWyJSBj/f7oOk8hVvV+w+NI47ivxx1i9QHLdCiAlPQJTkwWbBt4rK6RtbGyLUE
ydPDAn7tjA5DevHRbQ3kWbrs6lh26RmXijCZKexSext/L5quzQpzUpShLwHPoCwK
zfkB6rH1DxQaZY03ChGzwLfVXzy15oCFwLL3Y0omz1g+LavmwZiz0QzP7Lt2Z5BT
tTqylZpPu5AOdBIUI+BoC6roLeB4ccfuF9uZvTTCo+f8hB8BmsYv99nmjRF08lCu
jSmtXuMC0mcRySnnrUnqN0BnF5sT8ULeqBw5dduj1OBD4lbY85f+mX5dg0m05WzY
fXh7DnPQAYK7TbKKTKQqLgeaKXZw2EMPM5P3dhLFMoKUDjNeleY8WbsImW397yOa
a/5t/dJMfnUSLltWEiOREv8qi7XTSGpaRF8uhlb3F0arE/jGrKyBI+mq5YUuRWTK
fTp7m+DiGPQLITLp/GnEoJA1XdNrlmYB+FxTls79XdqfdPvYbdxVglg2rIbGVUBu
82uGT0m+foa5jX3LpYvepoLXZwMHuJ/sjtOioOqV6dWSrpKNf/eXYPUvgA1d/VUb
UVB0D5zy6G4d7Ce73SQbpZ9cq1jF3ntDGKxnmVHvcMgwF6FDUacYMCfTpPs0pzSl
fNLies+D8FlwyGh0mPEqUs/8yz02dHCfnhIMYk6whRg7LZRlimcq06haGfGFZzg0
xjdV1c05YPA5pR9WHSVGfS6GyuGAP1c6jqG1gz7AwhPGx+rfwFhZRM8AJZZeYqE+
reQ+FX4g9sZUBWi+BBbm8AJIK2D3lvFH1I/NxwymHueCEnZhX1qJV51pWO4QE+54
YG8fLHENJI0ICHAtCR4qfxuN3UEQYKoyXTGgDZ4N6AuE7hpHu4UcwuGZOqW6Rb4A
rrp9SOV79fgHFnBtAK34RZ+8WQzk+gefvblekZiy1wTPTQHeXjglqh1T+5MUkcqL
VPC1YDBHpHhZXqhgCx7IBvB7j4ODgCTWSdih6bAOOCnmPB0Rorz5X6T0XVqENk2X
dhg/HHCOSeD3idNIJNW5TgOL99W+g6H7jOKlhPnC/U3jWby11b694W6i1yqz5sqJ
B9kY+BM2Kj8Ya66UrG2xZW26cNStAqqjq1Im5n7eoGOI1nH+fmiX363CFlLKOmLs
BHbeo3HfY0Eaznzw0Yvm+Ct+MXdbs5ZG3QQr9ZRrOoe0IK0RdGCotOF+21n68Ef5
rFI3a00pxTFPTfFwR/2G+verZy5wYw6wqZodrAy5N7mWyInC2U5UqF/zChjCuEPP
YXZdQP4vK9BAN1JxG+q5dc295EItlE3ZkMxHsEoXLUOo6L0sNh8xZ2ZRwkdr2+w0
v1+oUKoJ0ASDrKIAN0TSwPsQcD+MtXXcA5RcrZp5Esv6riFjSs8Mptu97hgtLlOw
osa9IboRejdTfLuRgggND/P+/HEkNwtLxI2BZ0cCq4am5j8gQCLAT00IGQF/TIAn
dLKOa9O3RiyU4eDcStuNCzQP/8mT+qnx2pxV/4hi+47c+xvj337HkJj6tCkIOWmz
fuc5UUwn0/5ijB97y6+hvdDnZUb98JKw+JmBge133Yy3Kvg20A3TQSFjbvKXkvrT
xSUKS+Czsb7WuVw3gPP/PKD1NjKij1dIJPABECqzC1uA0y9HnUKW87ZTccUwrC6b
Du1+0fJ+aSbRnP0kSJweBXoWPe4k2xMwAdPKvtjDtH7onCoAg499P1saefFCigw/
cw4IrSRPu/ed9ZEK6xrAlJq4Pt489so+uu/KmRNAWLG3k1lnRemp2Aov9luqJjWI
6plP3c5Wxo4u10jVl22dXCOXpDmZ5/48dJ8NoZybhLjGHaLhvjKb/qbl1xR8Iabq
BDfvNcg1uDKSEzrpoGK1k0Yii20LNw49OU792vFFpYWxhUPUb3iS6YICu3PxDzVA
4rkJFfa5HMny3+pXz/VMDk1t4jIl5Tf/OBmmJoacyvtLxkPEJy3oMMMOXObsL57R
s0FnR3/2UUJeKF/m0J9KeTL+3Rz/bneka+DiexWRcVl3td/CxD+vpoBMFeY3612A
Z3vUrX6b+prY5yn3J+hoV4qtO+UN6UH4Tf+Oo2sQKgrKFrovQ/ShEWZStCPKIOQz
+6cKFIxs/xLzrfT0GoEEIFtAqlulDwJ4mt6noJGlfRF8d0V3wIGVD7ysm6iwsBjc
BS4PZpONUd5YRpwGibj7yk5i4WIhrpoYC/q3lAmM7JHNFMbM1XjUZLPB+Ftl3gY1
xO1Oa63WbLY2Y8TiEhSF6H20GoY1Y1WoG/HBKVsh8JyTbMojehHVnwEewnwzauip
XGvO+4vZlIeqLld262qTTbJ94OBSRGml1IkCQnmOG3E78yKRTOsGGSlWm11GQ5IS
nQ6ggTfDqz46xwq8iUbLbAtYX4bUTv8igtA9Y3mXQOutq+nYvPdFxMlzD1N6O7wN
L7Mt4yI1GunWa43Ju92/SzDrM/5Fiu7mV0+KJL63t/mkwEzRiKWONLc8qF17fBoS
cwXyvStOgimIL5Em8GtK9Fxg6iZfmleSuZiTLhK/rMrpfumoLY6xRsAnoGgZIiqX
mfRjMLCc85hi/Yyn5trx12Mt4rkvD/JWMJY9Nelc2focK1Mmfa8ZddCFQKdS2E53
NqaI+2YXh8h+DrVlmM4VCk3DbJ0zHrMrMdmUZypYmZUeWI/Y7/ArUaeZdxa3UEaR
T0XA02RWrUmexKsRCCFEY+ZKA1zJEkkxTby2y8f0fr+9MGuM+gQ7tzSwQ7Fct6yk
mYbmDlwpbW3jwznhZeyAlImtc5R/L4e9KIFjNYHoCiquU4DxdmUrWAOmpIYiu0gJ
jzsHFa9tMeWsyfGpdkOwdof9CEILaBKdP2mflOaaZm0E09u0js2gW4HHDk2OHgeL
qInV82QilJzl17eyoiQtjYrk7UQtfmFFfKR/Gfl7zoQViWwao5pdnOsuaA0lYos/
i87wixZBeydY8YVuYw8hY96WjFws/pN40vgB6fJUdRlyYhSZjM7SaSwQMMoHBwvt
80PDLvMvxtjF/avXmgDgCCLTtjv4cqpOBgNZP17VlBhSomghCI0aJ4BYycuKJ7hs
JbBJKsmuF0biHmWpsc4bg765JM0P1mnzbkDQdb62zTzaTLX1pH21rQJD/ZJmjxIK
7gieAQ6M1W5HnE23oOYQeA3DYyoFgsMdvNZGOtCGZq160twtyRfMUwzZjFj0QhwN
uPXRoE2nRzLmICdCOMMVb+gAq/3lC8duQmBD6h0KFGYU9hnuukYfQ0TQdWaquRzY
znc/NsoFlxYfVuNmE0E7s7YgjQSC+i2Z+WMN4iSP3j0nzmW+lQ1StnphtNuoIt4O
vXwno+MlM3YzrfbgfPCVsKxPwNVeDFdFELJ4MIc0KZ+z0mKyovu+dXhLIiCCXVFo
4HzdWy0Zyv5ewKApIrrD2JrDH6YvQEO8HALugLpbofJ5rl92LNFtmAgSh/mezem3
OpqXxpRPeQGEBkTpJqvitxVI+c4EAIAgFAG5rBRVkssXvlpy9ifK24lH/RSWomAz
B2mBMvk8BTH6ealTkbcduNLtHuoWXLrkYlveSabP404yFBzPPbXtYAfntBhuSMGJ
WcIJry8UtiVcSaEZu2IZW9ciXy2q8pWze0bGkW+v0oVsNCiDocYNnIItbSlk8EoQ
sIibdL95ARONAVE7txd17mvbDe39KzViwNdoPfWTgxorccT/sLoOLHwChNp513Iq
gdRwsJgjcMqmyByQ9dsXeU2M2ke8kt8WuEp7zi/cppy9fAbK/PfbDWOzuYSXejXs
x92CVo3xi4qnyQf4SjZB4ZuafASqjeth8kU/FVKl3Y+QeGxiNQOmf5Y3+/Qy6E/e
OhU0O4kjG62CWFbJ1CqGFwkAbvr3IVFBANmEATlebZQBZJu4h2OVE0EQSIUS0HyL
/Tfbjj5+dxu+ywh1LPuHxnHxGpd1yXNfeFZ7JgvzcohKRicue4f3yn+uhSnf06j4
uno4SksjY5Rso0p58EUg10daddufUsTOpFAuPQ4EngUQUJ18Yafdn1djF+Gx/0Ao
qNNgW5rJW9Mu3qEujRGRwvVtPzuUqUwucja+jbVfGC8gG7WXIneEFcgt8lSvxahI
mRFsfaP+eW5OuHXcJzXlCsQMSRn1pXaeotdZk4xfC4n667p5cMe94lH2iZAicD0K
GF8bfSnaF3dcBYx3NRbiwM54skL7Nc8cWG9kEoiv4uffPr2Iy8L7MDfpIhBjf5Us
1/vPwKr8irTfXNzP6AM1LA+6UJrCS3KyXWgW/Q8RzX11COkw9TrSMWbyW1rH6bWw
vXGrTnydPzBeASCJAKo67EYylmb/Juqnx3+oPPfDlgjFezvox6cskTHR7ld+yvJe
s0SSdeQiZuYEsyXAVdQ9VtsSvuPMIoleIwNA8O3BMZQCqkMoeP0Kyh7VwLGSr85D
6tsZaR669inoQ7VzCQf5ejJG5IuV9guuOkxXe9DwV76IWOjtm+PRXoI3LHx1Z7zl
GH+lqV7rf2LqZ69lpYzfLV3gy6MZvKqLkXjjgLSBLUc3n6McL2FbbLsSGHUEZJu8
eGP6sh4V9W2M4HMXB/KiEAkuATEKK2fLcBSuqqkRjYZ9xpwEr1ePoOw4mCILxlJ8
QvbH9XPPpi78VHphB2ca698T7Q9x9tsa7JgNkaQTTShLjEYwdrXcso2ZKT5teFel
2ySr/aotsi05bC/lZg7Aw7UqlU7m1rXh2Ig0olk3WDKj+Pf7NZ7L+MDlutmr4ldU
uF/uBU2Sq9ljkebAfcB7AGKuF0auEtPjnnAT3aioMz9ToPzbVoobI6L/CHYZDKZ+
D3larU4qlq+7YnyQKw0W9rO186hA5IydjNjuH98iOj1xE3vuFE6P+QthcKwyceQb
G08M3kRITFkILvbHWv3z33LAQwx4SEhoTQe1vSizkFMlMirFpabBy1yBtG/W4OZV
egnF3Fr1jbgHE9Y6MFZcAqW577C11U+2JTWXs6unSd6RkN9g0Xmpp+QSj4xN/j5O
uby9pd+8N8X20+OkMnMED/AGtSaE2RAZLKvo7Twn1IKcEyB8S+GaOffy4IfsbZ1J
e6NyiPp5I5sP4h/+dU3qHNb8JuUvXCdjkxGiJlGXhmmokyBWTOwKLOGBfQvL3nZX
H6qUOy2gp4NjjKmVQWWXaO7NIFZYu2V5Ucx6l7OM/o8bprT569647WD9ubDUCQkv
J53DiKlZFZDnvIyQFChVthplIrL4Tc641O/usqfCT1DiSzD00KfWaDW3vnWjOvJ1
Yr9jM4WUTb7qEOmsWLm7sEaRMkKQ3MifTFgiKPMiOKC7qKI9evGLHDDEmlsrHBCh
wdbAVf/sDzPaUqMUugbLZ4XojomJEhy4DiYrNTAgBCqCCQhzb4vf4MyhlRrj3Qfx
lVJf/FvuEKkslKQDW6tm80jsrwu//aFY47VXBEZVznThOoyAnUCgPvrmi9iXwj0k
dy/16yvRLa+fDjW+qvV2Ql0Lsv7a2LKl43rqxQZF92VaFHcveGy0PnC1G8cqG+N3
DeEPAImgmF2+2RR9A3pkUxh8e7EXn+TjX9Y4G1bdroB1C8HZt8wi4Sfg/WbmVRIi
g2WHbhFk9okU2r+YbsVi9AdLPa/oK0znmXms6U0N0FixDI1UrdV6EnCap5FU67hH
lbq9HQ+JswL15phoqzsZT9vx3vWnAhBw7vjQWH7oIv32ydOwexbRrxUhsZHXdaMs
TnYPgfBdwa3KtKh8ZXcxEfdojGoBbcht8+Rjz0gIJjWtLC55QsAFTFj4cDtNxQNV
QQbIVeqraKdBSGNKa7mflr9DT61pnzOejsyKf6tAGsNMgLG9jsXsjwJzGBC9wYz/
zl9moPaVUMlaUcJ2eAKPUggb2hKuXHY3eqkoXUIJNtpC9yBnGSkPHNDoRN2kmeiI
nEI8FrAMN02Up4/vtmhYuvhQI46ZVCNDofI890dPy+2Z1hQ6WSoSWYacwbL3Babl
S+T6HwkLKHPqqDlBpa+bfQs7PVpYy6Lzj1KoIoRYf+ikPdu7V70ru0HC8CQIqMDL
cXOopN7/PN47HHFRoc/dEnEri+2DPoMQuo5e9+relA6APru1BQBS1UdnqL9H1F6b
k0t6JB3u0h+0N6Mo/3nPx4+6PsZRiG1BMGEochUcpwewCupkGXi3s6H2j5v5UKBW
GHoHBIilgLcY7jMGwWnlx4qr3FUjeJ4PVBLGybZKq48y2HYmm+hXI+jBvi/GfYwy
lSLUFCEtAeD2x2KcF+K9cV8eVMVN4cmk3kwIdpCy8xKfz7a1rhcg+0UCImdmDX1G
utwqEcSRddnAiX7ytCapwaYOyV4FqrILx3vlx25HWBEfMapazTxoufl5etXrFlZz
70zCy4vS71PUgDGevEcrKv7kzlJ9xXEiWZvPgH5/XBJ1OqS47AY/TwAM44vGkEwL
rci+O2zbdGb16IZbO0l6yOq1ZIklFbyNnizyMJKFby8/fFClJ6Luf7DvsOjgsj2Q
Ats5qhnxP5bm1dt5gsI56EnrvbuK5EdVULBRBcbIZLEAeZc9csvvYjm77HP8wYmK
eDUvmHlXeLScyfnGDb8BcBuF8x+0cFCwrp6oMUE7GEPBmZDdLtaCSmRprSWawVb2
4JfoGB2aJOX7hlKelkMVCWOd3aQzwldEzqxPJ4iiccJ852QiSVucVelBYfUO8GVG
rysMuyiQCsrtUQi90lXqRjL0YvTZjsx+qhLFAAAPbMg7s7hwK8YthbwailIBWYwQ
Uc2uFGWXf9Ye3UYg6mSZFf5q/t/byfxYGd8gRO5OGKZ5/bZfYjx/xNJapMuWGGK5
a7TLmv7Y6bKcE8D+CObXETWY3TgWp4Q25HvDxga+/6goiKleAq9f537Jk/dnXnYg
RUNxbbjezniPGHHg9xjbc1RzLFB6wAD6i/wpgYqAkQatUtAdvX+S5pihTGES4eCp
KorIgxSaCYAgxR1yFp1fImmoBR70p4Yp3JGCgBE1TvST04ok38hmzBbdsxOuwBIX
NMsUwk/CmnFSl1sYqz9apE3+PLESmJt92olhqqqYzFlirKeo6S7fJO3O/8c87v85
iBsj7RJC/0up4+RJYr8DuJK1AeV9No/kMWNhm9x6AkzBMUdxoGv6W1cE/Ob5PA1z
RgfvPJLkbzHTvDH3yZQCJaEu2L6kFHiKYELft+AKVnLWhMgHphCdLgIGW0lZicLD
PGdzANIco0LwLvqnCn7sMV1NX6Kbg3RNB242TJc65Jn6aC9yjqCrm1BpiaB81Ktq
tdyzLk/gW/RkYmJaj8gGoQKJh24YOk7b1KmNJ4W1fy57VREue9vnIeFyWaXu+lrr
WfFoWBeTlGf2BwbB6rbhoh7Wl3K/GF4bzibto2nlS4IYaNY8P0dBld4TihM1MPfh
rLm2QffDOHpWQduL3C7+Pmb1/hzqSgt6Mrl/TNNc7gSsHvfyJYQgyRQ/hAyePgke
vKP3ya3uqDnrLvbJHM8eyykf2rp+4behJR/DwobkS7vmjdplW/Nh1MYq8bE1qL0O
KJUAeZJI09jqwfVOS3uYDHhbELyZhnFnUppbzd7UmmbsFwZZlZJgl9WO7HYQS2Dw
DXkeonR2ugkqIlAUbE0vbmUp4iledUvJzQaCP7SCa0K7w0e4swQaV+C9wDx6Cp1/
Ql7OCHibsV06qoh93xhDk6Zpkl3hSQjzr3Otg6gw6Qzj/2/oiRY0rdUfX9FZLW45
ueSmQmm3vWWjSYZiar2LWk5bBu3kKd1pYuR6v7Myj1sXUz5c28gwvn7CLXxhw43J
V+mSrlwbJgkGiXYw985LkozgQcBzH0AwGfecVr+smv4mxC31dD8X9vomU2pGOwiP
rBL1qDRXNVlPlNdvNqGFQ8/ScxYVXjYevpimMeNaPwiSXCw4DA/3+RyYWwWwGV/D
g2DTg1z5HOVve1RxMlUmEvopLMy2+KKqwjA4rYoe6IHocBwxe9uQh1Oa3DX4BIHR
XfifUZiQ+wbm5lITK4cKRzJ/QrDV1GeZ+6t7fol5f2WtF72ipMHeH09yhPZGng7d
0hWBOyBAX/eL8s9wUiHPqoIl/Ti/0VKZKFi1SgWusgG05urO0Hi9fx0othF3GMIN
QVrrSSf2FmBYJ2DpY34mfE78nglfSbhapXt68HRejmhxkcsJ7LsiT3aI7iSs6Q7h
96Vg9yjPip1eX2dBX7ZxMgkO4cpF9V/L8MdLEOILih9f929sbiJ16YLO+L7AJKkV
SgxDgEkyeBFkPjVVpmVeJGcgKsTzz7mbNHbyUz2hGmKUlDmcUWJE/qfT2sJCH67E
9dM2KJPX4ekzEhIEndDeY2jImZALQWZZdFZrPyKOxRavP0H6RCQLXfR4p4vKsG7i
HZzRb5hIfYYoKPGNXNE/6d9Csrfdy9ydQpCECnx+iyLGIldccabCIrVujIrmSejc
NbC9XW/WyQaFnXN2VBUK5nGzNgXKDPqneBJoKXuGhyO2dM2X0G+i8Hcax/LKm2jW
hkBO9/rQfImVfsxajLYNRVigzQkzv7W17+UCNRqEsJbKG+D7FQBmE69l0ToXkg7V
uVtkFyz92G1YpxzscVFchBypYTcHfZ+5fBesTvnzPCgllVBLLXSp9idrs8/e4R0R
SR5uheJERwNB901QCF7zmJddMHPxAWNiq0f6TaWI9wjxC4onDSwJ/LXpY4q8/c3R
NtrIv4twhgukbEjpZ3FJfKEF3xPTB3TfHKrKIQoKr2bngbKv9ct0y9dxkA902ixh
z8Av+504VxwULfgrWHtYuOE5A4Za1unNWaMRW3rDcaPwWObu5XkqVx633ofEQiR7
XjUO9+uGwo5+sHpXFsG9xUKXs9JI1gJY17ShhIUduxfd80Wv0UlIZiueT5MJB/vS
Z0Nv6gQicGnQU+VST2/mdvoGxwpEkm9XsDvtHSiEmGGdFrBQ60+6oBMilXSB7h9R
EDycIxkpzfF1XHvNg27nW863u8oWeWYYtzZUGxUbIYSPg6dhe+RGrstUPd4mdE9v
ddd1E3nh1mT1OkNAqxDmDnna6cGHDVtr2pFFroYD4xy2jabaSpp2u1sN8+Efum86
2RZcpNJbbKUh8tp3Xxwkk3VJu6fCKlHD3GAneKA2euvcKm+y5lP4SkgWs6v/PauC
0hHEVqAFF4Z/aJLPp+D2h1Dm6Pase/9b2FFtBxbiFHnoBw3l8NRfHdpq28j8zLRL
lQ5p/zwUgmFc2PrWVh39FIYbQnm1ut6LRAPp3B3ZXDxe0Zr7BqS8YRwQ0UFwAulH
EnB0dyk/WGt+KAe/wUoRrZMWNmWsFeL3D4W3kCks66QSEahulY19mBLE+FVbkcJF
xfG0oy9H8VgPMfLQ+n4Xpn+xuFUVlLH5KOYU1yy2s0GDrQK7us1CGbgEJLvJ2JsR
P7PXL7mL4xZMSlgeY8MCI04R6X7hEbj2Oha9Myz/AoNbPW+FGbYr47ZJdmqybCDp
6jURmijpFSb9iR6USKb2B1Ek2IELSGSLXD+wBbLdYh0YPrFxPfql3M4ZCv3ag+Ot
iEAm1hodgtXhqQXnVUuch+tJSO2csXouLy9dmeDUZfegc41IVC7NppfXEFk+uI6o
+qvsChynZo1MjVlFueEb5Fe7ZKWssJdsdqdoEuA1qKRP6tJyezdk54IvpGK/6IRC
piTEDy3kFw6iol5abszqWP0+UAOOTj679NRKCQ/Md0uvdL/hqizajWGBoGheqLNb
jbPMiRMXSysq3QRnRpgrI8XNMLhUn+BcaTRgfHZpU/sCbXyMeahbv5jDTUNuBT3B
p5jaoi+euoIAl+8cb6Opa4xkQYP3GqUQFGc891C0ntAY+HllTkM5zlc4ksNBtJ4f
Cf0AAMR2H/4kg8qwIQ6oW8kbPR3XkmAoIMdJAJdu+JfEcIWNKyrDSLROP+VjHsrr
YWPSVVk6n1K0MdTjGvDOkcND/g/PJJzH4mLRtQJM/xwmLB7E8Plbrj9TcuujHO7W
LjUWuqOm+liD8aXFlaX+XPEv/hsJY8if/1Fv0H8nz7lVDPAH5SvMCVK0a1COCM2J
4TXjGGg90fy6bL57cSCs3mEe3f2nWay4AEgTIjXpKFU0wwBo7RejxqqRgbgzJrh1
0BcBbEY9FPLuiw970G93f69blfkMOpB1jj9O5BvysR3egfnFH2OkCmfoIJVkUFh1
eWoJRvsI5AZhrwydK5INteBciRQDTi5ezn1+cahTMkL7pNK8TCNFh/GfgU6fRrXG
JoRI5D00dEzOj0PrycDAHMzOSVXVHl7YswOIsOnivQONSKu38uIUAHmALAtdNln4
QdNaK0fqUtJU79/suocY35jtST/7B3pIVj6XQ5lWriTySTW2T7jN7HAi9EjkdyhH
zuZL2M7sdPEo4qSOY8AeS6L03JJjYOs6D6aSqOt72Z9EurkgmX5P1OkBHz+Hw7RX
XfUPjusqKzmCyVtzHJ3/8ljoGjPOejPsbCsB7NMqsOz2CfsZ5BndJLBlPNANsv1q
y4KS3o8oyOwvHyRumcI+seS4EsRamjxy22mKgkyqi+sXGIn+/XjjUOSSP3XO5mBx
tLArHy78PXKsBS8gNO/PVzsBaLY89Cbf1t8qoGlHkOPlUKfevRG72XGH9wxuWQqv
owFu927oeUhgN3PJhn1PR6im6+LHTPLdRE4YppY1R3JMOO+0GPbP9bfdHFse/E3Q
Lfn37H2qpq/nG5Hsv7QIanvASNFDvoU5mNmxQTPpFM99pTd97dXKxe2H4Q9NGN6U
k4T9hLrQb/kboYwBqOZORovEJWbMK+sbexB9+hJvsDr3zDfYKufKqkEfFy6fyFIP
KMokrIHtSmleRUU3AgZlZmqsHzvONHMqU90Epx5ngLO7d0L0Gf5ejELF57wieIAj
YpBWVgYOR2kpjmv54A47/C8TbGE2lWcgoLmjFGsKXBH3y0VuyWblA+hYxEiuuZ8c
GkPfgshCxGpSy7cYgKSizPF1p6YeCAuhM3yYiCX4Ygvfd2SCPmw8qg2sHU1vptxh
M0EyrrCVyEQoK0daZ1c9iTuvIVeTEqGKp3bejFhpYaxLLxXJvK5v6q4gt59FHAS8
wP/GUBwn7iXOUPJDxIf4KB4FbwyiTmunn1CHEF/IthkAnvc4FB+iW5E5fi1dhrwt
z7JI7pdaMzlbNmSTKkkibXLul/5CDxHDf2xEJRN+1Zt7xpW1wXhdgi5iKhuzb+Mu
849RqG4sI3oP3BcF2R3Mow3kXYRkr3tFrbOuAIDnl9sUDj6iNUeOmFi+aBhartrm
fScu5j5nv7oGteSOZ1h6zDm5XjxvUGYK9RMiacMa6+fIekL1Yz7NK4R1HuvLyHCJ
mhRlXli0meB+3sRKKtpxj5C0ZhAgSfx0pT53aFTTLjnApPIRsaZ30rEoFnlJuawn
mfBwi29t74r4ppAgob/j9F8DEQZYlJ79Hn5sez8PLk4MZvcJwW6d0GNQnQW4TjAp
qkda3BNC61LDkL3trGU5B76XS+z/bMyWqYmGhoGyaXs3qstlPnXWUZ+19o2e5OCD
zmrZReaBvILzPai3VlmH4dw/B+Ho4uH+gTdulNEA1rfyNiUQ9zVQXI/NByTMstIC
tCZbjHhA3Ux6NW3TmkSJZSBCtdF4uDV1F1ETVLcDxcyd7KdS/0J/KZucUKN0kDOW
5P9azsEX2ztM9MrfGWGNdpIpiGTxUb7v0+GNtZXQytZt93DNKXc+1n6qurvrz8mQ
UbY7yD3MRcWksTzdo8AdW2APHh5CSzBi0z5L1GbaOSR2kRNjEcLpYEZNgo3Mse4f
8FSf2x1ObXuv5hfDflZyRmcRsDwADayg6fDcC+TPpBG2n2DoYSrHsUYyYXxUjgec
UoZh3g8B5ZaYfugIAlU9pjN2ZZkTcc7QLGnOPfAa/Y90SeoYmwEHZ9Y2ZeoYDgg5
Gz+hgD37GEZyYlikDtb9WdWtMjfu4BG1o5Z6GVV/ul6MUrrfo8Y6e04QgTpzvejE
bz21ILxjPkDI4bWuFjzT2wvvIx+1DcFD8khHuGnDFtzHa5tu8jBLJodIXl+9ejPE
AipDbVfErEjGQCJloaUN+RgHJTdXasBYhwM9FAfeBgYXWDRkP0DQ/5mOzcxE+59Y
0W01ZwnHGe4xxxgR82WnTQ9+RDzD6Ou3ybXaJ3Q91nL45pRRBeiQljDUY00Ha55r
oZO8Wx6Rx5Fmb2swlkjHh7KI6IZ9yx1yWXP3SFDweTgzETvCOG1sq8+0tf1Bxlrf
QJE6Aq0pD8F5orYKwecUC10iPsp1HccQm7Wri+zANXnsWHJjBeflK+zEIOMn0nFb
JZ2eVOK+XZxVttgkpqj1jaShNE29t/yF53SYHldopFMwc/uMSzqq/YgPrpR86Ezm
ICXMsnUxwkoPEQUfs2MMpuYJ9d1N5ZeTbGtn71zpOXQT5Sw/vdfDpIGDvSBgZBkN
XVRGGUh3KZIXCx+4BTO0U+ZBCLQYMOm4ipfec0nsbK7K60RzylxKVrwC4hVD0a5c
IWIaffqPi1l1TXYQQB3kM9Rzb5/BGA6Few4XBFYwQPJH9nbv/bp5TXkFI2xs1x6D
pBLVrtVNl5zVPGohwYQDUkVhpaHyqxNeLyMGTMsrGOlYTYys9n36oSKAshnGmOcs
w4RM25L0EBRZ/edI5Dnjmer4XFGzGVotOi97BAzgrmQR4QrXsvP73VUo6M5RH2jn
IL+asLbaNcEOy4LcSjbEX0+YPi54urA7UF43iBw6eWd6SJ70GsuLSSUBvQRV0hio
bDeGOuvbmf16QxWj+lNG5OhwEZHZFUb460qDlk5LGDOFGRIj+pn7AZ2wpcxgjYqT
lIlwBzxtDG6BrqkxkOoQFWldoIpsyJfnCgi6c3Xma6kQot4hY9qOzOli7bjveDmR
Wljo0hfV9sasXjfkLNtyOCEqCM0JJZwHPVWtEBiQuvcXjaRztdT7mveZkg1SGgVv
iU1944pSyvct1wa4GqNku9VLBRzhJTRgs+nRaeguDWmzqVORl6ZVtul2x6pnyvRv
iRX6psJFq4Fm13mr5EblF4Pe5Q0eQuPtZzGKzfvwMJ86GHizPobvROtRh2dPUD0u
omVp41VsXSqMRTlDWai+J4EXgkTFrS3KWhCg2i9shNu94RmoQvgL2l8KE9Pgt5KL
Y+iTzqYUcBoR3z2zjFsf1xEP2sKWKALQPi2NHJYbQLTgsWkxjDNZCzEWKSHZg8ok
0acSJg6i85iy/41+bhRfAoht5aM3Quv7ktsv7ae9Y+vhBHCj6i+fsXmq+DFf5O7H
s1OiHNKBzzLMevvPK2d/FOek/qG8DFosvMJwdpi0zS2WyQvbEUSZ6jzZFPTpC/kl
kVWU0hwJf8qEpfzHHwc6VlanrwVOcCoc7SakF2Fl5GYdW+xCG3TPhHXY+6fIJ24z
4bV9n9rTNlNORH3bcaVe//BH+g1yBihWPvSjZNNEcJM1EW24Kq3625fhQWoHxXlb
qS6mp/SozNbjDCxdGUgsfG3+hSgQwtH9lKSoPbHlHeUPsDBGhtqe9fHHnmtBaicH
2dh0lk4NmA7XnwRXPe49D19djBfYAIWCb/aYU7SKmR6O9Rph3AOKz3jnmPWJ48EK
dukbwtziuO7W2yfFJ9ZC59imYLB0cEcFMY2ilQkZW4rMT5Yyg4zS2tBxo8e2QDHx
bq4xOmBAlP3ECabg18bpriZCMYclkRhBmmQhNXys48e8qY+KOMFxW5Sh1zFJin8P
2UeTx1wtbgZvOXQPl5ZJr6L+7PWiNB6S3zzwEoY/GsSLD+KFQNiCYVR9msvJqH9W
GajWrwACCQmrE2wX7sJj/J8OM4qR+ZgbIBTrV4Kee38vwi1OMY8ysW+sFscubIhM
jlsZK8cEEw3k7MfJ5RSfC/z8nL+hlSCyXTriaQKxC/99aBwEKjhMWs4M0XPbbESo
Ioeyqzbfh9N0NqQ8Fn0iSrD3K7pqKDM6Zin+FUoiT1ZBRbsZwdxzPfpKGVVtyLhG
gElBuK4pXXKoJQ7AHTEaFzuw/NWvyH7EU/LDqjhfyhG32UET9uWHCy4FzciqaUXR
pG3ISCfOIlnWRLvkn4YR9pVp/lSss9qIV9MRbpIBJ9GeCmVcgTRjqwGFVRG5o1v9
RuDx9MPHRmnbs590Fy0qE11XJNSzi5hrbcyQsXtdRgPN12/SHZaenrfwVpsZKx7Y
qIAiWXw4x5A+2eh0IlqhafRbEusiOoID7obDKPatXvJiGWazxvK1O7yllIE9NyHp
U6bKCIBEQvPzfEt8ECRRT4pKGGgtSzRH9p5WlKYobJ4t5ld/daj1dGjTDPQRoZEb
YCtv74jsAbh32Mzx6eHpjFJeQNdk0VgH622eh6x4ppBBlvOMD8BM/D/fzGLcuX9H
RLakoLXWw2vyCyg5tA0ooK09kBKlLta23t8eGn7uWBahhKtdrDWQxKAvH6p+3mwt
l7FCBlo7OdL6jMXWWYbpmKNSaQU6a/Dr3SKFNh4ubUS3/3weJ3HtkVG6zqC+w2t2
L85hC7PDOFI6L/oWTGXOSN6tjq3m/7M+ChaDkaxlZZ5osZmtght3czjsnsYwBwRa
Oz7i2AFTxU3DswObYSFfLnzOm1dxFjw9pJ/bi/dYH89FQXFSnjfjR5WHH8/d9m7O
TM+5HPgHw7Hrw2LXVFxk8kGi60vkP4gZjo0mai0p5JfM/zxdJeQeMawivHVPOOTL
9+55Bonk4liKZt+tX6Rw052vvSH32EgLmaszo31daM6N8tz4byqA4tIWQLdAgYnQ
dG4obINSjzoVCJSB9Y/gW5EzxMEtiFMsW6RHgu0PMDwlDdiMhKrG0VxqSG43S17X
DIXVd/tHDhQ8ei3oK5/0JAmIDXc1ZSrFBSuFh8sQ9PsTfNuRsQUdvBqHltpgs8oS
OAAaqu6ygo5DOTl78ws4oFi8dMtyItNQtFm0+fTbZuTOgbioCkciNvO0RwXtYrz+
4ATvNZ9zkU7TTF3HRoxiPqijzz8GIjDBCCNPKlbmPXPwWTEqXtK+DqZofFUkfllY
6J7NJpQDR+JoPqlcC5LSQelEVTbdQ6wrUVo4R8pLVs/gxdh4Sk8Ro0N39yYgWYA+
UMuuDsx4BPhtViOkeRlq7wYk09L0eYG1Rgkpl8TGZqGKGGFiWqF+CeUkgsLC09WO
rafCuq9Wm+Tz7pxkx6TDD1O0T5HfT2Y7NNM0IE6lA3d3Ilwq4jQZw69XntbWZK40
SVaSCj4wzngs6thZ6ol6oBv8yaBbd5ra1ve+Ics8zNvY47Wu6THxmXEmRKrGhXEm
9z0P9E8ammBPYOjAley5TR9vwq/ddnSqFhRJe/L8GZ/1tFqz5Yzd+fGYPV6ARl02
YRh1Wf7QXbw7G8zp53YlGCwLtn+bhibztcj/SGhSrfzUaxHlrv2H8PZhZA+ZxqtD
w5jaV/yr+Z3igDOiCd/Y67zIIqpBY6d8ZBz6tLSOAKf4PEOKGunHN60ol2L9aHWQ
IKpe98WIfbmU8J1vNrBtrZaRVMv3U+dQteeoUG9HGLPVUz+QGN82T+Cro/HAAHiV
5G73wVdVGI+L9mTZj3gevIVE6M5ZWLuzVwkjJwgmjOBz/bPGTtBz3zFNbQEDU0iR
VqT6fp6SsnVXnU6U0wI25gbZAxAakUrBRGogmAbDU58CyIF/Z1lMksOTrwohbE9x
Uc7v6j+6R5X7/y1CnmX3m145+6XokRsjZsgHdmXDpzMCE9LcKHlJbpbg8R4bmrfr
2a3uNX9bOomCWcPE0tJJWXqe+qzUVDjVQ8UPgyIzO7g3IZ1eOVCL2FWTWiWdyMnS
skEyeDUQRze1o1FG186tEhqUhN1sSoB1zFWpsIVABFeNMoPE1cDcu6iXwExzcQtD
LTwivLdxODkI1l8h6v51yNv2QHQA2qRvkmsxLryR4Mp5E8TkycYtF3RzkbJvQn3m
s6/niWNLghB0RPhY0JeHJZbsFGfj1nn5Gm24V3b1hslDNyGEGQz68geEtwzS5WNr
DTrmQvZvFX65YrHaOFbg/58AAZJUZMj7DIohEK6Ibqy8TdpNgmtDl3B2XIxTY+oT
ENFLbHCAKihNYd8SN4DNCQnDh1ulNilhyw7yb9XW1mRZzzjUugZ2F+pGlFdy6NZr
n4R2aRLq6eqt9FbgnBQWPC0k7196vGYt5yMBUsYc9PVmTMmur9P7HdaPM08ZJvXV
IyzTC+GwwfObTYLuuhJDp7Y6RXae1G2eaAP0nHWOBO3z9masQHKL+hc99eTe4wR1
YDlDyuE7BYaxnykyja2Cg3fUsEaWo/w7biuVdpSJ9ojBb9qHA2Bp9CtZ2LFagrOW
bp+iqE67NplUbTkItWD97Cx17MmzEXDxFf0eo1FqcUE9OB8oD1m7aRsrLH2KispT
hufM4tuqAj6DD68Ue61vizG0B6qDT/S0ITOSusVaB0LwVvBe/wrX2rmI32Y7sNqG
BsdrIJPMeln7IHZK5AcDbemvAGvZ23K8gpeReI6YMp367TD8pd6pEIPc2LYQ/mUy
vawF8UpcsbKfJpzVKdd5MjKdoSeIpNqe/csEPQMJa2j1he5g9KW7j2gUeJjOOUCG
alyyvHumQ1gn/s5OEsEhZeuYBwRw8Hf3eSpAFv8OvskmOWkWY0GqiLpVD6ou2uuz
/2cSKA3576NMN012iLzcM88r6QYktp9D4uXp0kXI71ZXa48+oPk4zAAztIPCCDRC
4o4b2PHAbPqraU4AZFVswV/LADMTQmU5BF37ISLaBd1yA64SYGxhZh2TzC9RSKoU
M0Td2TNnO/u736gQzVUWLgIzrQ1qW7PA+HVwTh9vPP/RflH9iZNYFAxJelZ1YG0q
b4I5gzOpcjYnSjR1gB41h2O9ccpVAwAQpap378N7xKxA8l/vHS+grL67ihc1lEFm
BOOjkoeoYJrJl9bg5AIwk1BmozPb7MiLAKnW8hUt0CaT4UhH+SNgp+oNvtu+ZZw2
uEyJoAPZa2o71zE5AQ/qdWcszNDDdjzmi9kG2J6kl52lamW+HGEjRnmUjPL0FFJE
gEWJykW5Ho7+XVkTC56q+FVsA4U0MB5MJS4/EZCf4EORFyU9szXYrk61wrDukARg
JuDAq5Q+OmcEl+SK+joBHxXP1krcEsW5y4sS1MKJoijHFRnKtsYEUPIfkRdnz3nn
botMnvBzZ67S4uIAgtWLhDnGUJQoeoJHABTOtvx5VGYwnEWn8P71+jJvHMorWBwO
ImfYe+z/KLaitkTO/HtWBwvW/VRZ48RsPRZQNWmBNF/GmzWA0Y9/vVCsBMV3QqDk
ccjY8h5EKflqfDe7iSghILOynXigHY/xA+pVRWey5H6cXmqz3WoOsZRShST/ITt8
JrEmcx0g3HyN1gPp+Fdg7E2c6qal2Xkh/GBtUAk9cS7Hh3SdyEQB5dMvohV+u4dG
QLMHXHLZnW8taNj3cIHY6x74l2NBnDgw3dmlDNuQ27EjDZ7cyCZNl+VqoAO9mK+p
Azg9j5m2WmbiscU/GFN49yinBgKo++1XfyuO+D9aCZIaOUl7Z1XGJ0K5+PEeyLEn
91twHCCU/cYibjNxE7iW8WmyHRFpc1BxMRKlnomW6ro0bnYkutwcsIAvy3ce7wNF
gZjFp2nJcJBDiKYT7FjLFxo2dyb//ZoohjFUIO6ROc/kzkcMaI8YAl09UYUufPLu
RpNKZ/BF6P0DDQKqEROm2mKVywbzhDtj3832w/QNfDJPa0yFHO6cKO/MsdwNgLo5
07JkTIBE3pXBa5cgN9mqz+JCUmW3p5q13EbZq32ZUXS922xTn5i/w846XULb1rWU
25VYrCRZ4MpmtSxaEdZfra4X1hLwsfIwfI5r2K75DX/oPu6v4rKvIC4Fzmb2RKZ8
rzw/Q3iGBUC6BDz1GfiICuESXNZRznFULiuPfZwttvXFBEMMUBBMjfHHtvp+o/lQ
PLxMbRdwiC/7T59kTSZVaP4Q9F4Ps/O5cp3DyWKbW5vUp+Up0aMpXoxN3eVPfm+g
U6W7jMvfN9lx8X9Lcbq2AFBIcwAWH2B7NzKNfEz3y4/9MKJ25C67w2SSB4tKbhZU
cwGkCB9tbuNzDJYf5pubaACpb23ZbroRnU+FfIMqr2UDiy9h6tgTvqYuIBjckGa2
6izC4MWN39pDfeVeOys0vqpWtnNjI9VKIbwEGzhB1Hqm/axWDZQ7FWOU6D5F1XHF
e2m7NFiLCgf2+vibFX/Wg2EN6nOItVCPWAnJVUD2RaFmNV2HZm5RW3UtsgCL4D0o
fuX20Rczkt4AsqJfdjax7WP3Tjs2QoqMmlwN6JqFGd296dTZ05nCY7xrM3lNwjp8
NvuUIvbfGwzhAKRaV6wurCDj5ya1zOc9rn+8LFG+ZmnDd4ZFA5yKSsZl2j2bx/c+
Ifa9xbs8al8z76M+T0QMe61biVJlUrQeZCRBQYTH16lHrpiwzCTHU6Bl7cxrf/IB
xQBFihaV0JqQi11s6fmnVtwCJgfrNRxMjBzWXUreaD4GLeHcJ/6Gc2l5pS4EVF0v
EbKNJOs3x5KQusyLqm4TdkJFpybKVDJB4ZQ9xC4uC8z2l0lYbgF2lWsILO43I0Of
Hh1/rl/hwf8HYMqixgGb9rOThCAz94JqLAXkRRHDRWQsDmDLztROk80fC3ciG37Q
bcyzOd1Ivr2mWOO2W2eOZXeLVi1X1a7X+bjyc1bd33B7O3MsJoa8CGi7z2QRo2S5
LFUQfplpxPYehL5pvAfAl8jft7/c8o6RsM2z/kf/SnWqvrqlZH3TNRYE1GNXLqCe
zeHEkHQkBHXsDR1whqc6v+8AOPPmyP2KMOnLhyIkg87KRrchXs7nLD9Wfybbxl5X
6XDF6Ghw9S/nv2wF+DBPpWYi/gHmCG6Ix0HsTYZN4vXTSPuVq4kmz2HOvLMBILFN
drArD7Ea9WcGzTjPupAeNYgyOcLMWEc+0DE/A7NJxYaeb2DJGjHa1NufYQQgFcnI
mWMje/OvX6lac5XSC+5aPe+Ym2FSj9J2KIaekTywUFyzMELC2Gwvr0O8RGWj2R7t
XM/EJuSDgg58A3QWsd2r0f3d2YY4+t25ji2651jfpXUYzubge23zlCXPqltuPdmw
D6tWkFX/BOn1HA3Cs6FrKNIXZql+M0XzdkPr9wIGy1/N1h3bMo2sFyiPcGPLxq5l
lA3tobqnihahxYGP2mWOhoOgtVDKeUMBrM8Ka1M8EJp0iDv9HltBgsppaIwpNYeq
ojrVzc+RwiPjD4CC1wpHrt1naYbmjAIAKTseXcHUv56NElZ7fBnwFiBW7cm92/N4
GsRVn49bApCgFA/+P1tuJsJo084kAj49pidvZ0rb2VRBVqH7tMI/Yq/Eb7iJIZZ7
AJKWjhdKdegA9GolY9F3hIyYuPYukoAMPVSOko38F/z80TmZvCM1EJ1lymRlCSp3
xEdFeO8QMoDjWa6BoRuQ+d5m+9kwRUjVtZypjiSODpWYypCQCFLtqtk/ELZm8J2E
ar6DpAhttlLWFEJWnB8N97HsBlZucrJm0leO/k21cevH/DlBtfLfKEyi5xVs0UBt
KPEan/NGhiXdZCpMVXgR15iBNlPRGa7rIGlnJefny/vcNV4SE6O0DUoBYs8KYmio
/mq2k4zxBT3XIX5Y0udqZz5BjeNbp2wiPNyOnGAWQtYjLKBRRpCkeGUJSFUnu1vi
4MpGrEZvPyRAvJZfzWB9pvQEFDfVIVBmDlQLf9vcNsolQ2FO/KhmFsxeiSwJyA6+
EANulJsoVvFdQUrlC+XtBSaRbyGCl4pNzo9SA4/SFJ8+7MDucxHlDl5hW6sd8D1t
sQ4S4jW7jg/EEIo8FWdwd08NuQMiICJ1/nahQQm87h0DLXZkYL2knmqtpuH4OoLP
3fw9p2wNEaAOj8+L5LO5z9mi05jYooz7AW2Owob+NlHs3R2dlfW0fkdtUwnRYWih
Sq24KKnG1eR8DZS4Jw9J+b3Ew6kvKtZd/R0e79CRS0KlZQJ6+OxRFwL3liWvfhGr
DOMZO7nRXtCzr2WlH9r7tqRLFHTr/OJlFAWsn0EBA4gJwv1vYqj8GknEnmA8lhgk
yzUWZW/6NOl5jTrKB9hXNOFaywJbWG7uLN5skrZewotQ6ZoJCNHEZFTupaKxO3kY
RuSbdq8XaOWNMy1FEDuOKaImxjfMsM1HgUmO5dLM8dVhoT0UaNgO58hpGSLXTIZw
rWOSitbdZK7axS0H33McUZ0kXBV0Rg2cb0GjAIaWv2IWtfWTyNFBe+tdqV20q5/G
6x8lwCrMYn5/gowpBdkZ2Do1LHyENrJ+3y5ebkDUkWCr5TGQtQoNUCPgVk+kYy8n
sG566vsPRZxtID4keAdn0ndWHmiwvw/Om+U30L+LVEO8dssDEBSfv7QEXodSpmhD
gRcI9h0Uo5HA1fCRKZySuSTbuGIfOu6Zr745K+19YUMOHrk8ziq9jR6+S9X8pi8U
8XRe4r8BHd88kKdf2mtWbjopMaqglgmg5CRotxtMk6jMbNkSyJVU4DKivlG3O0E8
mmL8RNBMq2cMtfhqivri783eH99EhpVmxUY8c3cYY3IkCEv91rQWJ0R7tXl3v8Bt
4hMl5/S0TmvRYYQO+FvBRloX1U1MuV+uylKbbzuCOomXnGv6GLhTqkpknLb43gUR
CA/EgbxnY4JD6AyWptoE1HAvysm1KHqDioJ9lvIapqyWOK4rZQGcwK1SqnA5M/kM
CQtnLRpujjQU5S4OMOx6e4MegSK+rxgkrTT9B5D4N7C9YAx8e/XE2rgneqUZboWf
56Gm011LhfwQ7Zd5yX1O6jvg0kWlXHI/KkSYHLSj6EcTA0wRO3wRpmnrCm+odWxn
i0fICLrfD0yi33xMDN+XrutfcIOMlCyCbqgN8QZby/8bYu8y3+FPdQdU9LnUsgpO
hU5qaM4JCpm+nO9sd2j+kd0GEGkTa0K6B4IATMUUdtlr/WNOlqhxjqlpQzavtWSa
aFUGu0uTKzYVBcTcCHxGd966R4VZ1oObTMAEURAY8KiKcy7zIE1PVaC/FEhoz5FN
jnAmL2Qob7znrHuG/spr4U55MoNw/W78O29jetlGZgRFEZrG1DMRc+bzhWCxkMeD
t5NWWGNWGageDoKdES7QFLKaUaPS6gaIAzSodzs4f/TRuDOsxzVcK1L+qlJ0sn5+
qVsT2Yct8m4dDgIs3Al84JrpaRHxPjV+7RIOAY6XWNy7YGP7a09l2JJYFjHJlM04
sxipTG2IstdBans1aaSLD5lUFoScQSvyIseqcQUgrCPzNViazgNoamKuLnkHKy/k
i5gbUuEILktd4x+lmamPjRMf5XVdI4KYkrIK1cgoGteApeUcPebGRshfNeWpAGGE
IFmPdOwVGBqIeCFxIONQKOLcukZdISUyzbxziow700u5Oo0y76+COD/25+LUCmqg
amDN89mbCTchRpMmxHZjlns+YZ7GVdMjvdgA/udhYdgiZq/iOnl6wS9wCHDtQlNU
gWGaIgUlK/xANWy+nXqtyxuj/T/AVJp50fv8m13GjFYlMnyfYXoLwPIiHubW9vKD
oeMfY5+6Qs932f0SK2inOm35/qWNdbkSOuorDonj5adUJjDN1/aUZ0aPFYk5RYFK
nIuGgptW1rAPJKRAIsXssdnr6dJqnbONPQUcjyUkVhNgdyLCY/U91ZONYY0E3W7S
GldLKr8nMOD8KHLFG4HlwoAevfA/BBBTnUcCGepQh5M6iVsrMQfWb3FWdS2bSFlP
ryl9r2V+9fbpDnSLsJ7AL5ee0iOjvgN8UHXY3NHKnYih35nTJRr9+Ry9v4sXe4EM
M53QuGpLpztHtLHGYw4TWfDtHfwfSyKpnp89eL7LwuALy2qwZ/eG3c0rtzJ05h3K
9mEyKMbgjiM5iNpnN0GBHkWLm4qEJaW3fVKtDhq9k/A1LXnOlp1k7rsCpJMA1FGR
42PN+5+ydKQ6qsT+dPleA9UNQHV6dAzR79fKsrNjvEULE6PCRnS5AkgT1t1qOK9z
noSh61YBkxvbbG+ou6SQkACi+/zN81a86UPlkipFnhaYVxRKFry1oDFlE0sfZKpc
mYLA0voN8kCSTzTzz2xjtMdMOOE9dAGT3WblnxD4se2ioFCt5f9cKusKYXFtW4ln
g7corN6jWThTa0BRRbbKGEX1CNoB/ercTdn1Ze77yYhiXj7QG9IDcxVqinGsRlEW
BG4FGKQYzqjI/G/nq9l1811dtk5yXKpJOmjLk2yPmN5/4DFeVP3lcEATyjS6iDNx
9zeeVom7d6w17AS6TH8Prtl986rXVFF+23hXMullp5NBlYxzXpGyijPsbPkebEc0
zuBjg1mu2VchqUqB6XG+Iwiqey8fsoWmnqE3XwQuX8FeF5nmD16bxfp74/ybqr7w
uf/GUjCYWw1QXASH/YMZqVH5hao5NWYHCWGqhko/M7T8dbISxm0glKUXNBmL3ead
5N9U36LNdQF96L36AuoPyYZIkn1ovbHuDnJQBkTL3B9nyViSJmorUNvcoEI39H5d
zxBTf08U4D14McTs/uKiwHsyKuakewwLw9za8/QxG7TainEQcTSqAmQ4p9RwPejI
T1nVc0lsoxFtS9QWmhCUsxQwufafta5Ymj1S1ari9L+ZolKXQanl2EqypkxetaGc
auhLStxiMUctr7f09CvXO5bmLnioVw30qCfiofm8pmY/SpvA8Px8V5aZtfqZa8QB
KYao+cpjyl0PbQRk+5bmSXi2+IvYnl0XCfvCgZ+1PlzyHHT3zvVuX+UMzKtpxYAJ
USowCDKuYRoEzzRdukQ/jWHWNIDrFWUo9JLc3/0wRmiYOG/Pz61cTAJcQiA/uDiv
TNuQDITLbWwoeX3DHuaugZIj635uiDsNTSALWCyzZAPnfw2p45gyBjDUMVpEEnno
0qEmIJAzeDMYV4fOJQy90udgjv83vXhEtmjBdOgsFT85dUm5phIB2jMLD/GtIU06
hzHjyajvKmQELFG5UN5qUpR1KGRM5ARkT/kFVYHEvDt2tBt8k5UTtQ40Ibu1WHOQ
ebxIIT1zanTG7kEQ2l3nWXdQZg2ESslsXz88vPvTb8G/mBkbveTpL0nW/32IPm1i
iHcJuPP1Y0b3/WjaasoUwhXETfcpi6itoJ4a691sk7vwuKFdgVylRQhafGprmgpK
gPeR3H4qThsQhb1HAzqFbxHWAfe+JlXrUsIpILwNwqcNMEMKX8vx5EcV6UA9ojNc
ycoYRrnkhh7TMbSdod1GMihjybiu2yRfHr9UhtsKCJgpdV0P7bpOlxugSFYEhEGk
A64UXpRAumxwDlvbLsJh7jNxaSMc2gdiW4aqDEPipJvaIuvxuSqBX2YD9dtdMGKd
9u7vmq3+0QzverlcJL8VrBX4FucZHfrnqoJ8AA3s0CeikpMPrTImQQQk+2lKO/RB
JHtO+DgEkfuNOzsIGS+pBq8d2FtULJSMHnja3NbgwUw8JryxuybKVjEHAAWE3R+U
sENmGrW27Js4tulJEK35ZtWlUmw93kJ136bsVx0x/s0l4kUcuNyAmxp0VocbBpmi
JTTYAjJehf2O90rMCFwNX4SDBXD11ehgjBGvjSAgUy2vGAKTH7b7JgE98U3iOEst
JOJl+hoq9VJrowAV0FtVK74UaFHtiYsqLYMFqr2jwWPBH5v3ztb95AATHay+uAzy
4CZbhcQwIHyU1z46BzMjoYRnP79GajxjNxfvqg3Xw9Pr+cgGEjgUNyTpT6nuXJlK
1wslTeIIljixJ7+eQndPSVWMKvF7AzDWBW+lBFSjd/r1zCvqyGTdf6QrmNzE0rPc
koiFoPdQBkyg8GWr1U149hfC/z6KlWiEjZKDAU2HwYufkRgEVmwQQgYgiHWPgXid
MAbf5z30KrpCLznb3zld/uhM9eZDjFrV4PkcqgFB5s4Fxh5zd903jqOlU/qEm7kV
HCPyNpd09x4RQFhb6HO63VIQWrBZAk5B83MW2orRx+FN9A7tGobGVLLUUYYep6ih
IaDquqjwd/TlW3wEyDDRenyXbKz78DIFCrSpVIY3+a3um/BNgcYTgTIhNoo12scU
TNpO6X/kFej+YTS/HUWk52xjtrrEIOJLHEuB5u22J5sxCTO0RfcWxvxMv9a/iqFx
1ihLMgve/1rpja4+Yu429gnRdBw7kbnMEhkTFAbmRv+SJHoVdSGfbP5BQvuLLmOZ
WHakvgSHX7cu/dSXYQdOcormtRbBxdF3Ly/QZVcmI2dSLdZyOOorHHKj+OPkutW/
2KxK46fEEotdGXU8DPNuuTjiT/wk0jhtM6j2ciiTbAjzsfjKIyg1iz/sPa/YnOsQ
NrGNiNvwbcLngZkJU0vqridLi4/GegFo7aDStsdtkaNzpt4tnwev33oGGjBDRlGs
9v9ijK4TxOxZ33Zhv6TIfHJUzGq7xEy+ugcCgAnHZ5nPt7aA0BmXkDgxee7Tvrii
K707w6I/5TRbdRXJdYyCUcTdRfC++v6Ot3nA5LEjeAe04YQsJ7Ns9/GK1jaAbZsL
dgsZVuxvxp7rwYKN6aHltzViuykH/f5j4/tE6qVmYDG6B3x6hGjiZSJuEM0CgWH3
xmWD10qVIthh5w8Z8q5nd6HFkDG+ZV9Qqb5OxuGqZNpaESoihmsauD66GPS88txg
jbugf+h4d2PIkQ1Ro4iiFPezlR9yVwkyDdE1nWrcOLdKAWIcO4SogMSog47qjw6y
yE9tj+dyhMwBLZOhn1Ld2pW7w6jgOkbx3EArCZR6RiaP33xzP9DRFJRGBkXxpkJ6
MfuD+TA8ijQ2m5WGkqKN6OuuslLxbWsZzr8OkMj/RQ4h+rWkTjG3GzfztyF3i6Yw
i4cnK3dDkqgnAmQCgnW1U4ubnXXFglVf50wmqMjTJmyeK6qOjQwAKJcLCzwexRxb
203TaWUHV4lsPox4+x5AQhRY389n+9vCCo11Fuop6YhYTi8Rg2CPIHT0yYc3w8qd
EwhiX5VIQwym6UTxiccVmKNDS+T8PQDYnX6R+utocyk2GBZMkrJjwlVSpUAXvx02
PVAIrOdamXt8TAjnRblSjzQNkPaEFiFRDrA2uMkks9eyJwCpREl8j6lg4KKf2Siq
gf5jIzjCOZ9IoG0zbUvVaesnh0h4T4h0ouOu58jbOwpIDAiPGpMpbD/csFcfRCkw
lZb9BZ0DAqISLl3LyOKryy81RxcKzhdkJM3i7z0StvIwTwiFoFI9KbwQ5Reu4HjI
87+7T+8z/8ge8/PFLPajdvRUvw8c6UMWX1eUDeAvELkCT0MifvvrlF3YArjTWQd9
LNufUEhAoSxLFtStG4E4hlDYEmCAanZDycTMIAD0j+LOUkzNzU3bfwJijPkWZoGH
NEj67JJETyeQrhuujVIkHK+8ttUUKLlyVeaG5bP3r5bMkZ6MUpdSGYwPPrCQMwp+
zD/1O7/QvKQ6nwwnj4wy2aqPQ07a7F+70+BmDMvq6arRtRpL1G1BFsoHDQPar6Sc
QxKQIUYKwAivtKygrrQ96QB6Uwh6a3BbRw70WjdAqpUBoiZKaN9GlNaGrxRawSTn
fE0R/fHYYdvS7mTyByTgHf8T2TbBPNnQaixnCRv9gVQVCVFNYvzIw5nYjdvdJ3HX
uoNW+loBiqoBDzNV3/wutCj4nIDddc7tHqPJ+OEtKlhK0Y8pxUT0TV3E2OgzBwZG
YU3HHb1xPtbkALihmOLuPPOk3YMbyJq0lfy5On7FSHGtnkad4pqU9FQd9HaO0iF9
9LJGt7aMFaUyQXYPEqEU9PtsI8I+1MOE1w2yj7uAWAHFZMfIrt2Xcbo5m5xhR+1j
lo7aAy1Q6EugjXCrzPcpfg9ITdmrWxDU11HjSI0kkvHh0OBhhLlGkzxwe819yQeX
4SwP1hWnnoMcxFSssUwDQxBJ1y70s9CAY6O53zA8brGCcy+74bdM9K7f7hD0QDbs
zEnzs+w7DJfSjnFhFyQy2XzoVkqtk23qVmXlSCCEqYbvti3/b49I1Dk3gYy0vvtG
rNEo7XVmMkzmAvzz8u4ided7LflWHZgyrnKLgQQJVKEXP2T0MPHGFd0grg+Op/++
6Dhe0KUhUkYT3/vtf41VbEp/gpeDdcMi5/ESdUM6Qz2SuNoM58+gILePgVLY0M5t
BY5+0aTbCObXwAWzMxSxvFN0HZwKMLO75rdwKWq9MNxa2LNy2t4OR+b2XKugTNUu
Xyi6U5HmQW6ymrZj5ij+E8POKK1mMJ1pre0Ww3oEMNALfvmKcH0Z3XdYflegGwL8
qYAWKt/MoPSxCROr/vwM6lb29FZIj97+tvc6dnvChXmcbj2I3gSuDa+64RCwF1LY
chmmXUYbCL4kET0/kbrVAO3QkydlXXZFzr2j/EmFBi+7rW9t2YAUETQ/szv4Vv9f
G7NBgDR1kv369OhbU6+XyiIGPFCyoiJbkhbpeli89ovl4FKOFdcKVwWy1FJ1hi3K
J3hoe5A6E+yCRPMF3zKYLXvqg3NudzGFsm6YJffgly2yUYni84QOwrxvZCbl98Wj
W5uc+z69cLeZVnQDiipPXw/hwBS8zkH27/jHKRzaKBe8rGplh3/h0ZtFXVWvpKRQ
3FdabNZu8VIuVhJK+rtE+U2tCQz3FgvTLnOKZmsSm5VTdhZTDnkV48QvCs/e5zS5
ze/M6qf2ty9f1lHGss3b/03vBUwW4Rtkab4gT74QT0+kPs0NH/POgRzUaNhcEaqO
JT8qx7TjPKPfeNHGRIRZ33NTRJHPXdvUSRGLwrPgcAd3D56McC6JQ1XZ3XdPW8eK
bP/yymq9PFucXRFbLqbt7v3ws0Tn3WrLNI27dkxtzhCGejbBIEN0ny+4unWDZXHs
6uPh2i22INYwFqywQrAt5ggwXdIuOdwpK46RP0G9VJHVaZ4GTGKhK9Dqotn4jARE
FhsF9wLWK7oqZp39c/aeVgJL60YIYRTmLYfmZsQDrEhWCtK+3N4SLhuplknNvyNa
3DKZSsrGv97eNlRL3C84gATpw2ehyPE5+4jURXUvNDzEDyrQOpsrMal5vKwMs336
GmaUKPmVVsfyvzxYvmfBKeeSds8EKXyizJhgMAIAll+krowRRcm/e6ZAZewV9N11
7/8MQgXjwhczgxVCIHWBwr759oe6FDu2n5x/R5rmqTdTqgOhmIRRyrZLThXo9Gnq
torYlTWPLhOyNIFCxgV8HckeRztwDvyfp91s4UjuQCG1WSc5VfVowW7vVwPnAQI+
gprQUqHWf3oSCMao4zajOexT9/5ispMfj5H3eoOgU/j7ohBvuCNbb0a+UieHwATq
cC2wW9k2VVYzcNTupdUx+VvtU5cztrqA5HWirbbXm1lnnWhoX129XBeW+bUQwFux
Bk30YsEYVUhqW5WY/bpKwxpT5HLsm12NHksyKMjQ0TnEK8uR4u58dK8b/Cbn7xgf
hK/oeJzSh5ztt/U3VpWkXYJCV2O81nLFqBW7bRNJOgw66ulLfi3aAk3mkgpBRmSq
kAqpm3A3ymlfd+pNCz2bUrBm53f1+B3vWLhp9xjuQE+SAzacT1vSwqIaMqlgFYHZ
aMMCzcY1O3w4RnDHZUAH2fagKeHjV2FaWh1yeifFkZZOAJSWJ5qrIAh/XKDcQMXt
Vy0xDbBjocqRCm09xg3aSPIgbk66ZWbKhNsg8UcNMTwm1ubKFcWCCEEOJOURQSib
ttEnVFTMYaV8qNByPA2XnU8Me0pilkMUnCnalglacGKDkTkQctQcGt5+ZOSDxs09
7QpZbOmbnLsqcY7TNxe0xDALKwPN7xp0UIcJV0M3aum34EQCS5uvmLMv6zSPWD4Y
2Hx8+BhkSJH+eXZyNW4NSyPUrl4y8xO862gNO5q7t0A/3ECpLkuXSNiLFeJQ3ApY
tX/WeZ8J7K8w6vlNDkgKIxoLzdfL8xCeJPVb6KTZ/VYZVPGR/GDgbKkhYT0ELCpe
ym/ieUH+sPNdJhqBVBktGguDBPKOkCzIpbxBFtoV/TAzYxS67oFbSAUVWbmtx9OM
TRPkZvKGCGt/eDqb2ASyr6+Cx8CtY4sAjFep2sHbodhmcIA9ve5VXx+0MT4nw6nT
/fDTlyOBrsyT95+RqFJIEWynEN6wbj2zQwPH4BDMz355/PTQBFyFLc44aGgCGUKm
e0f8BsNJlyyCrs9gm4ipaIiXQulnxEy5D9qo5gtPZ47rpkAI296f7Cj53Dz5Wskp
VU9P+OxJyLrh43yV4d3E2VCr/JsU7CLLlwiKisHLL9n98YJk5KOh5jFQcw6VtFDO
q/cXFIrET35w2wlsDkVa5Q7xLbm1ZACI9WhF0PotKzQr+gvWqBU0VvwkUoa9d1gG
2CSylo1KA0HTI47NR8nnRDpN8/dBB+v/9SL2JhpQGSQiIClXoMuJ/OlCwb21hfwa
qIPLxnbDPjrWJtlNTbwtGsNt/N26fAFTgOd6bMGfu2lIQlGRYriwpU4GWdA0ZaYd
osPpV2MDH7Lf6dLr653tK3+XYqLX300B8gbuD/vJ+dsP67LH3ZG1lD1lcoLw6nWB
NQWm8CAq3p+Vfj5sxa1mI1k3EapNoIGLkWg0doVP/snha02/VKtQFkuMdIXO9Kyd
4py0mY/Re3RkZmKVOFJmjTrA/XUmZfGAXPlkhawcFKwnROaQUxuv5eZflSXqCZRr
5sfBjoKt89N3jjKxNlJzo6xwJUhKUJ1oYrLEpQ0Yv9uIwWqwbGFcRFi8eI6QXMc5
5dhfhdO1PuDhbe2hKYbqpPjFmNdEb3BTq9ImHod/ipfXkC4I02ONSLE7AA8bFSH4
1e6gZG9Zu+UiSV++i/AD1x36iR0pbWcChCiaS7LykssGhL9VMI6AyLTfynx7FQtM
cWRnuHMf91StGrWnzXG4W+oX60D2mfCTIgvkQDQbSt+NPCBvtxW4cdCQ4KJwChzF
cK5/na8sb+KdMVNcA/TMME5IFksoupHKikKFPIme6TODtT/xP+oqzIaRVtXmMx7U
lruDj4v31GJfA5T20efqkY1i1bkHOMTtg7D05Hzkn1KrcO9wk01Q6nt4yHeoVKj9
C1yjAqPsWdJwfCt+TmVgKs7ax1nv9TV+WipRkxty1tjFBBL2mhBWTYFAfMTbhNZS
XeF28ngmA5dCu8eNnbeZRwUBryTy+wIQ2jnJQUHogl4aJ7GBmT4rnpfUfgxx/gCf
2tFJVktCPnf7enSRbIaV4E59r/kM1hV733QBpT1KGasP3s+Mrda/Og0iqPXRJ+0U
+HdF99jRnAnrNCv1JEVh/gjhWeZMhJQo4nWGbthwcTHOJf0qGMDpx5ewAM8b5UCu
MpvPuWTxrzb7SJdbrUl4kG2E9je51MpioIP7W6K0Q/ixmGAyAxfL+JSyA+8qkz5J
dCXaQoilBrnAcoTMfurO+ua95a94Lrbxh5kdrSGaZ2alB2L8CzZAP7ZrP5aJbRmo
5dtlyBG40+dPqaAX51+oTqqESE0xlrtQ/3riclXA91AIKvG1rj+GVgK3bN6JogY0
0kggvKPLhS6nOKdrZ1XkRIUTRrQllmOlyNASB3uMNDrizPLqu7IhV/S+M1ZRU96D
62IEI6rvqePvJ9GqjrAE4A4F74aBs42OTeYq/W49rH/I1MpPEXvXOokr1VeyXawu
iet/6Zg3k+ZNtxFhxliaOa7j+tVaarzDSw/gkr/IKo+ufBwZK2gRg283Efsmg5qK
+pPF8F0Y+C0SYh0fCXi79oU0yuXDk9aVyaxECbba88BUY8d44Gx4hUZZD1aii/AA
p14Y2vuHoxAqfPw0RqdATvAuhYsp4sHBsZl4xccPn8fA2g9hZLb40EmIZkOdQmRr
vuoI4UizFqhTktLhuMVKs6k8fZ9kL7ayooCgHXj985Icenh69wbbyQjBu88uDHVJ
w8/ZZdlpNT3Y74S2NFlfUnuMXX14Z57JJia9ZQKT8QXWWQb7KotXIopgmytsPPb7
L227rm+P8ueOZuuSfkeaoPrbS3SPtJymASh0UYarlTkQSYs562DLbwHq+BZfvfG3
vRSFakx04C0YrXUmIH5LJRPyfNzRA9r5aTbRcNYAvV/v9xPN3XZattJ6eK4a7s5m
tdmsSMarRKZKYmnU60wCIdQPmylpq4qlGiSbpG7XWDUd2fBSYxTRVfmBNViek2xm
zSM0eHhyQSeapnJjkPN9+IQqalACo+g25hg6UX5dcC/iZqykSmKY4wYyLCRZp7OX
6X3a5OiItUn6ixRR796kbLCtDBG69VditMRDHVbLxoZsKJHAV2B6IqDvIlhlwKHU
u7e6z3ZNaNC0WqUNo8nDiTUys8ueva8IadqYbwtrFymcl+ZDnmS6w8wltUGwvHpw
ykjoq7uT65064cTUZAcL8ZelirQfFpf7i9zKrKW2rYlA5qaaNaKd49XzvUffwmMK
j8QoBkMERs1SG4h6e65YGcNSD05keU0gQYYNyQbIhlVddltFJVMoslUvD3lvRjWX
82JKus66OegqsLeroKwe2K3RmPJIZ5QbN0OTBAkGoM/6lKQ4KYF61oac4Omk5Foz
TtLpB9A+XXSuhLEu5u8eUS86SuR+l3v9NiC0qiUEb2Kzp4tSTiGkgblL1nUUWSN7
eixQeNj+4rOfVHEpVdD2Gh89DrAQSBiFp0V9P8TswIAyVi7QD2iwfqhVrOTfY1qr
lna+pAJqm+NLL67tykcZfw3UZSSiaowZ9MlXpyclJsCCDJFuXAv/48KG0d5Bt4d7
h8dr3WkTHD4ogEIJ2fLa915Lev2R8UVcBcbQ2IwD1O5GX3ahaKX3dTLIsLbiPe1P
lsjZAgyxszTNnAEF+pZ912ykow1SnvMiB8W9sWLct76ZDOT7abJBWLRhhww41/1m
FQ30gZlpDIN5Z92T7J65i8ouzg7490IZrSOXpeKQ5LQH+jXfFZzBSNkWeKA/V03B
4VAFQTDmEqW1gc4HGjocYq/MRTixsaDP1mtCmEj8FUs5iaCQkP4B2k8kZABpLzoN
OIAvDI0nmzwAaTo0Yb5dxp/GxozOaJ32BVNFIXts7DQL82FmHiAm/rPkcQLQvOJd
yYywdW0gn33N/S2Sf2fRCZMF3YmGINJ4DwErXTxX5WPl16irEPZx+uGdQQ1imjeN
GX4BLyu9Xu0usfY3RomP/O+LcCdqtWfi8iScGb9ZIzIRSN3LovagFLIQnoVhIbf0
XdWubivTs+CnyEALVFh9o3wbq/CvCSb16G6+aKw0K+n0lG+04TIv+gZkjyXc2uyr
FyQ2KZM+OTQ/y29hHqesCPqsG1KKlnQrWh42HCjcVxOFZKSRvARMYhtTF1Ys+Yah
0SDyFxCXOOPbxRwjpXRrTPQcn3bqwU6DxT+ZMkclqiWWQv2cYqk3+pAD7tUmhJwl
ORYZtim1gr+0mPEkzqBu3qkxHPzq70jZrCxsxtUHqpHgtQCAaS0X482ZsBO9NlM2
r9kD3lRXKczG16ukQahpqabbAXpTYhdWJjWkcqCXo+UVfFa9J6QH7S0hldIdv9tu
dN7UO87RAgb8zzLzavIeiVOQ982XPepSGfgh4sJerafWZCIKVRZjHdCeogTHbsN0
i3NDJrbkKkKopS4zKyiarYqAtSWILFOM2/DpaKRPTU9Wjy55jqgko0VzlVFzg6oK
uEUgjZWY5a45fK9UTeFYIArcJ6pevCvaSxuLRu70v0LEVtrG9OSI9iCQ1QXVRl9a
/iWTQ5QFIqDGo9KT1SzVKOLlCKNj7PWy8LCBl4cJirA6epr5PHxhIMJH0GM9+ajb
ZonZhTasjCPmzpUvLLFseR2PvDeXtqdVvlj8P8JMpokxUuBT2nZoWn0AwkdXMmw8
j3sgTrc6nrziDYS/85gcIvk+Kt7TovyFnEsJgugW4+z2K8r5BVU9i4C9E+ZyXrou
/KRRqGhN2m5VR3cz0SmFTAJ1wd+kj7ss65kqmVtkGq99gVWNyrM10muv1AQXSdKB
7LIl6QMkjkLDFX0oQvhCX6btHlRN1I4i6DiivIO7VR8RDVhY2kr7G7Wf8jnfAn4K
rDQUWkeWXDdl56JrGMhkNmWYAA5PVhnEQcue1rHtWm8neXq1weHvlIz+ca/7QGk2
cgorUcKb472R0BcuN69kBpJKyHDqO7otKmVHiBE4zDK+FBry19rxNZHryMg+S6U5
htuVvWZz3HKqsRjJl6wJcl2rkeU5btjLqpY1LQZgqIn/rhHn+lOq3QODOLvERVO3
C4vgO5MPJlowfCrNsSbsufhTwxIN6ewJiSAqZkYyjAhnS//1ECTiGtA9UHGozjBv
2ynx8uaRCsX+hHO5GikxpHA2iyISqt5f3bq4WZ+fRIg9MVr34kUf24roohWXWblD
wDDMbOtaBOo7usOA5a+jt3iSmnurht8lAwnHGLHPT7HNHSNn47WGvSk2kPSLpkfr
dVKKSQTVQA2/H8Hj1tOziOzfBr0t4a3v/s6qwDoVAiLaw4wOQtZB6+RW9ySyfOEA
9FG7Bu7ohaW2+ak75gP+lKGqYD07Wq6Qt+jCEj/iTLbXb4xfabYB7S4wx4YyIcgn
iTTlT5iezUDpwZJ1SwXCk98V50pfYKIEjDowBqBtmtkz8zd7if5EnPbbSdQoRIMx
n4supGpuS4DHqXhSbo/CLGvvWzujhSwoRfNTKFTyKux2HOmYK7DQJnzncAiCq1Gm
aI6dH+iYul0CvC/H0KdTTk2NDZHQSVLGu74IKS9ANC22FRpcA86HbLTto8dmsMER
KFBKzQeO9ctlYXwSH3bqpOH8qOPcqc7Nj2XBM3TVBj4IifH/dmNF5x9GDJADQCWk
TQMOr2PHEmP/Bu+g+i5xKxAfVPyEMq3JD01Tz69ON5VdnRSVOTYeRhrFR6cCi0Oj
T0Wv64JneRjs8iLJR9MmEneLHfy/OB5uShB7nnRNHxaBQDALp/yFZFBo6WiasAti
iHX0GQAZR0wM5uW5HzzutgFiakkgD9dYw+x0aSskwe+RqfA8j9TJtRlUeH4vzcDk
FMUXW/FD5gdapcHLutllUFJgcO1Mc95n9CnlF/Of0yxmcEEqAp2i+mONPETSnHuc
haqKXtiyy2xalFlf94bWk+e0D8zP3u2qzDqwVYqTyQ1Y5F4D6b68x0fJL1uQMv3t
jNda4JJTKHFgcJLMpUm8OywlXwbyyCcpu8OjTDE1erFbYg2mz4XQBx7TfplPk5r5
0hnyLt/NM2qIK3xKLryPjxKqAe3y5fFW0guLWNpfhuWItvGDb/xvilqswqe02JnI
rljWSO1B5kn7gArbZZD7XB/CbSvTXUn0iUBwdOhw+GkUJeRr2reJ7zmGGfBZScZR
Hin+k1at5o2ngB7BBIim+eLISF8Onbh6lob3WI2hCFHetV9xHAZoukRFoA70pWmr
1CrKSJOopxJr+Fh0RjbE5GbShA6Kqb+peS8yEcHVsx8bfEnPDz3SadML1iUNiY5T
PWjXmsFZ0LX2lcQJzg7+htXawyMhytm9n+zradQVQ7dxXGczX33vy4s1tkUwyPQw
aThem4XPGREbQmQUN9ocGHm1h4R2pRDCbRJhxbvzI6IQuxVM2yWsNIb0cn3tNbXt
iaTnGWV2o9U7SS4wVIDVLK2Udzg85pdLW2me31YArCsbWhJ/VX91i5fvP4Kl20N0
uKEp3EdFCpFPJJzGXxHGcnnOeihyhZBZBPfqsWprH9HkBaEurq5JNQfzyPiMvoo2
GS4QIrKnJmpVePGvStHsqrEUXydR9pLR1+/I1jryA+IOIOIyk3KxdFBm3wTP0Cbz
6JDRifQdBMauJhgw/1N2Gx/vTqMg6TmrLRb/RvlSOngky2BusnzceJvJXmWUxEHU
54nDVluxmC+x6YESf4ZXBOBfkex0N3shdTvuTCBmPvb98cvZNlKh0XPjrKphqruz
1j4Cl06CdZsDthJ0pcrL6uH+DCvk3jq2rqJxcne6T32OhOfV6Meda8usjGi1Pbxd
ia2HAPMVyNHNxiJY7oy39aWJEYPxEQM1AcAzmPyv4zwBtF6Yb7C4ETT2y5qAgH2P
njPTipthp+S3wrg2+zbIOBJDPaoTyI6t4evBj4+aTpi3GamGS+QuMF1TiefPQear
wDydcBENehlzrKaDgN/hX/k13lljG+9jLrksweT78wvPaOl4ETpq6K1I8t8JmwAn
DwdpOt5dJ3AOTywaz+BqrgW25BxDXRe7J53oK5EA2jPw/rzigmh2DMwZvVL6Qoej
fxPrvg62NQUxcD5mY9jfxY/Pl6iRfpFzXgcuY79dMBgnxDwJKuyKQGmhPQu4QCZE
fLm3gV2Gy/cBqTNq8O79JBK2DDeNsB+o7lemLMZpB+ydvpCjSAOzwGVcpevXgA3C
LEPlhU5rJx8XV6qbNJFOuv4LEEj5s2c/6Rl3+ymsXDHNdvb2isZEDnBemAS0Bz5y
PqPYA0ICq2dWc4i2+xHs4DBukevKk60CIel6ONqQMpBG0DPOHmd2LjISrY2BL3bF
KTFqoVGYcpwE0iRR9W4m1e2l5WhGmG3IMNMg+6ZCBsNg0EW37zJiJHzpGPKFQWZe
TxgTestva+e1Z8siG7SUxYnOzMYspDQ6w6Ier+CS8ntNfxSAlz8HzIpmIm3fFkUv
0GP3xRBgDsGX1SiCybsKEMkOrmb5o9gchTcVJWsMijO4/3uTM50x2qaMNMCGhdrm
6RskVcH12fFh1oG5AWhvWutG5bX6Y2beaMTVpKyKCUlG84VBPxuGtaFsoRuRu75T
XmTJOfDxcjuRQymt5WsBS1cKYahnQpjq14cyIYaR7QywqIaWSb2PJ/Yc/CNzP9Gv
WPeyaRvy2YKeSxySTTltjQIYgLp0CCtJl1iz8CdBrrQAg1+81rGSPjGGEEKw8EqU
x5HNhFwBcoAb2HrnltQ9Up6mXddHPY+/h6FMANVVqIswHgUsbcm+lOXaN4gFghdj
ERzVooqQ6N5ht5UI7rNEH7h6LFpJ6sLynhz7jXkcQXdNoR3HyuueRXPp0OeGV2q+
CzoSJAFqA8MrgeElBmFGtkTKBBmVMXYIa4PchpvReqGwzZGZZsZTFfySx+IHCo+K
X+RsLk/z6iXOvoXrIXlX4ZywXp8q4Cpkqw/9qxGzG3/qtBTc/P3eU9sVwNvMuj2a
qU8U2i+4T1RFCgY5/8amtrHkBciSDOJ7VadYBBnGEVBkZsa3qqfMVoe1Sx+UGZ8p
an7sa7OIGF0oX7f6nKwIWc3r6t51q0rpOQ9SPKWAp0YmFgUQsc3kYSekLCKrJMT5
oNyj+oOvuqyWpxmWKno+X+xF5dFrdgZDnYyLwcJ5B4nwXpztyUL242zkad5vDWKB
gtfI+ERBwfV6pHl6j0jSdiGc/Y91TylWRf28Lt9+5UMzrMzUipkcuDRvg6/YjRzN
+gofqKHzD73VV9yGlfEMjkCY5HfP4528QeLceXAh8W4YJ30MpxwDTKXH+0nfxRLf
LcWmw7cTkNvxSQTvLdKqwGQgV2ic8eU9FqnB11HcAZY1ky9mGOMRvNyD1opVeKpL
l9X+uBUWRvP9rEIkf8m/ZdTfP8Mh3NLwIuUIgfDpztE+SOaKzqzRPy68oZIpk6cC
zVw9SjTxfI7+gv14Edb7dQtNPwaFK6fbHR0wkWTsva4fbl6Hu7Mdr4kOvkFdK6jZ
Me9r9dN6K090HgKsAjbEI9tSA3Jc9T/G7j7Jp06x9YZfF5Q0WcrfizGz3kyKFt1P
1mpFWQ/KpMPfDdzY9LKl5TS5l++Nmmw3KdHhPnoAC/nkbD3LFYPmtj3GmtH/8jAL
3FYtUrlJKtTSvO9nwwlmOt1HJp+AY+hj16HfIgW+OH6ooqK9sx1pl26iP2OSeGp9
jx1D/ECaWRfOLfDCyy8TT+o7yGrrF3FxuTn1wOWVLl9+2kzwaV7kU0IYtcgufba0
8lJcascRcVQEKd1pAhAklIPxJlPEbyXhTaNoI2TYLZSqz94s+4URA56G8DDU6kCL
p9D5OuNT7xRhUE2gleu7xFDJ4ximYjM/nyAPC6mpH/34UsbI3iBboFk2lci2u3+n
VooCN+xudC5T9G8ADcpdeWx2a58cRmlx8l9okEj7n5648UX8ho0R9R/nj6Ti1WZ6
6uQhbSkurZWLO+y2CrrIOLvJF7QEvWQaV1XdpFWeEJl3Kh/8vz6DnPxzI3N6HsDc
T7vtPA5GHnFIdV81LAlTNhXY8ZENQlHJhSikbUZnNHjMWlUw74YEsfrgpHIv8m9H
1AX1mxx1rdScVZa7iFZfFUmXbaUgo8bP3SW3G7/oaNcChwlzYtuGbY0+8AZ3rRlV
LTyOTL1pwgo+PSp6L83OgCA1R2Gney/UNuoBQMdGn8QprSEvMh5viGoUmVUUtxkl
D1wOYWF8SNfMh2pTNIapLR1gichIz8KcZlIhHqIEUU++zyCFmJkYT0nqrpI5+0Eq
S78YK0cRGrlftBvzKyGzvdyf2c6ZGPtq95SG+RuOYvMkCcVRHeK2O5Enf9PluJxS
nQWCMXj15bhv8Y8dffiesyRpz4Ib28EZOf/iYRWoU2GW/bxSfg9c3nS/Z0bwkFY3
/Jc6ld0wyeGysmMVbfCj9S6NII6QncJNy29NJxZCOJDlY+t2eEwQ+5T1OUF+4adl
NH7rU1c6ojq8P2qWFqE88FidZaURwWzIjVgzixECTMzA8omtzrkocmhLamq978/i
b1AFTwJjQxStRpbZGm1+7XXh5ddTg416lxSbritTTbc62nCfSx1Vt2Dh6w+tniPw
lBLyjrhHafA7KTZER+UxMnRx1RDNThAkVFe8TJAvS8kRBy7vXPR4O+hKk6x1gfWY
e9BfXU5NXzn7WlwXeX5S7WZQb9uhVdN5TLGVP0OysENX8tm5yCov3a5tEUgiI5oX
iMd83jREhWdBwcVjBnrAGtUROmg2oxEwfBJbJfj3noG0b3hAZpU9G6mAz9MhS+Lj
kjFtzmV4j0kMBL9EFo4a2ylpoYGdtu0JHEsWIgMwkLeYXR/+dMhApkERbCXuimgU
GnEKbm8LNr1aaOrjH38Ob2DSRueVIu6NXSQsraO4vGmF8p2CY8qixgpUHE1Y0VkD
0+ol+M/7x6EqRnRN5KuO7jSCkXmwiQ1iCS3BN3PCTJ5Zdg/FsRM0IgABGwVuyuvP
hwlmVNYhS+/1pbWRYq4AmdZnHmG3dSXaUtdVczeoQ7+Q4f2hW7uQJWmLDBqwPDG0
lYOOuOELWjXbpoCGq45SbzYu+4qjTYubYLR0arSqDId2+50I9vZBna84QNRSf5do
/PDhrj4RTA5vRo0vuNN+1HV/cYuze73tfqriSRTj1awSfGUurCJVpZD5kK2mtmQC
4BOWcBXKcX6V8mkpeWB7sMngaRkETGUVyfBbxrZdV5QW/fIS7fV9QUCoNzSINbW7
MZeK6VnizLH+qk/4J9pJFiy/Bd1cL3/Vit3bVLvI6p4MQ4ftO6lkXRLqf/Kc2zsH
0N+ycXiZKdJs/oQFoZSP+0wmF/Pl1O539PD86Ijft6KxCRtzo3UCVRspn3CcIVi8
sU1LXPEq/mE/sms0KLHNz1gmPL/rVA4hPINEyZfyXbrFEtrPihz4HvKOxoWn4zb5
ejq2X9t9GxsC+29RdkAvUhgwFZkVDO2NZnC6hO1C1pwHRh3o3r03gcg67SICZiEt
ngPYQPZQG4lQb0DpTBtEcB8VE2bhSzB255o5w3d0BScu2q6xHleuOq5+hVL31T5r
1ENud8pyjn2XcNZg8cDEh5if6mZlmwQqdUdsnZp2Ez+sNAYW+zaDyVAIBfarSnyu
hS+ob6bbkVyT+DbfZogr4HEHYwuJBJ6ZlrGism3i/uWMoX8OsOqVYVdo3p2lybY9
CN+m79V4WH5U5Ix/F8dodFZJLmDf/jSGxAj9/RrRRLBU7FrZrVzYleCzZYpyttK9
gPNYWo9rcbRhrGO3maLKwGKarhZtA50baWIe0/7B7BGZUhr+kvjnt5AW6mh/dc7Q
cMHctpfioSgAk7Qlpg6h4LOENCt0CK1eJzZopkX5UA5MO6pQ5CoA6/tnClScDvC5
QUvzZ/cA0NnifZncKwuPlJSVjPI6nbyuu86T4dkiYXWbIOZPuRdhSVHWI7Cx+iYm
msOM4lxLfaUlpTaiix1q3KC/kGE5lucr9ZJIU7e8IlWHFaT0ys0Vnglif7X7Oy+A
YD6ilgrYiZV7hUKSSgZlLYq5JtAGAaQoE/1V8MvMbXobsDlgsx67X1dLFU4kFWkk
XnpCkRjnch9XSYgOCsa/rEgg4Oh2d+E3qxPYQP9SHS3mjd8PRrIXGqpSmsKD1oWP
MxNYjPqScqNAP0dXPv1ywige73eJrUWzt6uYq0vI8ZDVVBvXOg1tY4N33VZe5GuB
T03d6Jr+jRXbOL0IppmYyX3qmGsjLIZs5d3Ty8gqublHukZSerE5aQyNYHYFn04P
eo2RQ6MU+cQJsRFu+rOwyb2T6SXdRPa0D/JkRANmp6Pz00C9QxykWcsUiTf4LXNk
IC8TFTWADCTajFNg/kiRh5agKDZK4OY4lN/DB+20xRu1l0lR2KMvfwTVCjrUS43s
e7eCeHtB5ItVz0/hDN1CrLjI1M/zZB0WoFxQjOaFIxKqbNvLVp8m9rn/IF4F0x02
+WLMb5QO+wsCX4EPJbXhF7+/D/pydkvYFhsZGiYRegItMk/ZLCnAxmW1rm7SFoPi
NQZdmAenUlcEThtd5vNB+dIFh5cJXiSAeYOhME5VNWTcvPzxoIjq+Lgei/B7wjys
Whak6DESBTOjfF1MnNon+fd0b39J+Swz8MQidGR1Qv4LTumTYJ6Hi25ioV5ghyGf
gCXkbnit2OnT8ciYMWrK6U+51EX4hNT9oCI69Dn6TZ5qnuzerVFzd+w8ziQEF0WD
8MMFNFhmyE5227H950SaNKpS8aMU6kMAQgf33PIOkkH3g+ZegctzbX6EYwKX2Q/l
ZE+tgjaV/Wm1dj0KbrqqeX689X0hQb8TU57Pp0bYXc0YnaCKW9ETtUwFVezg5eHy
11lj7IupMxD0/U4q0tdhoV51avxth/GLkYJ4mv5ACblInW46Mp9kOIrEkMd8PnvQ
z3/2VE3GmMTPCAwkW4NzbcJ+qJOUt9PQJKk4jqKHgZI9S48MFwlnXLyIB+fDwh/e
7tayN5QC2a6+skpYRFmT7mY5d3Gtf17aMF20RLY3FAXUKHWKBgfPfee3E6jHCng2
1AV2ZxamTyFSL65i07VPgDYSNSSLr+H1sFF+E/Eyp9m4LyK3t37pAq28yudUym2s
RvtoK56RsrNwZbmaSyDlsHVVmabdKvymNjDtY1qrM1tIJZUWYq2MK2U3ehznPZOu
ZnR2BSAQ+HMO313tT8Pm04rgmIr8sAmY8W7GLy+K7gOoHS0QpfLKXl6zRmDyQsuT
LVHL6uEGc2qQkbLW8pBCl7z84a4jBcc4Pnd1cjbgTzpzpTAcHVrIxe/ZM6IjYIFk
9SUa2J+Ue5KNHOXA5bP7fzT0IgymRuYt9I6ntMt8aMgHt0UVLN6czLrr0K1RrLfI
LgLfzyxcAVZHoCoy7bKpG45PKZR1JzcfXK+iALwZqWbP1KI5hzDP9xE9Th/h25nc
KFLQu2GuEwQvxkLTKmn7+LhqFCpTaIEXhd6OI7xR+2i8AASOdERfwSo90CIEWMid
kuIiUb1EQWMXMSEGL8J9LdsClDy+sGOiNLrml9KppJZh3j3zLVFTLArw26V1Mmn1
BVkN+X82cob258pDU+cIBsfkvb9UZ1RQM4zSh8Ut5NiRs9atAvZ3MkJ0xWt6dZko
Ac7xlD/b8AdXeGUGd+FZ6EFUwFPixdV6Y+sOfqvblUkv2dcMUrMhvz+3RWmLtuA3
zbM5R1B+yRrsPU8V93tTsRXmxt5WusnGf5s9XpcTX7eLdNrM/UJacsZeBd4qnThc
siMvT5Uxy3x8Yka1+1a7+ZKx+k8/6LreEWtCujXEzewxnMSXwrRq5KtYUz/XwdlT
kGL+Vt3Wn3/dwmh0sZhKavF6onj1imb0ue1IzLDFt7gmlzaaTUjpIloHeGkDWzzh
oQmTrrYH7YeLcWYiQStD9gHc0O+xrgu6Tpn4n0ff+z5H+LgCUKqkLjk5zkZUy/cG
8Pyxt6i1bPHHT9yTfwa2KdOXnDHtSghM1zRR4m9Jg6pTuYumUcjnKVVYtQSVftmO
sH0OV3VwPuN01p+FZxuIcicpvDrajmhegBKXRMO3Hgpp+MvdXKWnubWz0kpFWvQP
ZzF7E8VnP3YddRIPEvAOp+g0a0DiL1eZb7GQlaqjt04ARGpDwI9Vl40dwqemYvgN
1eMFHybrqG048oH0cM29AfCVXeTS5lLi1gLcEE4A1Qj5/ZrQ3IFprhk0/3LLxg7F
l6mYEoCrnbz9+oypgHIo1XElBXxZ6a5idiUCCHQQUbnMzspZ/gPHcb8lE6CYSVBz
b2frVfMgnxMYCjkP6QCOTj7eLt1yVyqghbZzzE8gSjvS8+wvxeBZxQ0hDXS8HAk0
VDUky2Zsr8sTwmRwkCmhJ1e9g7/YiFlcm0CoIwS1jY2+0pHXMQ5iCiI/4zrDtHB6
IIYjmCrfQCRqH7/Syo1+pH8DuOgTc32MJfFHWJw3JNmY5MXEHYkmWmvO2IIHOBjx
ULeaw8IXa5v4ahYg9sc9eNTpgQ9d9DlqELZgHd0UfGcNLLnxmZq0s6wOI6QWC2pJ
o71sgV1VDl7KIt31XpDk/LqZx82ybE8Zvj/zf70sAGMmCkbpU3AuDapZDwEnTrm8
CtsXfzJstq1uXUsKBHEDZpDK930zJle5hrcguDTFukT35piw0BGJwIYgAhKJFO3a
mZCbyz2ZO/yzm6l1E0GC9So3fZqvSYSNcemn0FyD71rNKsd4F+CW3bFBdMETWiRN
hkuRdWdSWSFK+VTGcuVBuMm0n8ch/zAVkCcAE/ZkCRsnlbtesCLRlKMrjbJaNr2b
llZNp3523sq3hX6BT+nYjz446l8rCz2hT6Dls7BMdtCBabQgbXmrzzLSO0ll+UF4
1Hef1LI4jJ/S/aP+O2UizTTVgYLnGgaSQzm8nYzJU2f5aSaOXm8nlEWF4BRMkMQE
drYccbTlNE0ERpwaaulNk4G+CCYltf04YMfkutCQYSuhhVyo9d5eEBenPfiijaA/
THLjkRJTt5C455LXGhP1lxFsm5nm4ViVvmwOkVbMljt0ybXp8pCmhP05BNs5cuIC
m65iT+eUj6MP9IxPNZAtTzgIpmKyldwIL07yObtz/hSg157332lCuzhz+npdrN/O
UTp73PgHzzTmJi5HEJrwVlXmfKOBjAjqelOMtJpyFLzBm1Jmnnhxv2SDdPis3VM4
UTwqyNQNuZoou2c8HczLnFsH6lmVfd3tIChs1EQR2vv+ayVUBfIPJIPnZ+Hy1jyZ
6og1RD0aetOAtPh2ha3jlwjoqaNsCbb3PYZutIkCdS2xddg6rnghtd3nIUvG4SqU
R10lkCVmlsax7j6nnny69iWXfnqcZ+7S7qRpHZCoyTOChztaIe6oWdbriMoCMqhy
WkMefGMyNrbrOuYlxq9gqkkf92a0IZT3c9210a86dv2U25RXWhZIqpN3VcEzTE3e
2fPIlM80jE48vkW/8+J3FsI9MOpO1j5F9QpubNbVUe1yVONAmZWzC8pW9o8ep3h6
TMc9kvFwC8UO3hhnme9Cn3SSqJEAtJQ6CUiQlbRPEmfGr82HNHLqIG508USRGhef
t6uR7Rj9anw6+UGh4juW4WZeYli0cjhv9A68umRASES5wYtzzrW6IhuZrhncSGOa
8bNffg8njVtf9f3slKBGwkQRb+ROIF1StSyui+xUwev2axlLF568xR9Qa3ydAfYw
IWdYX10DZE0Uzz0N6/TYvSYTNmqBqJieTgdOzQBloEodm9ij9asLRJ+umJ0PgWAv
hHMad1czjXKzlGlEfM5E7agO50PAM3VRdc4jTjZCZKoXYN3Z9aMJXwE4sYNyVubD
wguD+lC0ySEsjau2EHJ4D+3/idguyt1ayy9TiTbrWcdF1A2lXMlfm3Lp8ZMc46FS
OPW6LO6s3LwQT7R/HEj+DHz8KhsOdqPywXYWEGe7Dcm3uspFoeqRsIJFE/cx9ych
7UYl8JFZdp2NXCbjCEAWbjLR4Mwe1QbZDiI4+0PbLvY04xqDgXtJT/wYEgWU84m4
ZZ5mh8CXFIy9pEU5R8AOa6DviXv+Pmy+uXNZ9+CcL/XMMm0ENllry5+7F8caQiXn
ikA2KqIbkBrkngZscc8lFmoNwiBSY2GbDmHG/e+U/Kx/j4Xhc8Rj81oL0tpU/ptX
19StYjczYmFCgHQqlwW38MxWqgOO85JokRVkuc7hgsERDkATt1Ssyao6KyCbjM6h
HGq4cDoIb2vu4QmvVZ2pAwsV9TliOaBztGlJ9ihNqvUpNc1yNTPgoJcvwoRB/6MY
Vuku8Sa09Za5mtcZXcZPdOKXV9Jiq1oSkp90WladcOMbqy2UFW5KWVlLzEM6XU5c
7Yk0o3go9nb8kq9SS183hE1u35kmARKooyo+4Uraf20t628z4xaiiKPQaN1EaKXl
Bgbdp7Iz3X8epfYo7JTFU6p1t7ClVUJd8jGzKQzlvIn21MVyXxI0bX4w7BB5H0Ox
aOP/FZNw2QFh+NQ0Qfb7Le2gjb+2o6M+MYjaJgoKbLrXCLR6Emqk5Bt9dhOdhkWl
j75LoYLTIYCB6ak+vSt1kKebadjnw1tN+oqt4Bv9bQNHQSUQpaF1D14RLCeJ4Upp
hPYkB0I7aNgiW05Gnsgjb0y+76z9EkVXy5XopfpkiupKxHmYD8EruD2ySQUYU67B
IOiDmARuVQUfUBWP13JZnSkh0yMsCcPsBirnybQ159h/VMmXepkQzFwqFbcHwRVc
XeuPygDZhEkCiJ/uRv6hgzxFLSTppNvsOf5DNqXEVLgcCC59aPEoX2N7F80o5r8e
sFJbEvQGt5RWKqlyy42h/OalTw8JbpFQkEGhIdUabEqPvpuhcukwZDc458hmSeBr
4Vlmzi3HJV/eeiv8m0W6eepTW7qhAaDm2aS4xpP1uRA2DZMU7qq8BPQWZT4WOPf+
DmiLcgNu6o7H69llkm9T8y7c1EP7Wsy4UNvEI9hQz/CZFY2tk0Gbs+BS2TPRAdMI
iXDDL2L0PmLoG4xi8MN883s+sp9KE0AHxbe0Sv8iasqGiYSmZ6tlUEE4sBKxNkbr
PjCRKjVzEOR8I3Jhef8kra+VH4Ecj4T8QbZ0ier+Sz7bA5RoV0CKa7hIpdmreZb5
cjt0uoj+m0IGpf2LNRhjrNO/nZEEIFIkr/pJwEW4ZbShxHahVkB1YjnpktLBFON4
YPeUgxKvExjqSJ3rT8Yq3+CfRe2FrqDhH31D90BljpQJwDah7uMEXoGZClBhruCg
XvdWPsYRocuwuJ8J8okdlDYCAEUWlCJ1KLVJzpp63N8LERNkz3sfg1tR8j3l8NL1
MCotc3clm4a9BGvJ32cCgbmC2BC50onUxkFmiGTKJAYGMESNZ7mPhr+tPiLvJj8n
M9jUrKjIkXf8owN6dmAgFxHF2vNHD/20a+AX8oOTLdbW0gXQtctA4G+ZsTFFJOH+
ixjLvqD4y3WAtjbl+ZrybXy8/k9+Xr+5Z+vxEu8lsGAjH6FWSC3QVgsEguEbywfG
YY4lCL12T4c5r4X6GNTX4e5G2CVYfRd11ISf+RXhz45SWFZOQBE3BIBmC8INIvck
D+4u9FWRWAatj/xCtUsg8xXWbJrpZoAyeJprcawqAD6/j6cCzxXIDxR0MsBlpzvw
lZAhND9YByBmRe7eqLOb+sAwrQYkGvi1s1EhOb2VM9ChyP002JUWDNHWSRA6XC0V
57sW8ZmvuDwXfyn9E6ZA4+ajQCbFgO1/JRMKKfdPyfi+SjVDgQPq33qW+bSEMHMs
Bqug9QhDSPiKFjlWiVxO6bdm/4lTcAdALA/rbB7t+01MOFZk1T804+U/dmdIzKuo
4qGtggg2b6TTNldN8HPJ70lMXZQUi46D8//3R+JMwknIl8/y3GQOR8A5gw5RYx+r
7hOXQWqm9rj0/mO0d8AokUr77a4mER3uCMD8mX78HRL1vG+WeU8hiUNibRFrNv4s
vt7RpqzZ9vKaul30C4JAZfnPq54ll8+aPafk5Ns+77IZmJB7SQDyvakxdO0KBSX2
8o/zSYmfIHTLtImzZWbvHmZ5ZkchBJFm9C/Sjq0Uc+8RjzvU7Dnoe2wnz3URsjk5
H25uwEJm0HcpsTsTPKwQABZLEYzu+sACZAket3z1G/il7k2n0Qxbqneyx53N5jI0
husBwLF6Cz9UKc2xUidpK/BGzqqruSir1ZlKH4lT/3wRgmdLBfQL6UDAwIj7w64L
Y/mMLvPi0fTAPspY9P5DEVoAp+bxLt1HK6O+imL9UMmzgJD7g37+UvQLN0rM7vKx
rK3noEG2Tq2+p/lnvxpbBFjyZjd4rsagsj7aIxBuHUhoUNGFiNksdf/IYQ2dU/KK
Ge1mUC9uYBhs8aGO4kdpLe2mUuJODTNe/R4NaH16i0VPadBHDD/8+Q7LYRFhNAYd
aAZ/+g5DlILHr+oo2PXBRk/JueBvDXkX5zkG4wzv1383ey2lT62EqTJQiv0Usc+o
VDLcoL+HRGilg6Zbuk+CY+YBQtyHcm8lxOia9CXz6uoghrZKDTuMcoBmvek/GeNh
FaBQ4thepWJF4qY3zkqDIlxMm0v3LNVWFvMDL8OVMGrbq7GKyo+1Kj871YyypuSu
QftqBs1W5Qa9DHlah3fthW2Qt4ZHZ17TYTfjv6o71uM5eewEr3oStYSqpjkX70zS
4+DkEkMpZ4qUVTREzFiw56LbAFb/fpIKcSTSEwm2336PuekX9Siw6SMGclLIg1S+
4tXpv9NbKvatKnnKUhLZPTF7k/G7Y1SJunA5+jCqIeRZhBbbL4//XVQzcTwP+Uo/
Cu7RuQgjl4BcH9vtuP/2xPSoFwkiUjJ0x8ps4nSAAhE9YxG1SQoH+8QsFF6fQkCJ
CyFMNlhSnVG/Xt4X+4fVO8deO94y3JauqeVdiDnLyQ2pQ5Dm6fYVvt/MJ9pDXpqE
5BI09yHJwGCn74GFf04z3yuDSq7uOeMHlsQeikkq/q/2qkFqdI4tAYLfc0ZGFU5v
jkx7+MZmK7qwI2Rx9ok8ofiHNylNubTq8XX4zb1MnzQCc9Uhya2wfVou9wn4WbsE
V3SX2HN52dGOtxazd0g0NASPgpVeWp5lJWZKMl8SEi8p3H7mqmgZBncA94VxpWpC
K9hfqNedesbufgKADvou5TSkFSuI8ECljU8evzki1/iHl9G14jRUDKLocpVBduVp
lFvzU0ctHeX1sBmKkUJpneKrJHGD4mKBY1WSfOCKsegl58mAdK0YX49i7Xsjp7fV
2A8ner45rUq39FW6a7qo3vzGBNBqzQSgd5djqNXGL1bXAN9nyLATfnCUAL/7ufLL
vcPmSEEuifB0IHfdmQ99QafP6rqNzecrQ4Vspc0r/AiBhEzyj0cxECFDYhWr260j
GYOo+1PC6xbS/TTXMNPkFuIcy7wMzyRsu2Y7Td0dnx9spgTWjRLefFllqJ4Z0226
xKJiXBse9O1gAnqqhq9h4tSnXMdVClOsmrRh40EJcbjEVqSwKFRh1H+w8GXDQsY+
ZFIo9p9L8qfXBioi5NJDC/6vs6167ghML53uYmzq6cYjYVv+0wu53GHAu8Q0DJzw
aK3YSWx6Dw8YEVdZNxW19qXMk3tiN/xtN9nK1JgBNrH4wSQFdUvfm6iYSnKvcT4R
6AhlwVdoyoByOOHCxyVbRjIBRzzYJeEi3SVGkK0BEsHPj27KA7VkMbgsHHYfMSGY
F1ndmcLWRQ4L1GKgdMqrl444u8DaJDs5ml6p41YheY19ePrLaZo74wys476dOSlN
Sz34bCp7sxfIjcrU8M7ezjC2rTtHpeuLW6JU56wK6yOhJRtBuDYYzPZv55kQ2Zko
nz6ATw1In3w55jEkauxrzwcOOzE9trSoWx5hT6f5TH6OfndZG/H6y4ugD8KOPYMN
TSwdd2V05hNRGJPyeW+Y76jex5xSfAh+Lb5xZa0ouZcQND6n7r1NIC3yApyaIERR
1q48SzhvczPgERPQ+YEmQCPGQ+a7HcGjfcazLNf5+FDHBwwOZdDrUUKonJi0uQ5D
QNyvJVg3bkuHTjzW0ccxORIzUKwywdlVillbky6HV39/ZYmeABqHDkxw9TL5VqTr
l0pGhDkK4R8ZvDe8z1T7wK54yGHNeK7Aprajf0X48uhy3srKpaMyEojtQ3Dz9fOy
S5Q9JVyoPC8BrePsUIgjhrU2oTOMrFyD4hy+VL4HPhwE2Cgo5Ce175iVzGa8lQ9k
C8nHPLhvCnewpz+bjTLegSfcMI+RiLTcXREDzVdvoHC58WWq3obYhN1cYUEQg5TS
6Al4gpOz7YEXvNeKLgFZZ/LAGIMETl14Rm8sZJMdVZ37M2yH9AZau93A35aOT0pc
RGJzLUofYmM2BnRra5wMlxa1Ofpg8XGXTIwPzuVzb7fcuGfHzawFvYLI2A0iRRRW
Wszl4b/Rbks9jpiVnFkIfK5scgTaBHEIfOXpVBjbYb8LROkdorw0Gi4W9vdSTfY8
tq+hME10LsK32feqpkkv+AXzVrWVnZ2IN2kzmYOzUAirs5EJpfUzxVmxAMHDIve8
LWirXJ62CP5swIRcLLWkuszMQXoH8yvwy9mZAHsRBfkxSdR834V4f/9lC1yz2lAe
3HIPtayVlbCvHZFTXkY71YNPWZ5dQR+Kl5unlPo3rtD6KQhiAFzjX6dYhoxUmDQm
Y7wToU2MU82+EqsrFSzDoL6+raKbORnZ+3OzDkLxOLbqZnx2JzLZG6CWRv4ruxep
sUeXZiVWh/8a91xgIKNDWlXMjeCXTIy10RVEw86wJPffARkSLj2hEZPYOK0q01Zw
YlexcQ7xNA+IfV0nMkSu51iuhgHWgVHr1C6ILDC8/hQAFYP/nWs+GjaVnc35D2eY
FQOEspHl0+vmzOd0zV3tB4KCVYzBbkeMjinoXC3qYBx5d804sPEModimeYdKg/+p
VmD2I623nxBcDKwoP3TSfCBUQpKQq3hY/xT+7Wl7GPpgL+8cDvZ3efiWDCRsTVrG
BCuHHRzGAVM6mcE2jErcOR249xMoT1x0CBgcJrXsEOTHB9fkUSE0dqLsOh+IFO1M
+92Y+yc8tpODL56djHEaCA9wMyJ+zjGF/NZhUB25cx9mai4ILl+8yZbgeIpRQa/V
FnJmaUq7O9wAhz1Zfe29r7U57pGeL4zxiDnRssgSnaUayEesa2EUpix7nFyCziQ1
BDx0YIRmH7wwyvT2PEuw8LyIhbHdUuPFGodf7ZbqWybIzeEHpxR6jVVUnaD5+vCO
vFphS6IdN8sm/cIT7ADFUtBEjVGW3esT9HWxLTsOdTkVoBrjF/KLYUaBmwftM4JP
U5R978dTAZo4fmSrleS1IgCnqbQPef1FuSgSGJ4jGw/gcsrLEaKmqH0v0ssFNp0P
GD2gEbVgoMoKGXtIq/ROs0ZyOnR832JEgJ31FwV21OlfqkArdiUwKPLPsQoJMpDC
TkxmAtH9PyGl77bRbSZAsRCb9wJFw/gOH04ukF4cxAhFu+Jo6nGILEyyLShXnPHS
gAotYNmB6qbm+u5/mGGxVlssZvIjyshe80rBZmRREnKxGXYv2YsdTCeXqwjj0HXb
XEmjKZJNmNKDH8qYkeVD4MMgWNKHAH7JSVRuG9SxpDTo6/RqBz4YRK2fHca1NQon
R1+jcJOGIeIkCLDD8kljs1bzuvi51xLNt0DzWW7Q0AJAHwi+WTH0cJly/HKCClRc
UnUBQp010L7MICEEoc1XUuURp76OyPwc3sX91BmVox8DZwJu7OpE2M5/q3Q0O2DW
YOYBopdC6IMftnHL63nmsvN2sj7b+HmSYWLml4aYtJeTSrU0zYAsOzYEC+4RwO+x
dYhYCl05vosJjBATZiF9pZCUnRyi6qAv2Zwbt+t5Z7jZkNXGFhJD1CSNNjuZzTB+
t7pw3e2DlxJZr4wMAAE6m2kTLrHNLLJg4d/ymglD0JdL5rP30vLe12iOc0evWGXJ
tl5xnF4lb6R6P91DwS8QVfQboKDOupGZLm+LESPbE3hiTDvpK3LCbITNSA2IXAQq
irH3VZk8JW4iOV/n3N9If3UcHSXmQJSKK958QTq5yINsJ0LPD7Twg1r4vZgezKCN
KOInYMKuU9i0Z66UJNLPPBLGRdeEupAEikAxbmTsmtK8ZNT4HKSphw2K73FDlj+d
lQQqtXoV+Gio5nKHeNKz2boY5hzJtdAaO4dKzPg3abdS3ZoMIGF4XXwOafLFDcsr
vNfENy+X5PYcnb7P3dOHXGA7VOwf7W7t6meFi5KJskUkGGCyqDlSIvbgYfbl5KDS
44LgoATuPuY/laJtWd+U0j9bxEvHCTcROKtGTr6cnbsXzc4WozEnOLMEgXLDnw/N
rsNt9b+JI7DVBv2E50k4z14IvUCtBantfi0jYxk0G3lh2ZlA+Y9/pnWTKGJSNcH/
p2QFKavOwGJSkQkxEsZFTNtKBUBex00Ggejb3sl1ZzA9ugTX+hNAqxeaaUF4pg59
MgnCNfWofuUNjUsVBogKqA5lZTV5qptESWTBg0/oaN9n8kInMwERUB4TdhWR422V
X5hDNRQoH4SM7/SeSTSHAUO4x/ZR2RdULadjpdiw7XIeBnqvLYL+nqDaSgEq1XYi
pAZK0cK5dTvkVjRp+kbv0+rhXX4oLxN3gYQv7TjIFe+8++p50u/cKhuhn/s2P1uC
Q3oalZCIapLI3vPsiyItBBdud3rRBXNdziKomO74snpeZE4h/N1X5mkaEYZgJQ1c
wxPTZ4X5zkSIeDx5dHeYwIDpFjBGFOgSmWWbkwzWqM1qUZVy4Pq702CHFF8Ul4R4
+ZxQIqdyp4dvqF8UgeN2cvuk4mVER+YdzMlzrTja3iyg6l44N3l/mi0uMMwp1o8J
qNHk37iHJf3Rfz6+vHK6KOn2ZrV9ItmU6FBPHZbJDU88MQRnF6nJ/TIgcJemzLmp
niYtssNjge20xj2R9oeDsPVXSdsiy3glyn2szy3dxEBF2kW/b5pnFNQr4/MIsjH1
C3lR1ok+fJ+anMmTllbRA5qq8zrkwUfwGCKtQZ8Aa4QxZVk7MAagKfYx5XSLJeHk
emhKlg8Ks1ZWHrnbJrtb7WxixhWjkQHu/F26H93uQgnJvhE1Q5Zm8mhUynG7bG9O
fumDLo9zIA1fgbkKZ/g8u6V1d+EwBA4CVh6XLQoonR9Mt67mPXjTBQ8PZtiMfbxb
fogqnD9qLauQl/8K6xalsyQ4GERacnhH+KG5GLpsvk5o9e1HKpUiC/gzx5rd6sZM
bWK1im3SIUlMzAS33sd5RXN0y7fByNKwt+djRk6vv2+UKTsZl5oBEExjHpWxgpuy
21v8A1RKr6+7kNqEaM/uFdrrhe2q14nGAA9KCIcJHf1CwEB3IqQvG9UtpwcURnFz
DoEP3lyx6twjWa+q2EmQBVsF5aSNz0Lv+hlP9U8RG6JJX813/lm/C8fJUOGx9Vsk
Fgj8RRsgGIoBYURZ9/Im2R1rmUi0JS1XD9HjohWHMcTkO6f1LjcVNMIl/Tr5GLOS
uxEORPaSR1AjBoU8Daqxc1ArJN3dXiPAljoVhNj3Z5YYS6uc561ox/8p/uU/ktGQ
gL0KOU4H/DtY0vtyqJ6+YAvmKS6lGdXmy+MkPUmOiM9s+NRPXeD8fOPwOLx4DLD/
uld01E0wDbTt66PUZz5r7SnlAGLijbkcnc0PtaNhVNDnCQh6IWG7R+3UGcaXOQLH
ur+baEYj0fLqb+Hd5NsENKAD5Pzbkloil2Oc62UFPKZkmCUrWAAbJaOkDGvhqHhG
V6Xg1C5vVScH+7Ydif07Y779MF0hHa1SToJfxGl1r17yzO8TA0ksOWoBULqjHl31
vLUhcg82/GUO2Tx7KNc8YTg08aYHFGjyAW5iPHHwvVrE48CPSy+jhAyTasuRlc2B
SVCLhfVvP13j+mqC03Ujj8Sd1Z17mlPD1XHyMJU061PmlKuF1VgsXIM3PvXI6gNk
T0Iptn0S9wpAtHMVBLRsjZTMHBZ7L9hWiJL0miOvYAkxyZ6JlqQ6UTqKSiQWdcu5
7Cuuc3LH5bCTKUlJGT5o7pFWiphRg5yMvULfBrgX0I7U5/OHbwU7qJHGfw30VzJO
jpUScNw8zdxTV7BBsYtsRsAsXc6vK90YqK5aQY6gxu2aVFUzxVcCqwofu2Vuws3q
wh61SBt7WI/OEdjQe5DFdLkIVU1K3DlsDuD64YzaJ7uTU8PTNW24+dOvR3eOQ49r
nYjeXcfyxxqp88wnFY0mGOgKrZ/2Zx/9W4GjSvwcPJVYBgE2909OT+uoqssgo6GB
kZkQSRL2rdiRZAxiYGTdudgVhXIy2lJBip4J8odjfozVNpzgYqKIePw0PpfnKrhg
hqSdtu8fY59/478cjXmcR4FD3Wy7giAyleA//KJIrhkN3Vf7GVZMZlFh61oTIHJZ
jUxLZwvT0JQ1W3rt1Q0c1pErNbzhrDaBCIVSPMDgRbsjH+P+LyqotcSwWR4h9zS6
6no6U1tHNMRD90RO9a15mRm3BocU9Hj1KkFi9ENPidFotOZMDkRvoQ+qbO0AWn87
6D5zIZo9HV/ex0Bg6uxtURDJTVpt3G+gx6vI7/GQ2RkE9dwN+VkDYgSICu5CB0pb
V6FSd6ooXHg1XXE6l2J2y+facH/2HGLoQj/PD4d+ZYdwYqwvw0LeKh0l/HNbl8Jl
MK1IUjfPzP9QfLB1W01paYDeFf6ZLedrr5xC4CNC+b+S6EKcmyg9adyaqglbKxLb
RyJMneCcxXauaXH6tf0rixToXtMQ6/c6WymcGZL+xV2eE6FuyENQCilLJ6+8h4Rk
zKF2wtv83PaBHaxdiAtumFX552PsWJV3wzSzilfFEwfIqN/a5xdI75+V6kueh8Oe
07RAHxVC/KCeMg33+n6SifUsR67KaVI6bJji4+/uvMoEZWO4/R+u+zq/7C9/1jGS
GYK96j5nFV5EMRKJLdMpDR7VbBlEd5KMC5hLb4opQqvj2VuAI15tOOcibhuZeRcQ
i/0kwBC3gf646f/4B2MwIrKGfJnaytCiUB7z5P9ZpJL2ip10Cvt2iKaDwtJ5eaGE
kXDtFtXoU00lk2mxLw3eGlfNDVILtJm/yCiPxIEeS7LlzRmgL1tkWV6GPRrayDyE
Z4wBBO0yoGrUBKG0ocDjjKUy7b2CDs6q2XV5mycCmlgIB7cYW3BGVp9qTBBf8QlL
5Q7nw+gxSAdM2Cv7D4E6C7Jmat8yTPRK8EH5pib0ZvlOTJQX8JykjuDYkmPO44N8
Gl2pMql3B/r0KXLdvxOfOPDpdfwAuqEVqgtc5/87B4IyvxuYUgeWjy6aI/J+ZOKY
2PrF0WTJELF6YFTNcxKEVuFtgp+/zy2tV6vlc6sowHLb6h8rh35nnOPIBLGWQmrQ
19iqG+pOrTuFMwlhK5usZmVVYAFyZbfQfH4x5q7KnVz3g8XwftH34k6pX7Wh+xOc
PubDOKerYKIdQaOrRwIy8qqgH8WYQ+WhFmKAtPITdUg8fk7jDfVHBAGmkAn7iafL
zSGwa7aul6okWJsHs2/Ki/GwwyL1kiQdCXGyiZdIliUzEOcNqPUjJ8nTi9eNh8r/
eGIuFv5YprQYi0ez+5/t73pBA0oLSG777L82c/g6q3hzHtdaPuz3m4VR+GLKzMh0
rOlfQturnYJiayn7whQuZIL8h8VYSBRu4s0SQbHbdhi9t3wantnI4fxkwTcCmHTY
QrJ5CAdJqe3/XqHHXmIsUGYbVNGGOjdzVYQFBXfHOTKqs38uC54L0+BIZtSoQfG8
409tHsJaaA3fdvn61ML1j8pUzTBXNu8ufdpcN5U2fLWKZda69/+WqGCqh513QDnv
WHYZB1rFCtT9QkpvaEro4StsxNGi2MeyLahJGNp1wfO1lGZ3KmA/hQ7rZRNol+I7
NKKSXysNhWTMA6XRl7k3kRxKDZ2tJZjYRedrlc7jk9zQuv6ivEtMDTMGo1K6kkYV
+Wi7dhJu0rSPg1oNc2009XfhaJKPDCF4XtLtWGz1kXDxMVC58fvn/TMpTONob06i
yxDuSA86KgS9JqpKq3CIjzmhfJCkhgARt9hHTZSul8bMWbwLIZbBsTsCN/J+lRhS
Xh89/HM+owV3YqHYxhznCfcWur9tlCOpJtMlHTFFYGIqm4AsWycvd8ZxwlVzuQ8u
o7SDA/S1266Bn+Wxe0TILes1PLVmkEAZ8YugEe2q4AQyklKuE2Pd/n7f8zAaxjxg
1L50sQXqDdyrI/UVlHu3VrKG5xPxKh4fqhZW/nHJdRnXMJ0SyLwQhYLzU0HWcGEl
ZCeDqlH/78j3CJE71EsqEm5+ilrOZOEiJmNNhXf9d1ePM8L6LdG1Bv6Db2e+c4vU
DVQSJRxlDciACmxvW7uy/k+iDkhTEB7SOEaMk3xNaHQKPsGBZ8/HenCTbOUo1c/D
5sdtWG0B4cbfXb0E4f+OOWF9ABIPJeVYS4XoFvE9o4JmmrL3dDXCEkuyw1VSpfbi
P2D80LYewD1QRd5cVDOSaE8I4zTkJWiyKOIsrVBiERZSElFdMsdkgGMF9p/8fmO0
Y4rSlUxLlRnIKbIh9hILhc/knsX+CsTcVzB74HX79wYHy5QKe8+C1dsIA+w0WPx2
U7CbFb24UR3RxpABiRJ1ONjkPng3XE4wCV966QeSmozw0e0+SWG2/+Em2nRz8qlL
as03Zt8ttpDHvCTw4+VSV3TXY/Sb9kcRZbXoYNetKLWz8CHFuelg4Si0VLvTIdLa
b7Se/DcQ7zSYpbr6z/AfQzM6Kr/vCXKDCqWJaiV1txUlEcQqtO6VPY97AXU5vaiT
GrNSI2nMmrBBW08tZqMUqPMucp4x/D5bUxud1NrAh8JViRIb3E3x+KAIO0oQYtgv
2eZxevCRNP2+jYidN2uLbqiyn/4hCOVRx9x5CZuaMi/jrZ83ydlVXE9L0Fix/vAP
g4hHcu5PVQ4P8X4M4WueTebUxG41z6ehczZLnDa7w7Ly7+5+D3EBGUnUDWUbvItM
8aw3EkejUi3EHyJiWl08FrpXpBWdPwjgj28t9ivrNnC6GQq0AjsZvcTAFJm/17Op
Bk/eLubECFI4HrKgq2ki5GBEDCo91USox154Ex63EgfqD6P2z+G0bobVQgYcjtzk
uPe/0wrlLy4yM2/ad8KYmfjVgkOtIhZuujV/u2Xie/VRCahHWCCbnTqVtz+Hy8MP
hSiGvSEsPxQLk5rDKqVwDMyRFIK8y2H5XScv0WfOfezcj2OOAxvqqbp/NI3k2h7B
1kEjVSgAu9AyJvxchU8cXzQ7Wx3Qt/tnfwfrNJmIhjQ99NIZMLf1YHHoIuHBRuYm
nSxwLcZh4uUvyBVeoa9X6Fv/5GNIj12Bgw07oZ/GYXZFrhwzO+t/qk9Kp88ubuVk
m3i/fFzKCu5P43pjPpbYf97DLgb4Lfe4+9SmK0ww2n0NU8+GI9WWe1M+5F7sizk5
3iGFxr3RMtwhgKdZ6aHzDxic7XAEVbhp3y0oRjCrrqucC7RBDaEXEt+NrUUHAPVz
yHBO09y92Y9GUlIB/+EEH6AHPRCae9JJTlFVQSxXo+QsCZ90JoNdPrBVJnvhq3WF
NBHuuFTSohrVWdscz/NnLqakrN4zbQcwmsdLcsmR+dnPrSkf0nFf1r83SnnLIO+h
8Sa1OqcU5CUsE1LxNwWbK1mBbLpEtvyUo/7+nALoET/ZQKYBRxUUEopzgPO5jcLR
hd0Qwz/YkJR2Bpibb9wnvZGFeAiPd6tD2R3T1viswSf/RYqRFp0Ha2gPSX3MstdP
9Oxqs+49sucZCA10jd/y9zK+LJ8SVg08bP/cZ7MotCKKVzWJUveqOYFvS3azH9sO
JDqSkWkT4kgDj9Sf2W2+qa3wnyJih2s9zhb0TBaI+36ShZVKbUB6fnDI8vNcWPjv
6qG+srDlDMkAeSGpXHyRALsdv3yxw2vSiCDbrXHB4vJ0k2bK6S+2elrEOzUNuLYo
QJX1GLjq9hvmMaOYfmT21kPJY9cG82ikYdDMCwfWlE8TacS7N2T9WZRvsXiaO/mi
GMydfGUVyB16LMr2/VYCsslGHI8yChd94ePKKWS5pwnfo5TDwfyz5AcCdkGRbvAU
kV9Ltfumaa0TdqHr+hQW0oChGQSpGL8ScoTq36K87GPDlRzKF4kPDsN+JSmUV7+S
HksAS9D9r/HTVkh7IGB+q0YoZMd9tTDXvwfqOB40JZCjhCrHO3cH2M0Eiaf6xaBT
5Sj5nmcIYgpzz1XuQubBC5Tlh16mrYJRM2JVYlgOraL5rAO6n9EXlCH3daomn+7g
05iSzAKNFXm8o5mWFbkfFUnMGXyeWuukK/q4DzdmRJcvAaJ8FBzp2AL1OALr+hrJ
5162BkEhuotgsjmlEzb3bGzqSK0zmv/0Tdmfp5rTkempMNa8OfQG+pdpVRvDJJBs
cFhKua8xb08KpD89l6wjZyLR0c1lfZWZXKckJmyispqw2atQRiBpcPu3iW+tvgE/
tnQjC3gygwlEhk6Ilo5C17sKdBhK8BlEhR8sSbUVe/XUiriZ8yiSiP+lYwjSh0AU
9V2Y8xseOnr1lomqP1mWYC1RnPRsvZWYfoEebvdVYqePMTRmKfz+MiWoVTkXueG1
2Dac3FW0du/2eDtgvw/higZVLpP8T3Yr3w7a++UPBmfPjeryw+uJxhHrhlmhYnEU
bepMTDi8epJ8P8D5DOlaDJ5C7UYw1Y0mapQ4Rs5imSyorYpwR1UyP3i8YCzC3ML2
Af7U7CqjeVFYR4sxM/044VZpq+3z8aWjZzJ5La6dH7LQ1JabNj6tMijRkbxnQ+JG
e7/1eCCKCxGQ4FNpgOxysJa6lU1GCN3paMxZFk4XKA6KCs51zXwSm0yT1CFJicxY
pODWO400Gm3rStlL7tpVnvBTzk4BqRX7atsAqBKP3QcRC6UPf4/B14CEmJdeicPW
XhazwOgfu8XljpaXtSPx6pD8M2caAw1HSpf/B9sVfxUo/KywTKxVOYcF00euFOQX
soKv/QDKriGSOgQaSLQnydpEjRJQgcBbTFBBPKqE2KRm+Q+onwpghrMsTLHS3cqz
ygDTAqSo1+EpnjfMGc3w2RtZnKmnPDi1wCMk4zwrxWAKItLGTA9oWxkKfCmBHIBP
Za2btwKeiXbtkrrBcHepDFNHGAaeKd/p7Sya6NCldaTjsuqWRa3F+DGxLDYhfZZF
P9/PBWuBq8BbS79IkoFcEXme/fOIFVWT62NRlqrSh6/lUzVYjPJ1paFATNHtHpn8
`protect END_PROTECTED
