`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UHu/V/6sMKvMpS5KmnCrFEgYiAOqXD8JJL6vq8LHOaAHfUiWdrWpDrURnerZF0bo
ySWofYt0+gSCH64iCX+s4ZL9z82VHpt54kJeCOhfX1W3co2YCxmX1Q/4utAh0jUG
xqm7gFURGewbrmI5ybBUfXNi9N/METdQDjZ8TFlxfq1082usS9ffq4wLRUeiK0Dh
+Nj09BLKmOdlnA7sevMRPxQtYbhReRoceWxpTkCTYvFvvLCQMh/9UKB9cqpYB/Js
VNIOK4Jep5NCyFydVjv56tGQo8t6I+BxrPEgVPlxxVDlO51gYJtw4U9Xxjq+SgTj
7GxrAm1bzcMBALUtpCRHq70YsBfFGlaVWNuJUaaUyGwrIBkRG4j+dMjhboHbP+Sq
UbRrKwV/r0gDXAOxa+ZuEhHNHqbdOonvWVYPpJb5BoVqbpc4W3dV2srJmOxtypUi
BDpAGmBcNm7yZorU8WIPW5LLa60DvfDbeYXCfvINX+6x38IeLcfJYLhCGQbMpynD
3YL3rTM9z0qIpvygE8L8ANxosTf+QpkNLBpT20+iEv+vYYH3AGiXw2662TwZ/3is
AWckM9G4G+3ybMe/IOwWYimQl5FolSgjXmlGnXG8B17mPJAhNqxjdBqKjgJhIJsq
sKZev/5XB+miaKEn3LYzw8pmHdMOTKxu2G0fkn2c2874ERVui6Iv5NOvMYbmWBuE
BYI3qZMKN4ceojVOyGpoFDIHEfSDErN5dIIJdaKslX9hREF8LpDjhURlezbrkD1z
1vLTeKooV6ExJTjOHksIMeF5uCG8HIgKO+k+OApv0jnSlhyjnX8dIV4pxFW5L5kQ
LQwr9Nh9N8CB3hS9vNmONqcc/FKoRKZLf8ba5Dqgnw9jkuY5Ttragmm8bQMb5hj/
XiiaCes3ZQCcJ4aTInoMjGOe7cCPeBdzqPiXduFJg8NziDMxfKyuAT6Oytu5wSfJ
EOnlFp1UWc5JMcvNQcfvy7HyHrPgZ3hLg3SahHbx9ZZMKHd1eUeMlT2S1DLkCGEJ
/cnTzrZWZ6606Z139eZTALrVPux/Stzp1U+6H3GDrY3dcTfVOO3LmFjQOHOaTGK9
eeN5B8ZYuwjLYtX1RNFCYrgwXA8+Zli7RBmqYRwoMhwkj7s4hp6u4A3uJb/YnyJ4
xO1iO/tfMc1apBgZGSFKwxg2RqisMKN2dTDzSMSDXGQNyCGPvTe8s7Bvwm9BoqrM
NoqI0NxyLabNvrQGjcIT+yRLu0LsKqXH7FyjtrZIPiNJPIdgGAgGCfq7/6vULX2c
rzvqyyfPbFe9XLbudkJS3JVo6rIiq4OtwFRmEW6yKjCuBlNrovPVvct3BSjziNSZ
ww0kzcRAIulZyPGiS3Y2MKeiuS9YGC5oF1TiJflf3RSjxnmu9+kZ2m1qsvJhZtN2
sacXyfMPQ+nyPOHuG96uaiD1x08NlGfXnkDgEPqrZSFVRYSMUZwppNsS24VgREBA
+yRTQ4n0TPJv9NIc6KO8y5NFsT00yE7cfjJP/I6FwhrUrAz483C5sxuQDv0Eanup
xMRFoyCY/17PXoSUZ5/eNJddrBsXkw7ru9doGrIuStEISdWlFupt8mnaIw5uXoIr
MjoinZ8lHSlHbdBRyjIsm4F3Lvk+G87f2sSqM829ZZNkxSrBi68HqLSlnmrrFZKH
Kta7uxn5dsLKLHBzBMpchWbMh7W0YucoMJpMIPbTr8NdQUSh4fWjAITDakiTsGsg
+Nhw8ZXlOG4Rx0ZNbPYMyGJBMY8pXL7tjJuHKBL5TFRxisDKEWHGUaDRMgY+qOf3
BLDS9SAd7zOsE57lnoyM08HPnmrJEsHV6U2d2N9Fb2WakGpXD0nods2gsli3gAmP
+8XwYJMN2uMthbEykM6YNgBLNIGlsgVGGhsoJaCwyr702fOZ/isSw2GvcwMdRyJH
B3ltGh+Y2HBAdLBraAC7ZGsulKmpghbAtjngMiJeRJRmQDDIjLPfCwLxYbsmIzAw
1Rp9pfKCyn3kfVWaGe1GdmCxmYirbXTiSqf5i7JIz7t1CJdfGgMnb+myVFDCRkI1
rpxL+qYEMyhtb0Pmjb+Yd4iglf0NRyGLyl68c1tutAWbrcikd4pkubeBK6TKxYo6
N9SCAd3n6VONdzjH39LgYkCmDOM6nMrNiOoTqcvHTDjhCyfWVeJGJY3563kXCOLw
wziJ5cF1u3Wqwmua4B9yRxMYAXl/di+NrPAGLUAXclQfOx7wzXSmg0GPuSTb437X
b3rmKUSV05RyO12NaPyxVIdlRL0RLFEsu8CezsQLr0aQAPY2nm+bMRpm4wqxabXO
CPR9aVzswxutFAJU9m4jwp/ttodRYt0fOqbJRFXt5k/zDGx0dhFGEtYQOwj56PeO
D0+H9xRv2H/1WWXQzUbuVnCq2RxZAD/tevvn+MdBE2wPhzBcZmdvBBYSHXVcDfFM
40mDV7SdKyJcPWoPQocORHHptUhrhCSmuJb2/mkg2ebYhQhvVDFCaLMqQKQDAM/+
EnSMiFhRTbXHCR/Oe5W/f5jrnVDTq4Fk1h/gAGSaT/J2uHYfvVEnWk/GoB6XROWv
fG492YnTYsEUb0vJeITYjnWHFRX3xesbwiz+WWcEfk/VxQwtSopAkpENK4BmtJbZ
/3g0xsFxXQrcFbJEKi+i8I+NXsJ4GANUJjvAcAY5Sz+OEgjfvyaCDeOXlEQ2W1g2
7oCbe+tOl0Le0gDJ5LKexX7LViUVf6NOyEXkpA+SsUyc2BOxebqRTKT77OnWjxGx
pbJqS/QBSTEiF5sXXL+ZdHPRtPAtMeHfIVKTO8zsMV4/DRZGxdWRP2EsX15z9aeB
Ad9E9J6NLm88w7qh5AXHMi4x3AvX2b75giKI5VpsTvUeVJ3S5u4FQUUReh978O6c
8kdFk79P0eYEQr38xXHXMggziWLh+AFnYdYoXvj69XE=
`protect END_PROTECTED
