`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VfU7oFygvRCCVfPT2ponaFaLo8dw6/P7wwHHfHN5JKMVcwntUH3IjadICxwne1tQ
RXiOdRK3TyKJA1osfupuI/lyCRDigFrLDBLTMeP2SL/q0X/bZmRkGkBJQfWqoxM6
Esq9P/BC29X7IXuhgUA/1deyzMeHbk7mZRKIODnPr0MJAyvfVfpTla0A1n1AuFIL
SPRySWUYVSsynqpgDnVTTYuZO1agiayIC519ik3FXXB4vc/k2Jo5tC8SLWpu9DZf
D2DKHSUg+7RwBtzDdX0L/s/sBOgXu1PgjotzO48J7xNaVaH94sTAs9bMT60hHkXs
xXoIluwlWnee75qmUaeFrAJHItAWvyuJkOYbQrGDN2w6ZXL9pjC2zqXYL8/Y/pRO
LTubhk/1zGxXSo7YxtxnBSq8+RLgeyjQhQ0cVhfCuc4jQg7Z0IfWtrXQVC3QRXyy
X8BG0o07KI1/jpTm8tN7XQSOpPhqjYIg2jmgA6L838XvE/tL8FMNMaNVL84ECX09
fUS1JUlwmHlKyLbcsDwkIjBaprnRBegQ8YCOAs+TVy38fHGzbXmLNq0HJPqRFLxO
3pNYjYjpFyoc4OpBNNuLiKQtrIEnIps7qC6yQ5/nLv9ySWa+dMxuM3bwn0InFcRd
g4JK8r+8AqziR+xJkbXUTvLkG0VsfphoBkaqRjFAd/OuDn8IJs/4XYEmRkR+kgMh
yif8EjX+TSj3AQSZ3+l3RFJfqs0nog1VEB8Ez1r+8iYNlPlGneFF7UU/+KSspcBb
SbhBdZPO+optXffvyMbh7DH7vKJRwMG+cqYmc+5y4w5JAOUc62axUbjT8t2Vj1xx
`protect END_PROTECTED
