`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PxCd0QP1tSgLN23nCtzJba4jgCjJmDUvEBDFByz2tIa/quRuOmaGPyJpqvWz+BLy
qNgnewNcGsLpj89WtEox8jQHoxgSTGjx4OjrnqtMR67uUOmn21PPxf/QGS8RLeTn
Q00D3FBSc37YJgmMRl6YDhwRPLLZjGJ5TO2qOfGAui5PilOkcxI84ePfgJVW/jUf
XtUMA+pWcde4e32zgqvPFkpGOCsD1TY8rY5TQyW3Dt3VhlJ2E9sWUMhw6Ivio6+N
yPC93irmMqDB/O9cvNh/dFtdKmFhC8Sc4vkrfuQSdvTzgA+22TlH3nNvumF9wMYu
vg/kcwdqYmMdWZoSVLR0gce90ERB32HBlu58j0Ll7dEL5ZGjZD+Q+SxzBS69xR2r
zQTTezczQ6omTzKu4pSdWwD6D0vARVOSFE92TBNsuSKrHJFP3RX9eTg6yl13jYM/
kAOciIEWu4nIGOobisfmwONpxg8jYQZpk2tsMGfwKojZ/KL/5rrckxhBZCcfVrGj
S03zFOczJXd+DtP+dFXLqBMQJeplFNXew+lNKiX7uGmXeqYLYB4HcVtCVQiaMoHk
4M7gmY/qn85SK8JQNsGIn+R0D8pygSmQ0FXFcAy0a09EWxxBBzwnnw5qt5bgRiMY
bSzrh19kUlqhcP0fD0Ci7NDSKql65WaJbXKV4V+bjdBT6nWKqaxFaU/SfSra6Ilc
WwItx1Sdxtw3llVlEQ5yJgMLYXtd5IPkMp6h7WPaF8PRvG3Ikgtrh1ZmO+c85GI0
JSEhi7VoKcrFNNH/+3ZusUn0p4jqOyxvHs64dszjuHer7T3WUeNBpmpdobI8ipdc
gLsbaIEulybntuyQvQ+7uT89bNQkvwVJTkz2rRaPp24i+np6XvKEwRyzNpl9k+37
fUpT0VKFfuMbbkqcmJfbnO+Oftn5iNHwNGjr6HpPR3kaV1qU+YtzlqFNXXNDhgsz
5mXOZkx0QW5bDt1KH09Lrfq+d8nUOCrzyz6V9giMlm1YcOtoc9k8iKU/NV1VEJlA
O0lW23P8bnBc0MrgQJXZmXXlMEyFSQ/HzLus/i/j34z27ySy/IMkY8IotuOSGhtH
jQYTbnoYDbFA6ab4aDDqrKYDZQHfpKQIjoQWKAmc5nRnH1Onl7A7S8H3JpwuGOvl
yjM+whsaEiDiUzyn9w5K/vkYP/xHEW4GyFDjQUlYKtpl+n8v4wDOSJ2fWEXQzTiA
fvU4I5TzKsQk7pcnv343aptXNnwrEU6buig30BvJjD2DUFK/JcZ4IAmio+ifo3pz
ymCVfhpeK9YJ7hSvgLSLfFLboEVhzHWv14RGLxptqNkhWFZpN+ch20PIE1MXs4Kc
2cNdJhmDbA8QeKjdpf/010y65fnBwNTApzlL53ZDdPEXBlAzIOhK6YkwdpFWNp0e
mSHeV6fGu14dy2aLjsedM9Idb91Awd3ORgc3FMLeAUuppYsNQcCytnLuZyRG/86h
cwYoa10x5a+BlO7DDt0kkLp1VJI4tkY/lvdgaexzCHeeD+bga/eFlM7XT/9Ef2k0
T3I4gUd3fdCl8ndydyZ4Jpba1lk0rjabMKHd3pwVez3hqMTF6QS598Q93oT7M7o1
AP/+4ymVSU+qa5Ao/hCocT6XZ0sXgHHi3uejLPUaztudn5HUasZXfyh9UML+Qe4y
KbZofdRwE5BLQZ9uWCMSX35vHPSzHzVFNTTMafUcflusr+hraNz8B39tmMsczEGg
3cU2JQoduy/oABWm10/d8x117l52FsktIKFRMv6x380J0nFC2eQEXzsUAjTeoftN
gHTmh/+86HGsdgrmbOFjJ7JX8kHjaon9ClKaBvZnfb1lnvi4DxcSItfat+munnRw
JIEOvFV2u46FdvBG/mKu+2VWWh9nGtOCKNzvmd1qVO1M/iAIa1S91BRysh+ycRxG
J0o+xt5b1cZNNYR5dr56PI252kOCxrpQJ0I3P7MeMLc3xIudd6Qd3KWFDIdg0t9K
O7zudYG7te8hgXkLQuO8H3LvuvFkKVkKDrPQRO/XrKUwRbXEX9/m9kuNHdeV98Ef
zPJrkyNGrW0sX+KtN0xBVlRz0yQXTwCLLpeDuDCw7EhYd/3CFomhXOns27u0/ohQ
hwRhDcehTzx0MEKteNrqX2pKOCmtamrbzTFEdcbr60M/7LlL81kLAyxOZuQRJe0z
PA89i4jhXxdza5sU6cn7Dm6yNYntqARPYnCQ8tmBau+qH3mHjncRmf8hzMc6gxnb
DgkbCMue4QMrZS81/AgRW0u5yvqq0wlFS9c95NoNDhbepNcgSgF9oScxoOEGjDrG
5BkAC44RalcejSuLTVpphTlSGdAABE0csofLFiKmu+laraymev3ZGs407dYd/nSh
fJgq6hFN5vIcI+MWY0VdZTXvWeq6m6pWI00WHVbh+mdM1orSIu9gVnXDUrcAFfAI
NCYWryGN35H09SHJv7IjeDq7lDqzR7e2RvlFpezuWDPK6uaopWB0VHNh4/uL+PZX
/2Po/ONBxJR/ZUFpMJrEU5b39194bzb0X0fA3xk6ZcEmOYsUroW/PkHc2YZkQhKw
x00rE1mUKvTgnapE+YliSvoPsmZ8PjuKDfpdPkTmXHG1VHa5KauqnD9k3e7owKYC
RllwRwXB4LeI1B/qfwZ6/0qHv1q4AlDyjbsN4TY30dmC50A2DR6ZxZzFt6LTV/06
pkRZOLkxkUqxCZEZ1lBhiOQea6I3PIzb3nMUzMjYqFzB6RLhiB0of/ByW49hoPt5
sOkf1kGCkr/oUt2WCo0QVSj4YnPEdl3LrVTPu/gZAsDcrhuk23UkKKNG8+xNKLse
ajbPlIDYO+kdAuArc9sH3IhhqW31cZb8rVs8i/AJ7bNHcHVOm4TzfCK6KWnr8tJt
U+OvYwG6nKvvKoYDowf1IpgU7JhOC0xpy5BrzgrIkVFJ11Z1fwW7ws84OA9Dv9d8
Clfn9v/lZEluQCrfoiBUbWsoKEwUhQZPynZKJQFFiyEgYNQ2RHOO3zFo6fxY8F1V
/isi39kL2xiJ3My1I7rnpSyURh8QNtaMFlOB0rzCjUgZKA8R1Cs/D2einpjgGlI7
fxaaXHPLQxIVZQToD8mLvD1kpiM8GDcGxrMljyKDHqEdci3/TQ9pLpNQjCNPtu+i
1gd5q35O9FT1ovn1Xh4F+ti8JlWhrhnqZHDp0DPPkF0T9wymCzHi7GvEif0aiPpv
U7RiRzKfsQ3siQ/JbeJzbgI/LnJ5OC12LC/RLfqgURoitrjdVJHw5uOIwcF6KlPa
kcBNePlfetEavhUKEHGmY5BGLdRnx+T4PpQjRVyZEXbrL5GdiisVPVTRdW1oexW0
gEyZ8j6kAPmrd6uA0s9sKaBultzzTKS4XXMQteQC8OtDACtpnX9vfOeyUxCcViKF
SY833kZiM8aP4L1TqpfKzIpGoH92Ijv7jZjaB2gm6F9r+Uy62b9kNfybS0RvJylE
FvCLUcKR0TCtmIMvmtMTTDibIsXvgAudW/8f/9MBvHzpUujwjYLDIjWquPEOfOKd
3d12owFSSgTDEAFYDupl+vic2q3yHH2i7eo3hmDSRzcDRh/mF0JOYKQn8dNmsQGs
Ay5+Sm0kCKraSiyNjLuO2p1fQPLvEeD3mfd4m/URhLtjAJjNPsfH/rCsU7DDIJg0
WIPWjEBjRN5CFBslRDBSBAXMLjGMtostkb3Z+3R/wtLYJh24bmB8beT+a5BpRwR3
dZ8y3Rk6wXsLQ5VPYoUNK9eAGBXNjAI5Qpp4mQCD548kUfhs6Z4IgCJ+h/d4U9KU
OI1EkGrLyaZVJZ6MEKysWheI6j/BV4tzsTWIThFIb48Q80uT1zG7KVg5+q7hySUl
htlp1UWnpcNvXaSqh8gCzoBlWNgiG4mhCwt+Zd8IAJRYjO3joVKit8WRzRycd8oB
bG2NhqIrZzaVoifVuKPxHWcfaaIpEu1+5mF8Y2AS85KjDaJcA+TNG0esoCTcXDCN
FlijjXRtsPuFAF+9yM8LAclCNp5iXeVw9Cm1tQh/3nZ0RHvUF7AVaN/BE/SWB4Zf
qYIjTNhDUq3gK3JSXjQIAycrYuk+2VaYL7KedpbjGFABTHN6Ga4ZIZ3isID3kqVu
8+5G5T1y2WVaDvmc8u+RS9p/ruvUy0RlnKuUPlc9cFQcDStLRYCXGG8QaVyqPTCh
0Qn0XLjq3LfRNAr0vHqsME2+HheNk8SO2VVxGs1IiuxIr5gEU532dFGGpUdVN/2x
IZATYurjzB1KPb0e6s5a9A4B9GSfuo2n7gmi1MFzS/d6VzntX7LszrqxIxDrJhjG
rORU0kAWuqwrRlwzenNkaLrNy8ICNtuR7OFVTDCPzs64qz0uGcpBn1C8ux2xk+yu
IXhhmb61RXRq/ATKC201djzOJHLUf9Mq21bPzjC6zA4jFxMZbEKWWPvkpqD2DqVN
YVOQM6k7jm4iU0cLt7tMcMvuYE4rCYCUuY6kr38XdTvDbXAV89FAkuNHODWFZIVu
82Z4LyCGkDn+Ye5z1c/FoodSefX8gYrsSDOQunDWOFL6UkeGmEig62qzXCWu0mU3
zjaSleWHf8sZk/a6bKDeHhdCIw/+wY+hFNRW7g5q/n/4laPuk1GV5OQS9modsYYR
hthzPlybGGnc4W1MeiW4T6lHcBAwHCRw4n9nGOdieDx1S8vO0D+9a4acfa/XFxDc
sL8iWEGUNlbksuaDxOFP7CEtMXZbFRPph0nVeONdv9emDiQfshndL2sdqf3Y7cpt
wVE5UbUMPWjFKuFw7aTddb9o+85CQFk+OMEZJDWlDDLa5VFyqKjWcbP243jxJITW
qbINVhx66cK84be9XgehHMlS6qnwhk1liECaQ7zKgCZWnR6UoKgsFghMsq5u24Rj
oLZakBe5CoGg95s5EunMX9qNNAbrp/oantzEDqxU6pp8nAv9o/tz4E7VF4YBm9rb
ME1BMEqj8D4Qa2Lo0Mhc4VtHnJVxaHWLq6+xlx6/5xp6zAsIQUDxebhgU3/N56X8
yVEPfctYoxIshpOA2ihJy1t6WYxY8QKjtLOMDxFwtZXdoZ63Jfcxwnb7mrwDTmWa
AzLt/Hxo8mbIBkvBvq8WnWhgZHfFmvbKD5TxeWynecsM5jK/rR5FguPVBvfY6AsG
6xk+SPSWwu5aduriqLosC5oWSq2O0ZDV0/80gmwoLpk20x75ffCAPzKKFM0eJ015
uM3+eGw/SWu/OC+fym8eGzTV0YoC3bZkjk83KMZI7iBSyqFeEsNh5uVC+i0/TQrh
6D8KUWOaTbS3Z3mr4gJbh5OSkERBnLSsRQdsXtrtTg8hBaUCY5UBinrZlYtO2ljF
w1IhpNzlgFGqJ8pgV0+WALwzS2T+QQsp9zYi3Em4kT8ZKP/RdyUScKgrBtsU/soG
5c29LmTMFPkQKyUpnm2M1/7kZ7D1p1W+7UPf00cbRt6Qm/Ya758/cHXwMe4fN+0O
MVJSDEdWG2phnpSyD1Pzn9nf1eJ1K/lng8aiDqlIPF/P4xB6kxqPBv9CYKm4jn0L
/TPB+YO00gso1I/IufWq42ApDcQb5L4lpSQfXf22b4FltwUeDfmNVmNz3+zLIi4r
Hqohx3EsHfz4VL3bEOz2njsLwaEx5vOkzhuKrHbEK+BGRM2rCzbI5t+YVsFs9E4f
21pxYxpssBI2luz+L6dnGBJoKyse0a5geKRLK6ZxM/lUxjOXxiuBMSh/UFK+oQd6
6xyG3TvfujKJNli5igIARw2hjpafXNzanv7pKxhAWB4fQ1AHopfz7HU519LCxcVO
sOg5udAgFYftfJSe9IcS8NdtGAB82XBFOuCT2BZwSkvrRWwzHdKJuB7TWYjQcV8C
WIF3FPvRTccppHtd229qc+grEtxzAV9MzDrejUC7DsLFQJvPK8uWT6Jmz6lC/aPx
IrjUCgtYTLR2LSU0FRd1uiUG7ArewCtMyZrFDfjhLbnjm/kEJg6Qe1MCiXhbm7o4
/SomP9OAVpoAiz3FthZGRL21jRpolEpvyhoRZF/X/ePC36cGHPUKXBzcU3Vb1M4G
788FTjunwaSsup5xK/PMw9tFwALwAYy0I194Jeh10G+I5+v3i10oKjwXMZrARYfe
YICM7yoNfeHSBq9PKRjnp9cHDif34F+G30TV5x3wBT41+5YZT7U7UnjiHwGWoocX
A+HFN6GLt5A0GlBybIU+i9DQhtULejU8E0MrKzWVpa0VGb/Nxp7yd5EbW05CNVE5
e3XbxjTj+NIZswc8KE5D4W5rvwl2LdFzfwg9QU3ZtMczfN5oOAPBSHdwnjY4rlU7
iuQPbuP3hgVNVluIAYXBDDQ7/Lnj8LkVnXqtHjFHYSVT2beZ27cjfwFyhYEpvlgE
4g9RF0AcxQVd0d+U9RUdZmPg0fDZalHp1Fft6PD2WDgL8L4LFlnwQWZqkMnw1+H8
0NHy3FJU4k9J0AGxCkBqEbRYsJ9lhT0nRdpKaNTudoOzSJnnY8MTXoZ3BwajFEtG
fCGdjdWnGG/rimBgnquw4uTBAHX5JM9zqxdwmKoPSKj29VOhEXWIb9NXxkjk4ory
fn/GjMePyUTCfN4UxQkJ2v5BgcFUTvw9N40UTw1VVCUNEzUneIm2GXFxkoNMHU4o
FYsPVGoin7fuK4NEEVleU3R2860r3YRHWIQZirdctnE0JzaQaO4HA1/aYuA9Hfk/
yIFG3kTAB85ShNfmYqpyIjNgByenJE59Ej0QfhLNsrFfhEN7a4Xmthdb6jyRBHps
jmGvk8pOAqRfUOvOnpCgAGhDFN769nE8PhIyKJ8o7B7UDkLuq5djC8/S3AdWo/bf
1kbAYbAiaw+QnqSxDEGcKjTplzqZN/Q6ZtZUEY1WIvsTNsDeGZrbxtiRByvKZJvT
IBrA5UsAji3TB2qNnMvZVDyL9B3EUAgqq6uR9lPYzthQfIhbiGGxbGdjJApnBy/g
YxKfnIqoxFertsEunnyLaSdSZ5PUwZdx6s+ev0VKDsFgtxjoxJOPNsQ1P62sTfNC
uWeQM35e9mSYFz/7KkOA9CKR885duENv45pJqZA5q4+ZE0gNgiQGlgwkrYqIg1nf
A14DnBvmZASicP14CxT0fVbMsdxH95hYss87Mj8GY7+6IQMp/cF+heDZnjBuFHgG
gh81vB8elBmDCe4LJrIJk5Z5D9Yf/vdlq3VukTdBnPzfeFPeqETGp6Em+S3CPLAg
Ehfbujne2FGr4Vf62kbZyT+NjGfljmi2XWl+tsu7BjAGPagU4AA1dYK9RVMcJQG3
Y+KbbxLd7PomItBU+8+7/TddLVbxECPC3liZvIArlZ65QX0ngE0H7l5Dts/2UicM
fBsqFHz6cBd8Ov0Z0Ygpuw==
`protect END_PROTECTED
