`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8zLYsmbDYXmMV7GbQ9M9OAdKtbFpiTUjp9Oy8plJ4vsHVUgAkIg09BNFeQnlSAK
rssJfGakN56DjfB2CSi2ikbG8L2QpKi3juV3GOAQSwVtI9ufvyRzfAVmMb7aEKHP
MuCgUKtS4lWRWQHWjuIZA3ePUyAUzIokWoLrJCqEeh14udksCTScMPm+zOkiP+2A
LTprqX88GqTL4e0WfWi8kGXvjg3HUJxwVBh2cppFpu/ftt0PmNLFzdIWeZ7w6+yr
SUc/gGDt60Z3yxQLg32/fglMnBLOIhWUXd+ptZ/Sb4VN15a3jWZYFu49GSFNSxtU
IpuuPEuWAqywEBREZR5Wbhurq+8OiEQupNfhMM4950AwVI9dRhH3slkMjwEV+G3B
zF1+erd+PzfxlqiN6gqPWOf0eQYJRcFHTE9oiiR6Ge0cb/OVSLEBNUH5hxRaXtIP
fKaES51kNuVDWixq5gOUGYQdLVzNBVZ45DHX0Wx79Wd6zzAtmoeQkkklSVp0NIAh
D4hUpXGYTjBqZR+9ThrNW2GyVaL0vSxeu393ZoUfICXWcyzd0J44pQLWtTqgL49L
usw4B90cC6difFEDYGC6QGnXoP5Ar9pL+fF9uD1DkxLKKEYgkJqJM1DXawdIoJTK
c+2vVDp9K7yHNtuhENKXNCq6BtQpqQkO56N5AOWJdUXThNyAaFTPNv1qgZvcUXNp
WaeV+5ieVsTLI/RKj4kJ1XDcf7OWNI+QqX8xk+56WQ8I+Ffxi00b+5Nn0+PWC6Md
WEfm94g7FAonWC8xYu9riWhAxhSl4IWdTKHmA4U+OPAUZhnDWuH6LYPRp02U0bdA
nT7Qby4Np7Srltq8P/JmYHc9/XSsGTR1sU8RdhXje47vlPDpylnyn8Gq4XsNj7Sj
UmVtW2yq4crxCWTk22lk68ieHq+dNIgjrS9f2dzcLhWIA1kx55qB3uOG98bkE6yP
1ymmPtY5htuWT1xtvlgw+XsBeRRWyjSLeBsMXrygCHYnjAa+gDACL4O9Phcsk24J
amyuRjMX2R5neNk3GwQ6sChc/cnfbA4JlZo2e+tdPaB2TbM2D/0W8DMfSPbT4FZk
GuHRfq5OLRV13JBsSRVqk3Xh4GeZhcFUZjhWx97fWjLDAuSqEClJ6U40Fl20FCym
IyTOt5J+/yUAOF2DSIeZbliRb7o0d/VZcdJlN7cZGfzoIIASW+vcYTDXg8mPHIJZ
Regk65WGf79+O7MdH6WXuwQUr/N5n4WtIqcTonEj+9nPbzRLEWOaqbleAgrU4DUj
dCHByumwP1dhAWjMe0rRvsgG+xph8V/HKrnjtWyFRa40ORhXFIxkqeapSDqNUMP3
QB5ra4EU4fAJ9B7rx6rl336Pl8uxq5uPU4y+xWiuSZ6DVWaKeY5o9MaQJNylY3zu
t9TPDqizW+tPRVa/kftV2ifLKuKVGjSiW50F+AT4pvknBxu6iPOxTl2i4qP4lZ/+
Nd9qZOrRKZOLMznjqTn/9koIWDlOMoLgWW/FwntSNOYyifkhUkyBOxXIe/xe3/5o
Eov9S2bql2gCtKCSjWFlxCfvGCC9hH594Rr47exHtDnBq0G98QwKqmzDY4Bo1wqL
gnPF8q6pZyv6l/ILtlUqJ2TqwH782oH8I2mVHaUxKpzbuinHvqmAetoW7qQo7np8
EVlCNn/Qc1UJibzFvvPPYuw5FWaqfP7jVA1sojOP3Hhf0OCPNCpF1YFKQA152lrA
+qbr/yF1x2TGXsKcypyTKuBnzs87cCpGILOhkwbXh0DQbUGGy8D0N4DjjQnveuDo
lbhZ6kB2j3I19VTp31dMI5E3zgCT6vm3PX/W7usvd0AY2wl91CCo7lRe2sv4BqZb
jovlu4y2KlhRB7RSS9CBh2S6RSP2RpqTt90W8TeUMRZSEraiuyd0SlSnIl3FCTkI
Tfa9vuZY1XnRW9t66Y3DAkmX8Ht8yrNmoZhPm1oYM5jhVPiw4LjB6NW5ZAC6m6KU
NfwsyBPipjZJ1JqPN1FZw4Iml1BBZWNWXcctX5rIJo1Spwb7DHrAZcwkUkSxrQ44
biTOrq58UjUcnTX0u6tWM5fIv1g9WCMb/7NPmgz7Sew38kQYdrOjTcJN2J1f+1Bp
8FGE7e7jsfcV3uLJqajNwhmTc7LDHUmb/iOyyZbQB9vgA5XuMKSu446kcg//kNIn
thE2EgtzIvktYvWbUHsUz459Lj4ACI1KKhHmo+d/nGsO2O7NMHNx5BTlr6U4RVgX
WsoMpsNr8dEBBjsubOP3Prh2Gau5/2eGVsJrfjrEYMLHXM3GMnDNLTI2hFZBG18Y
CWKkWXNRTzGE0ipUqlGrz4Gwi1q2BfCi3zgrfYqf1zxgiuP4pppe5ECp2CwKJkJW
YECDhYqN3l4STkjcoTcW75uc4q6rkFPQ5Y0/A/RhNeEgwGPcW2Lg7pvhJdPQBhFM
61XFYOFc5ScvPlJ+V5J9BesBhGET4waVkFyo7DShmFh43qujpmf+3jvGNeIjVD+J
PNq2rNKsi3ucnOezNUiGZGGM8WkhHXJjgYS5VWHo6eiqAzoRcEIHTmtqzwqoBM67
wmJkj+Id+BPXcNv+BFOHR3S0CiwX2kndVLk2jvAWz5zD6qVFAxdeBTJinREfJxPY
3oq80fg/44bhSTqpVYNCdfISH4qkon75ygvsCsvrvwQs91P9xXvEd52KnR7pkolN
KipWSKcvebHGG/EhU5ZjA659BUmVFtstC3u6gr184/icgnmoORDqWTqFs0SiZuhE
qgygd8RI4N5tkvw3G9UhGC7nymz7cxNq+OvC/REH8o3YnWb0WNUSBRaSFqhdsYLV
1pYR3AMSEQAmwcB7G39D2+gNS/jhLpPfbBnZmzpTzaZC09TkDjQ3KwigxpDLc6bY
wJMkJejvUOoBlEWqicx5Nnx4atovh4ka9IhJkGjBZkeeeQ1MwEljFbHgmAe4uZ1p
n6O54NxhoFUdekc+S16SSqnSyN1/AnKaVzD49LY6RppR649+PlGu/SZDR/nd2T3A
JkDty7ylY/3HUoWML4WugiTpWU0kKEBu0mym8VSzPsqc2qHso19RNSTh5V/7jOxa
fV+ge4T8ZH+uCQ3g6fP2QRRzU4wAta16jNDjAlYzSpvj8HhtzajL2OQo102jkasV
HpU0KUpG9DXmdN7fjnENKfx4dsgIS7PCCOdf8ofhup7q47sx2tXsIF5qAIuvZZ8R
14voPhe62ft/tjtIlGOuE0LmtG9Qmct9Yl9bR/2Uk9gg6KqbYZUZl2jEYiWMGhS3
FTWcDXi0bfheFygzt/7dryl8LRcfohwpVJZnqDKOOokNX+rxqEXWq/bVd7fu+nYD
yE8SKbnLxYoxL1Vo1xgogRBGcZUsa+yQDg3IzfZxbBUT/uInY5YLBgSCLh0kJOcV
zSSZkrDQu23DBgbO1f5hG7DDTQBZibzbm4yQtK2POIlXOGouBgqPK5mepIa2vSKh
6PV//QW93xcwtQQR4gC+QfSC6ckz6e+gXV1BaPdtto+Bay+YIj+jTHkqrC9R4WVn
VL3uTFqyl1QOZ7d6LYS7tSPQRLHlXt5yFJ/C2i3IbtmYHeOf5W1LMJzYpI+BtgC4
ncUq28emUaFc064CUsumXvU1IxKTFTVfMPLX/nqBP6+350Jt+lQOw+CI+TZpKtYl
4ma3v9ogsiuMLO0DkLbHmudLomgXuAkuMLDaGy/pOkyY4cYrs9SIDAw5WMCNfsQu
ILbqyaCXYfRHQP0OMHnuvfXRpWH7Ct0RgUC+ACTSPMbW0bxW7YWPV75JdcFoylZP
6ooTYUCnbCU74zGegMoR2tzjFRwcnKrcz+ADL0sUcR0fC3zhMzh5WXqPWx+0DljM
HKvOh2+GtrdgPys+9UQSibK/2nI1qvX6AWJmh8HhuvpFdyK1Fwe4N0anqp8c/qxY
E0HxT2pWMhGfVsd/l/LvHEjkQQ9Hy0a9hINHDKSHXt9jgHLktBfNx8YQRYoZwXod
I3QM/f3gEKeIfzQb+g7IDwbTFSr6kzjswyHW20QTDqX03MEvMU0WTRBBCnqOl5G/
pY/veVRlkBAugMzqxUAeYq248pcSIm7DzOYnmQI3Xux2dLqYYYkBaGZ2qn6Js3ya
LESCA6As8J8yvIdtHxpR5ejSj1xx4m8y5AhTPPbf98qxJsGbE7zuKf/C6QS+Z0KG
Lsee65wk55ilgXzso+WJmAV9FJ3a1uR7lcl5ZXa/5qvNi27Jxa1JZsjw83CY7aU0
BX2fC6Zva7/skqLCV22riDT9y+kq+mTsapRFAKHP1ZdSuNygwlUduT7CJ0JXowZN
VH13R0SXw0IApejoNrxllCeb0AHBf6kjYuhU4Mdo6T+IjrH/9E5puClWE2Id+uB2
OsZytpsXX/tLbaeqsYeW783alqq6zpn1/vRiDLG9YSW/rjng8hIa7jRplAZnKVJK
3n4ej7y2SLADfLDBrh6R9AuEzqLk/+mrNuh15cby0B64Hs9wSsdp65V96NGXe6si
NBfh95MvT7XQpUASmMBVioKlrUWm5Qg/B097Lc7gcEbwJ8P9t98GOL1TOrGEyxI5
7Gm11T/esz+TlkAOwZBNxH8Js/+TixwysGGXiN2h397/pWNIGFXwkAGnrDYU7SZA
kXwfIDkkU6jZraA2qGD1OO/mMtFKjZRdNFUegUya4i8LOeuA/jmeQcl8DhUV5WBe
NnuWs3o5bN6VRF9KxdLHM2B8qVUHsM3k6jwxmGjiVB4jIoVg6NGKODd7stYLeaaY
FKctbFtntSuedZ/Rem3z03U5eufxzhjCHhtxj/4b7JJPcTW8x0MG4xoVfwYpVpJT
YUqCuYiXnx54OZMBUaYKCYNuzAG4VT4QZHKlsesCBgpR5nb5/ejIwNzaMuAI5CK4
N9zR7JLwPEtAOJccXanMXq93u7FsAg7HthH5Pr57E5mS7bs/QGxX+6pSlZizW6FX
udaM6nVFEygNbLzh0TWvDwnwBGcyG9abd53sPcyS1xIz7OyeCgOU2zsmQqVCfO27
eSmuVyYXFHudPViF6ZnaFhKor3xhc/BM3DwHCeKfzSKKaiz+XAK68EGyT8/QAnTm
fWTuXWs8tFbLNo5Oksa+tmgIgYsNXg452PvZ4s56rM+VTdgqO+qlvcbq2PcODMXo
0WOUo8mA6Pw+q+U08fqLsf1g1FH+6qI8K90/HTgDrBbGDr4hqDTqPrp1py17NI5j
OvpgYaWkljAVVxPt9VMATGzK5bxsfMgTppBGP1EwtpbYjCz4JuYkOfm89XZt8drn
IUUvRKgqg4fRl+F+sb1LYAMv/2EzyFmX8+RavMtBquWUFxkQaQ1jZVMErFsraaR1
puGnIVqwY9p1DTomCllXe7SmVwMNSRJN09GG9vvPob4NZ9j6UAacslIdLccRIIbm
IjcFSX+5m8DRQNxToPA4/nnpPLC16y1BerYgPZjnvVqb5ydPtavE68rG1VYsN9ZK
KFKY1rEFJbnm/09I0z8juqP2ZpxEa3advJj4/x3oEJdAvY/ZPzAGOm8reNrtQZ18
V6YR9vnM9V6/jF0l7FYwu1nOQobn9DJQbwwZZvBV0YyUtgYbcIoZ8slXmGjOLZ5h
LxfModne6CvoHJhc7Cs2CMhC7Z/lKwd+OHPxwZ8CuRDICM2ruXo1uYBPl2mCjdRo
m6GXXGQ/llVIbEuJc3OJmrzY9pMYkIrrkJF1j5eHav70GIOJqKSGIlqZGF/0JiDX
WMlTqwb48xKt6CTGvQtRJiHZqIL1uPQVa+Ukkm9G+eh3m7ERUp4hC7lbuLmKL32G
t/fBeAJISkqOGdj9el9fuPG8AXziob57zpVfWBzHDucCxHHtSJY3CwyrYAb2nsJZ
48oYe8ABVy99M9FIKK/cVU3EuG6e2XF8nOec6q598wdMCnKz4H3njCCbShJCZ7sg
bdgECGhnJPqlKVkbokuRP3a7/boS1RuYi/fEh7/WpvXPzMyp/0GSHN+ADcoL5/lY
OpfAQm2pCXI0aQXUMmAJtKAmp39YmCWqNbAf2Jpwz2et2+W+EIBU9DyKjJ/b64zR
Np+66IzHgj4TTh0xer7CAKEJJL04I91X/NsIFC0D4RYxdpYK2OWHsDzZx0gkIaHm
Xhi/jexcmwZIHBm+G2MOfCTSfbdzfRjfI9TA8c87IlfOtrlhZwFb1cedDPZmufoj
hAravV00Bb6svLQfe4vsluxuTJB7rm7ppX8q2VmkCmYW4fibW1q7KNnH1GhyXa4D
u6Gq9uVxwU+ukCexFNSrZSsnYZ4vvVc8+Ygr7l8beC+ap0MkUWIbNElxCf5JzqOm
pqo9aV2zcMvxQtN5+VQD2aajTvPmYPbb2Yk59nU6Wu3m14eppBvnb+XeRqNJbRVh
4kiC10JZdo/V8IG2/+ArAVNkTlxpPTP7FxAIP9K1K8HoWb/DzHYkG9g+Zsh5QkKM
Pxq6mKRTETFUtzeKh3BW8VdkaC2E0i55LiLpBZAF9g2fgyGh0/+5BLG4PXydtYZt
uJS88s0blO8UrKPnAl2LbDjZYkQnCxQrag5jyYmAHAMQyeSqEJEwMXXWPZ3PlY/L
6/D5JEP0zQpICo3534uVqrSB+9dz0dWaXf3cuWN/Cld/m9mQVhcZ9L/rbF0GVMcy
nXgrJ4bi458agQDpYDP/ewe3/J6yB7ll1Is/9dMyFtxH9rudxD25ZVSh/wTVT7Uy
cHgzDjrmETHUvqaQShITRTCQkY+VCm5jihyZ1Vy2C/G2oA2Fp52V61ch0vSnPnZJ
tD7Q4Z6dENCAL8CL31MYvRPIZ5XfJanQyPhtJ5kEg7GeW8fmfHK/dclsvBcudplj
jtWDQohveFQ27MvNIWQhn5ypHnpdMx0OZA16jZF5Q+AwR0jfKnqpP9Wl4Qql3tcB
9hdZ1jITGlEAR47fizIBo7B+GzNso3dQ/HViUsl+dd3wb13aknmTDsKs+vrBmu/F
GkFQVAe1k7flC1H9Y4E/1+ctdkdTse2uNE7mI9PwEMbpYKuX56N45cvDXapRMBVm
tatK94yFFISy5SqPlqC4LWTlOzUGpAtYo4zxj/tLIka0oT5dMLQtvstqlgYDQiVA
imwYE+miFpo3tm2ZPsV1rkc3tf6JGZUHNM/AUmJuxOIlYWbf2/UFhFbr1eU+c+U/
ct3IroX77jLFHzJU/eW7fjzIsXPhFeP5j0L9uiuViSFsOJAEno+evMlFiAwE6oKE
hO5SFJkhe+G9TM6btD8lc7veTmCdzpW9gYLW8CCfVasN51haIQjCDZOcQ8WV4U2E
FfXs8usRl+20F86p6fKEa5uNwqClE68jE7WgoVrz3EGScwGvJL0mxAVcYLiR0kzD
eEyEEIgDDBR6LHhfnTMbA8/aSSkKq7WclNLDmI1f/zF8bZ40g1AXL7KD/yAGn0Ne
9ooFaW75Zhehmg3Gb0eLp+rLncwQlcz0kxw7qFeU8sTEIMr+ezjD/OVREucTbCqK
PSeBKAIYA4UPEgcHoLH/hOFCUzRmQRqIuW8h/WC8rnqPa9qvwRsEGuWGHjEE/Ybd
hQgkWxAxkTXrpSrMYF+CGrU0k1HiREYG3gxKepMrevorU6qqYgYiep1BdHBclCpL
BkjzjeL5IX/8bueUlXvQqp8ou0sWhQ+DBwGh9OWRwE9Cjk+JraOgsdCUBDWxXNHT
ZG4kbdQPkO0Hjd2/pTffs/NBGMVSjpullGajjzvzMHYdi1IDRr1wx655ryD5SUhl
Q/0PqyemqMH6enHLrLi7X9B73KL5TlGpIv8e4JJsaaToBJ2goBUOtKj0cEy+mMzy
uq8tv5hkkqUEQlLDlbGaO5UmeahVY6uNUVz6P40H5QAxnDcYpsGUXVIwlzS8DJcN
LXaBe+ZztWMR03Y92TYyUvLLEDZuXNUYo+60lxvQbsirlO0DITp5qWnrJkEqqTIN
sUo8w2won47jreV6cy0WNAyRriDq7OyAiSIf7/oW13eojUJL5TcvA/YWTVTcwCi3
WpsxQMZWnm26GD2wijYPoHfuMt7cZRCBp/dbhrTVD/8au/1+NB+UufQ/u9gadtJr
S51NQWpq3T4ttVUyye6RAAzIdnPq9WhAMfIM060dtGPC+JqsINm45Xyd/dpN2mvO
hU69jlkVOSNgMBUsOKX1GMG5UcqxcgFlbhqHmQfb+Mz4aubrpFdOO3GqVX+NBgiw
ErUr1dxQ4nvOBIyWm9mD24ocp4nfMTsl6dOrAOOq+0xhIMKqKdDwbhOgaJVrxwOg
1nPW+7CT1C4skpCIvPqgMmZQdHkGviuHldqNEKA4CjlV3z4cHJxZL72bZV6jJFv+
kv9ydr2TinVXUc/XVeXdE0RA/cD6SqPi7MzGgZM/4aGKYtLFZebG9d3biSElqYKH
FO+58mBW5Frg4d/5QSXjvEzwVDGmY8JhbFenl5Jx/KcSWbCYixBUn0Xutjob0s1x
inFy8honNB5g3snBIcHaPrDpbj6v4lTuQvyBsOWTLgh1y45lu03vnxywHiLOX8Y1
BSJiErI3hMrYuwsnvdCa117Khk9q2aJrwRgwnzvWSGCenOT6vRGfJdboiUYcM/Rs
O6IIIpZSs1gkKNxig6va2l84rGPW3t6c0i4Si29ZkvnVF47OhYUAxa8UaFY3QYIk
NCOlbBQUmyWlKm2iXu2Mg/sLdYJXez6Bu1DcPLajXLE9HcN64St9g6qv00009Of8
NkUt/vVCpoa71sl5I9Ehnti00arkCTW3OVSYoOrVt9e+L41g+rgEddc/p9f5OB7s
fMGIfZZvZTJRvAu3JoBUCsnNlAQpJwftxkfv68QHikc+5OwfQyRf5Ne8rO3LtckT
IXQPnjgrEIj8t+oFRuf/iKGlikr+hfMNtRC/rl++XNHMDBzddmetsk/jrhJVNODH
r3m5N0b68BQ9PSHwmrZgU/pXPXXx7F9+lZcTrQwAIBkwlOUlzWB0j4Ms401cLU43
54aiSrS0H+alD0eGlieLm8Lzt4A6+4nDA5hYDOQNgWtUpJgG7lzbhq+WobDH07Qg
6sR1FPPSzS/fSQgrovVmlOVgL+8+XjAofM4ZS06jOCJemkfx7CRIdvGhmNLx75d8
AOTuS5bXnxRlrYpR0GM7k9bDkn+lx05cC0esUTocAMqyvBzbRCaV9CX0+IZja5hO
b3XRDRgH/x8UaXS2Usy8bPgh9nMeHTNSMB/WEpfsNg4y2ndZPPULMOntJ8HMRkLW
3jCmYTy2J4DKErPrltUr9rJ6KsnR+kZsdh4jewGf1DEGrL1WvJZ3QEB/SVqUUg7w
xSixzdzYGjQK2MJRui8jd5omAmcNitsh6LO2wU0ZwkS/Is+qEP1uYB5FlS90ViA0
ov/CatPK71qHC2YMHI1fs6F1gnmLOGQ6hFAD3hyUICjPtKyXcg4L859x/aaPv7my
11U689eEbC4IC2ZzHe3JxTDj2+ca3x/Gbjh9E922S7tXfHdlHxASYl1uGd2QjrBB
LF2lwOJ3Pd2YiKmQXa4uwLeDS3l3pfO88iy6Q1Vp0aenegylwWSophhTD/AwSH7F
9sWBpNn7ksK7FVoSgFfgahrxtrI7AQU7wMhs2zTxl1q+CwuTt0kO6VmDEcNj/RwM
4oAcdBvqEMwnqlCnE3Jr+aFhNlktft3XDifunNbV5WAVR5YvWTHrUy5SUhY8Vfdz
mhkq3+fdiuLsQjDvlGHeGxEfP2YteiDLt99vmmYrlv+o/+tU/ASkD6zp3BlTD2hd
Rc4jTllNzpnuGgejW5TOtUJv9Iw8io6NKft426XwMwZoWdnHc1QLiwVRbyg4V2sm
l8TcviL3hXB2hMxN1eMvFSRsCEov6tKziXgpLsG/yDrOvqUGZdYkjAGbRE8SiMUE
TkPTGOQoX5B9pN3eoMiYqPxC9t/CarF+IDVjPbfhta2WYRNqpWwypduxm0eT9Lzz
xqdoc4KCgu7CwDYq0XdUvPNoIcvdzFo4jdWYozmrUB08jSbH8+me6BiugZ9w1KTz
WbZ1rg4AKZNyI3B+RnnazwBpCUa2ITCdWA5HILMbYrgA5Ey4YDCLEogJPWbxVK5w
5KH2glKijNivTQxnKRXROKbOoh9IUSOVPkXPUd4SeSRm6McO9A6to0/V7uFDAO/Y
2I8T31sPfZd5PfHpb+MjSQDrcgWPvzmCyCjFpn6eqLx40QnetOM3m4PY/92sA/jN
qNwTnvK58sRbK4SAi1IEGpXUVW6T72KBdfv0bcKR5QozHxyWybxCO4Sn2NKQQEUj
IdId7m/g6lkIrdGQlF8tlrn8GDTTQrU963J8Yook2g2L9WoSfEtbfgtwLgeHmuQg
avDVIH9Sd3Vf902c8ONWUCDBMnlilqqyqSrbTksgSnATPXFFCd9dcbBvLbW9LOrP
UrVxmR6c8NDEVEmu07Xi96/WejFnqyBdBT1mJ2yiLB8ySsP0+rn0cRXzbA7awdil
v5LdPrdczWXy1c0aRJdodfbRiY3P1Qf5QB1g4EvutO9Q7oRFhgpU2n2gy0WqZ0Lf
SlifSbz8vSSJ/+ZTsmbUsTVpPPTskuVXhBXuGnKne+67LJ7Kxecr58mspXjeUePo
dRf2ClagPCFZqIFmKH3afs6yH99AvRhDNdaLxMEMIc34am7wmq8/0JfC+QZOAUP2
rKa/yGlPibHXdfk6Tl7Uhnh2sGu7O2duCa3PlFPhrwJr8c+lG5t5v8zvgmPN8O18
IJbgj8tSGSL2clpiqENKAkFnzBf3vRkQRd5+cfpvVyxyks/uJ+HD26CDyHSIn1Ar
nOkWf+2uXW8Pw5DvbxbOiVe3MKFcD3DCfr4NX0Iz9v1OZhkgD1o8+SEwVyJm/dvk
ybG8oBXg0Wivkx7Ds/iXYL2LlWII2DsdOVz67rTGt3inNcZP1sLY9U1BZOk9o2xe
jgcqjBx2xys2Uy6sKZloPFk9QG9c0eKvgLgBvTQaB0c6IGy7p4cy8LTbIQOEUShb
vcLIYt5u+wpkObHwyANoF/xCmzFMNjN02aW54eIWieGONbYqNj0Xtq7NYCKF5iYl
DLBQCck6NW+kRRVaj6kuGUKGeWmXmZtICkvHVhM4oj0RbQKEt3KUpBf1G6UD1PV1
oMBlPXBZ4wlx91vgtq17uz1jdmNn2uaymPiWC3x+FJNh6fdC8vPVH5gPs/58TSme
pWqsGDxzUmDRUZhuy5IRF0zh38U6tDRbLs2DDAxWJU3wX/lT7cdsOgUlxDagAvyc
4HR3HJO3/CmtNF6Y6HaPlyiafsQXjECC/Zl4ohLJvxEQT2t88Cs5xILc6wN9qLPa
207M/Tqch7TDO8GE8r7hJ0A/0F/npfEhTUQ4b9tjRePtoTXj2fF0jiFOcQORevRM
UFfl8EzE8DIjeWNQlQTpxoqEofCZ+OnRjzJ/sbsg0QXUpqFpNzZtL8LsA6TcifYP
OqhDxX6j3B0XhRSNfEsJ7pOK0dOqSEqhbOgUgGddBn294VPN9ceoL4GyJ30CxTyE
UUSS/nu/bGc/5yLuKiiVCawuQXRRr9Fn4Cs5yug7fnt1zRegRUl2YH868SyxgiH4
swlwIObNCMdWD57sCuZImJKcHss3T+qi/HnCz82enN7NDV77XiIXSIK+Hy00PGNQ
URBpMZPSs4wMWY2B+fiLv3AeAEIMKC8t7fOc8+Y6bUAooameijnXytmtjYe1msJR
i8yxOM1OAu4JyQNxKFgb4GDpUqr5xZ9cpZ213XSS28vNJikRUwGYbcvr759NJ/Ur
WcYaMfx4svPl/3KT7cp3vOdKddP3JE34ayVPpZN57cQbtOyu6JUj/v9tIh/KZuPI
JQbXUe1ZKOduOnLMd4xVpMGrip1MNEEWDsycnKYn6XVwYcFUzUqzA9rO7V2XlzTn
EViROa3PAPS3r3m0XuZnLRybjvwOueSd79aZiqNVbG8ecrnv+ZkXYyt04agUtc0h
oBKjJ2+dtGKXwTuaYeFd+FIfw9eKI0Yl2ypw8fZXHMuFCtRhlOiOHvJGYIGxF/PF
htadnU4CUy8u2Nddrl3vFZ778zZlIXv0++I1e4+JatD4HsGF8jjwxQxJdnZz+bBU
1XjmgzhdY3ycxSTayHj48OA5UxRihmSmkHH5bV3jzPgaemczRvEh2F9gSUbiFDms
+OUzx4vc43qd0A9PIRKmA/PmGt1M0IINXXakH0rzM+RbrNFcyjnYdqJLpvTLoGwi
9HPybZ1qDqwXiv1aNtpYwmtF84lhmd9/1E78TUnj2Vi4+qteIajtRSKzyuBoXfb5
g06UshL2B0xxCdJ2VQT5WI0QhbD33BnMvu6hp4vDBa0JSXkvUkcMoEgmuCxBY4Uq
LdedN8gyWxnhbNdcpdmzBP0S7D+nLtIMycbAuCjTDN5vOgUJlVkkEJprc2c02G9g
FrRFI/+rme0uIpb/i6FUvCYSSJdWP1KJFXorlLYQ9U6JnEc3qBE6OBOy8Gs51IcE
Evd3xvWk+EumKbP6H2KKMZPW22GMrACP3cfti6IgOacVkJocQyspLqsc+E43y43Y
Ct5VQJzf2a5dWGJ1iwoO53Kq+isn6x1zgQ9biS2QNayOybAtOzTeeFRIzR0Rjtd2
UJuNLr/OfaTUk5rh99C5Dwl1ofxSUzHHTzExg42ZCPE8p1SYraygVIe6e61jLBBu
aGKUaZ+qTAdsDy3w1+hgov1yIU4kwfGEt+gMuyD5qEeCS0iH5pMdeNHXPLw+EJd2
lX0alSs1m7wrHLIpUWWaw1Gu6l8ck/Lafr04Z49APVRQrRKXbc9ejFbYJPQDcVIm
Kg6bwr61hi5JT/bdmliLsGRXMiYVfwwpf9ghG+RPXMuZFlR/9ocCj/T9G8kX22PW
nYYwIyF0iQXOdKIjMHW0NE5pJRLrgxk54ruT3eltXvwhwcW835wSJbGB5axH8P0B
F+EXG3M/zkli61IOgaKXfxAkI4fFkGkCyufBz9lhm4Nr6QdHkabYkmG/J7PA4K3p
zGAaFL/17WZvk0NoGjeITGMTYSbwEtwtR9P0RPjuuQjVsWo12IIzWYTNHHKXLLGN
OE/jggDsWR038S+BalnhvEmoEN3O6s8GLBB8XzEB6uspfR3vKyzA9HJlUbdPvIWp
ktX1zSOPQKwz502bVzNffJkzijnVVCLHqy/SGGFUq5sozBfhMC6m4DJcT0pXGQzk
USwXOiLPQrUgOQhedbqAqVinTAtVe6dzaqM+Pn6j/xApH3OdPdu2hioJ1amHSDCJ
YXUzfN8pSHjbCD4RXVOfNk5gkiPPGOHgKoCE9twmMuvc3chl66rPhXEynaFZvKkl
XXpoT1WiGLc1HlKS0eZtKlFGrF43Mf4Apu9DDkVE+iGzAFrjZNKDnN1SRh8uTtK6
3008myeWfo1sPbg+uFVecMQG3cVAQc/mX19eTkf3HstJGHr4jsGneaQKkU9dCv6B
4pGq1Jysm09z2AZRTRhye4lM4rbM1iyiqn3SLS43wx7kjZXPQToPexnH/eXKf/Jc
VF1F/kDA1zT8gxFCuGA8Pl3R6E8UgIkfZvSpmpTvTT9Mj2F+OgTcDRH1gnkFAB+h
KSlqpygVjEUqNq4Rehp3NDUd4hZhBc/Ykahl8TRIIFl384ofDrUg4PEnswabenPO
2I0rTiqDhKDkf4sKhjEPLOIPMeAbPSuqRPXSRgF1PySwqPYufgWMGQ0vG0T0u2NY
Kmb7Oqa7LNX6+qZ1DC1HnRBjr1yZpYp3TEQIGmW+1DcmBDxI4dOgkFVMujU/NmC1
J5faXF7/6hol/ZTtvt5nZ4Q0kmWxvi9xsUG1hfq5vCmKDPjCi5iz5KEy+VJVrQc8
8+lYCLWn5TajnM9wDqC9hSPE7LW+nK0FxANwkAzaQuRGkq9Cm0fhDBnulmkW0a5I
z4AApR7R9n9UYB0dw8umTZa8TYAvDGnbFrT0mtPYHIc6rmgXhieEhB9zxttdIlan
CHi1R0daik5jnv0i18VY6Vg6WvwFv7j+zHbHAmN5oR8Km9kojX+KbHIIcfyLUUQC
vlXVksXfuTJTC+WAOR5Os0KFGRvHsH8KuNFZAyyXEx/MPWqHxoSDQB5Zy1qD+Xl4
/chxhT6LsT4cNZYeN/JirOF7qide4I/CU0iIky37bVZk4UifeAyABTaYxvteB7XW
TXS8773Ook4RR1ogeD3HRyRSLw5E/5sbTIjXg2lOfc/Y4DepJ5jbrwvtGpl2N0zC
jKd9twZ1n4eTsWL9XitVHONHTocJKTWg0JJx3DgByCvyLDN5w2d9mjXLf1EkNRRW
a1dUDwdDghtBUrUWYNnyYI+DWeHwGQw9O7ppMTMlGQOgkKy7p/g0/OhqBPQYR542
92UyesXYuNGCQ/i3WkLuYIUsLk8qy5OB1FmyULWZ3b9NsAcapVhoSlY9LJaEYLX8
e9C33pLv6ni6Crv30gW/9yQF+nuQk5DTkMlGxPSOQXFFVXl/wTypXjXLVIuKOIKH
+dB4jGfKOTfiiqxUT4vbb+KZpHPMJxGym+2aZcdSIREI4AMN6u3KZ6GnUc7Ndl/B
Zt+3xF61r6351QzGx9Y7KbP4WO85dXGMJ1QjPeA97pb4w4jTmqj3O0/o63QJdGk7
ztpaJY8DlkV9tFZz8zeB7IfL2gOH6Fwqm14gHJwI3Y4iF68vabL1jEdIKWdI684e
qcSTg/FV7j3CNc68zp2vJw3Xb0RDM5XsIbp91KVRVfigfwp4pGIhZJ5+p/y6Rl2v
7KcnhKwqDGU4SfOXYeeralWfRjexxpZUnt/0qDw/Lqt6RDhvSYeOxTdUJ1mvL5Od
fR8WyWd3Q+WhSnoc0upKz8V3ncSDECRwEZRGk8VXnoqEkqorJ4fEuMLrO4dpV4pD
RaXIULHRuFruRTLGLB+xSmwMKz7TRk1P9urf+/u6TUUIPITS24gXM/NypgReAR2W
4NNV2c1VDNYOdnbGuGtY1gYEgVkAeAzOjFUF5sIQ61himSy20BkJqLMcire3BQU+
d+xx95QywNuigcD9J+TauPvjII6HnSiNHGXKx2NHD5BXziO6Qmrty9ju4emJjP81
LsTfzyFtDv77kZ/nXMjlepULdK9bA6LkvN5Jm+PYvJy8/u25UnOyiG3mESRiHWjJ
l9RAsGKmAVs2o8+OXkSRt7S4zJSig/X4Lk+Hz8+MSF+nEblqevq14AMJOa8hF4PP
QUH3+8R5NB9hv3I041EavrOodmCo2+EJD4mFSWrNt480DoA3m8BppgS5jQHEtofm
0xXQHazYUrvpm/6/hhpVqB8bX3AITKBhIltz9wDDOWu6kx9lNKqoBfY3GqNwPh22
Fy1DQ9JzcDa7JIjEvVuEnClLaMg8JBk0mw/KkS3CQtPd2rTCb33jL3TyJY4CmXrB
NZgSudgjcEYVZ+zawYgfOh6LvNSlhOcyDw8aZF98xykbRYv/whU3fAtVgKQPHPrL
mTG3pYDUcr/z+LDtb2pgm2nur9cCnK1/VF4CGdUpz7LvMjfXqxyMUL/fAVgXxGzd
nlF2MP+HVdOHRrHq6kQDwb7WZuToaQ3fmpExQbrM0cOzWsjyDv1Po+18SLuTbsN5
CDjY55WyG3DAanscPa56f6YJhty4jPiuoHeZfEk5WvAid2dMYk+7Fgls2oNzlsnC
nqa5Eg57rrrj71SHHJfeidfnXVg/h6ajmmvodpuQ0ZhpB6D/HuiNJiiUKQq1bzzt
O7VqHAhuJJglIQlgmljPiFGAPbajE+FkWf+RNqLUfR19hGbelZMIzt71o/jjDqvF
u8aD07MtMj2lie273jnYp2re9mog17weLeWbQO5FhD63nY9Mv9dXVzrt3u81EUxx
jxXBeOpN8JFfpR1jkgXqcev1i4PKTkJhM15MVTk9Z3yIIuyenh+PHSFCpRKKqbnb
VsHsK1SEAoE8wD6gIe4sEn5wUZ64UQcYR2xUiGLZKmBIJYeNCCq34AwnqNajXbZs
xi01wAf422aJGTrflc2QrEgr4eG6s9BxAccvrnfpGyn1wGNdJeqKblyDunrk4JDH
ZL7SSaGf3MiuAELDsyUpTx38i0xpmQhgNLclcBO3GJMtTQWWfGXCz5fsWu80vJZh
r6ZoU9NEAMIlBE9uW/PqENSNPa9y7hEWOt3fuQ0sAMf3GqjF7rN4CAhiat1N9+5j
a7xXVcPop2QX+yFNDgjVKO+3LxJT3T2Fquogf9K09xS1jMbTTteln6XaZIZz19Ta
kPYTJRzVnIF32iK9n+EyoPFlE0G3e5p2D/deXW3Vu5x6nWy24odN8WlZkRi0ixE/
VyS0LUSZIwF8KGy+0iohBcDJNEmWRhqb/Cz9SsWHvchHEVVGTT95DRyRADHukaTw
9MLwESOmJ3ILuRmv93Ar7i/Wtk+Hliu2ldhcyFSrKUQK8RpFLcvBrktwxNi1YXGN
7v2uA4kiimwA6IMuUfbBontIb7stEYq9sNrdPsePEtzr4FJuyVsVBvVS2vM+Raw/
uyq0ASjjT23m69P0KStLfQsoUNfTcENJ/fDOgOTo/15i7ATWcYNgKXM2mDXzt33d
5aoPNuhFC3zRndvyOoFquUKNVUwJPdyFI/49kEfN+ZvpljbjxykYXPDe3djMS2yf
4rTErmqPc2fm+IjrJCGxtHs+hnJ1D3TcA+XaYUXsTGR+uCkdvGjwxoUwxlLxQA2u
Ej1LJr0MVsZx14FraZ8Ix8u/V4qXZiHtb1JE50wcJV4PH17jDlEUWyhjKuwvZiPa
I/xbq3zzjehql19lJEh+LkViuvNcbHS0rCdpL/5SyCz78rPTdB8hzbAlZG/dGtvo
BVwCm/tZZsUS5I9yR6bMnegRGtKmRDTT9Fs1+C//5k3zlV95cXSpxTfSdIVjqxGf
4rlv0C7LCe1DkWk+DdvQ4HJyn1E+XVCDuoLA/0Oi7NDTbncj1gJ5pdLucXg/j4SU
JNvMZpdQl/xNANmbDUCE7Hq+X0y7ZN06MQZta2FSIjYvB8IVb88IZJJujycLa9dj
qIpPYKATRQaZYd3rn2BCgAuYcuSCoZWOHaGbk/LQ8FfWAzKaaColI0jSBPvduL+n
p3O5+UWHxEJEaxdrKzCkkR4GXcVl8Uvo3FYLZ7mm8sL/tiPYj7Gk6tWiuZ+x07/d
k1vdmcBc8p5jQQ/oH9u5CPKhXkSn56T83PhYjs0AKdtIvA3iegLSCFTnHbBpyANY
KA7IhqtMsJ6EVwe+Mh4R+tu0MiyQY/YsCEtt6byzDuON/e48333AkrMrWc0nXLPr
7TZfyhfgq7s1gCMP0WQ3v4gODZr4MH78VIECEYETjDLL3iwPJA8pOIApIz6ySqxF
gm1rXvBCvEP679hVCqwgUcGvFYEVHiZlNZ/xeNOZ+Rin5MhRbQ1kUkxn5VQ1YW3A
RyPuMNXcqCxb5bO24p/z1699+sfxJgC86aWzUp/aU23vUlGQgnn/k36QgMbDDpoS
eQI4JRyd5m1Pm0YCLNUauWLJ8Cj2RNspLHoo7sYRcdfUKW07XrS4f7B61w2a4df8
wA58Zbn0JMrfKE1334BSS+pP96mvDV7DtOdCi17vjXVYo+6SdDqEtuTBjReH9nIR
QE8r+EGInCmkVaJc3wKCaVYbK+f6TFQM2YXxyuV3AYZft1gwe1vqNjlb6FU8d5L/
Toh27kqQnM+FdELnnJEBAumwqiamBL+Id6jLfXdar9RERPQw0yznYkrQxdIR2x5M
mWvpzP7/xAz4HKshI/51IDY1+KVhjGmKY9E0uWESKZ6JLA3OV06HzPtrMvLSOJyC
CkJBa1HijtnilFo2zHUE6zchdqb7tjZfNcdo7xhxmsiP2rKT1G4zRoVNzRmA2MzP
kFdIY0LVx9bS6O55fOk4rv+xCLHyuXatLehMtIf3wU0zI1ez0pTaZKc3gktkEENO
QK7QC8iKPdM3s+3JyUvdU+UvrP3+BxzcTeGQNP5NMuJje69oO64jb/An3WCyJ7M1
LNyBrOK4bypiWvhB3IhRegQCc7x7OyWgGPfYcpFhe7zxGgbfEsW8HBQh/7HS2f7u
rZ6gdqsURcfNtyjpweZeqlV03WYaWedgDfFKOjmcU86/EH2XOfuzXT1+3s6SV8cM
zNFhZdP4HNe00QPCUT5E4uXtkHxomkw4HoDpS+l96VOTo3qK8OVPLgtISHX8VfpS
D89RaeEbXbXQMQjGTsIPzvHkANvQcD4aPNGwann2a2zbyQVJujCC8gvF3HkdaL4k
3l+SxrnmrJJcTgL0t9Px0vgBsejqTTyTV9zNHDxdS2ntJnw4FGzpeodRLjVc5N0s
/RdZQtTHFEAk8G/tNxRCHXfNWAeK06TvuvWD64uKiWpO08P2NDQA23qkv5HXPTrg
cVQc4FZNXGdRHqhtTkY9Hz0Qt5T4TSPgsy2KmW+LxbqCI5iNae7tfWrD8uhU7gv/
mdTRJhmBIgq+3s/tTopagll6/q+pWQbIV+AbkSCy9PPzi0Tmoc+3Uw8x2nejhm0u
+AP24OEXLK1gFLIimVTgVJ0AVjn3Ol4ItPFtngeu81apc9P8CNlEvASDDOX+PLay
2gBejxg/s33wxG5EF5sR/j0nmEvMTDwv9RvcdXqXocfEWBQD6N79bGPYr/fdRJox
UwUla9wdXg+G6cPySU6FpgVQ5HOqBiK5Vq6T1gpMulp8YOzeOt4L/cRcv5iX3geG
uQ5DmWucbBzmy+TETfNc+/ahR8YFqkVFwLJRBzL+8FnEjIyjckSBVJC48dAkB7YG
+tfwmctv57LwrySqTDx5cCc3WmxH7+QmXVSC/9gT5rzl/cLgWMdB0mioDwNFRlNS
FrHHBLd+5q+006h5FEWOsCCqOe4D5gxV+ge80I0NEwDw17ndiwctunyCcQI+Nida
+w6/mfLyrm18OAdZD6nXLGhieQhJ+9oNBMWtxGIDOFTXKfEBvnvJ1OmIci/BsDqH
TufnMaqAP2PEgSyGCgxEfTWoCXLMEf+pMSzGhckpRx0gDJHk4cEmodQ1NvosvCc8
s8HWRq6m2yPygAkZI6G274uAVRZO7SiCWcMRzVu8zY53tqiYrjlTeR/yrxgJp5xm
bBQepjN83Jy7Kk6KEz6XEXrPSU8XyUr6fALNDyefuPv2Y/eWV1ecaauF2NuQx/WB
rCb0YMhoM0FovfD1O1wel3nI3srPN0QE457oVl27BQ4aX2GRpUbpalWRTDVJDQ8Q
xDf8vVkM7OrJ/xkvdGpjbeanXkk9qInYDfrln1Jitcou8+7mG1sVeX+6iFA4RIEf
oFJ7LBw2h0+ZH2J1D/E32i2KFclVhsmDrHIcNB0AXNpUb5tMKu3k1BykChUJsLb6
H0rc1tF4OsvjCAqICzA5wQ+zx9BzmL4kSARD85S01CUYzONKcFgok5tEqaFahIm4
8ulmnhVF8JQv1/Sf4NT8qePm6iL7dgjcif7tiwyWXH+yu4sbpGQ3yUeedFFU6RBy
UPYoWZ43UZov0er2mZdZhXIirGoY1iQIW+JYwZOT+OjaHeOJgcYRa45tUN+8fwJf
ocoq6CH5xrkvekCCSlQ4Pd5ZxeXefFU044YsSdNVC1wtIYCjDQuzlvBSZf4RRF1u
pOb8PAL/AXmEZWoMTFOYsWqSPBSM9WYtAFk4LSgS45KgI1CwS66Ppg81ZtAPQx6l
wfHrCrPnmt11ZbgLFfL6VF8fJ9fWZFFwg+iuUkrw0e6oMurBotYsznAiylkQMdZG
OmXfcNOupQAXiuwtS1GY5Lah5TKmmz7v2hjwaLgykm4Zbd/Mo63sP3Ko9I32W/dx
qtLC+jSJzQImgXPNaYs7VfO0ByBP6D5QVa9qeEr5IKbR+R7EA7ERVQokYsV36kt2
nwam85AOhwii3rj1og5S5jUZV+8RSLmeARpO0W4mkT6nfZ2mMst6Cr48GCXMv3ph
cvN21kfSCe4GeOnkDykvu4I+svzIZ58Ap9BSR5xE6zPG0epUN72LPZMND2EnUSQS
BcflBwkp39ftoC3vfcxyeMLYhCcBfvscnuuVhMl/K5P637VSZGlX86OETtJRjg05
OCe5mZd+MjCVOl4XqAabjmFj4Goly2G4gcYsTHfErrq+X8ZuYoIUXwjuOPO7bcSX
/4g5mYIsWmrpiLijWTgX8j/Tcq+gftr8RLjPRzsJvab6A6yvSejImeebSwMDVEMm
39nRJ0RICX85aJ7Idgqc27s64FPBRkTKKy2MQEvbYgBM4Hnwmf2CS1HuLs08FOGg
ORnZs50s5HMmrRhuctmJPzNNIxvRK9UEl8rktd2khnmeAeLv/wUK5dJCOg3/NXID
H+pblm1BTOl/PaXgXo+ZDpZbcyoQl2/IaVt5KrW7syVgsJpXmplx0NARYt77j3Cs
uaG1PA0NI7abozamgttLGVgFjTzeNYoTKE7grJKEzSxfZukbLMIyC6M7IT1KJa69
JffPAiYAIITcOu4Z4tBoO78ZkSnVmsFH7uICh+c6m8nU1/vCE0Sq/57mt+Hpj8CX
kP8iTxY596z8vvPx97D3+GpTO6zo1B19a9Rrk0c9m5kwUmGWQZr9PcRLC8H/URkj
CS3MT8C3KPjUjif+AinD1kfW7nNUVMBOnYoaW7fDw8rzVRL4iDclDmqyMMCr7k1w
WRfGhQ1wusgFyvHT18fGjTLlUYfy8fsheJhd6QGHoADmx3bRAFuMDJZllAtC2kj0
pyK1ZtMG9TI00BUDsKVisdJcc0u343l+uPVN9EEl3KQs8PxmHbvf6i+Osld9BtMl
HcPpIBzFKAhzPB4vzRKmjLqVGt21d9AHJxvl6V2qtw6joDNgpKNfZRqHmhi/X+qh
6j/Ep2Dg5k6a6nlrbSafxlQKjM80Zb+8XUvr7qqYZe7JjUE3iWHVNieMk7v+mqmW
EZN56ukfcfwyV+pbFaNRGISrsoCEpRssytXMYXVoVj+dJ6owog4+FHyJmtg9Et6P
Y4EF05axd2t79HURckXynHqjNE456sZO2gprZBCoIenM8SwXQna8/5hUcQwiz+Tg
qBR34lDqcpRMEDZ5gA1kVVSQvSLFlzhZ6R5qfomufaBCo/Jtskt6kU+2yOcs2Z4b
E4LTvEYTNZBw3/yh/Pm3BQXw+62BTFiMHMObnqijRQHfehCr364hJAbJN+Jxq3WJ
OCSgTxbp3ZGj8CDYRLR8YZgBPgjWaBxkxiiSA5BXc5o9MEV8wH685xa1j4y2t6yc
4XiSEogo0vdkDmx7kVxzrATBBIaSNvouyUMVTmq2LIZhNTBP+kjwoQ57/LUpIJNa
MUqwn3YpdTdPpSqHtT8sKoRFUQV92UDEJF6yfeNFVhEv9qetaUWJDYLDB27IKK3W
/cg4s6CON9dQXuSi28mGmrRyumiGVO7BEHxNw3vj6aA0SYQ9UeWLDqlC7zTYGiwF
ru0NoGXhm1iftwmmTY3Uy4+yD595scxoebQuV2KlyjFZEEBnBmBag44zanYvDN28
c1xPzmYy+Z9yE0nWTat2VHemE/Ur7gDUgXOc6ooZlDTOhFUW0kuBoo7qDfIkAZdm
ec4I8QVdNxZh/V7VuAIDnXHr3KmRmkqnFQM0EGMXaoVgFdUsKpCA8wPNx4U2B9LR
h6uPqLyMk/K1YcTSVyA589YhZFsMRJ3AziDgBMgVD7xBAqqXDpY11Vo6nS/ySxIQ
t/Px72gw7Sv5OP3XkFA9AvW6xyIcI5MiuvHfF5uThRDdhNoH6VrDylH+Gmsnxd/J
VZ8ourWHPLygVdwTu5gPQ5ybZY9HM5e2uEXOxC80W63KIWsdyT+swLwY3ozLf57b
V/sbOwe6pGJ9NdgWxHunyrz/FRzz6JISRL+39GORyxrrXb9N140fK9WOdar6eqIR
JiIt4nKqrQllSe/9M2nPywFjTDbFJyvJKYymstuOvH69/grZEoCz2S4YcMwOyMk6
MrXDEl3piQ9/mj3cnoJW1xpWwDqXiIgCA4Mpwcx+ZQU/sWLTN554dMxzrxCZcROV
fEUQLe96dGf6YjGGwg64X9vGulNBaZ4Zys8HOQtM1piJ/YFXQT+hiemmTS/aZIUU
pJTRPYPgoiK9EVKzh9Caq7ABT8rq4W2fj4Drwl5li7dhEIdz/DD5V4LbRZyjMF8N
j3yrqolH7tIHvj/yfVC/SZ9PyxDapPHVPtjr4IznozYvZfgDq1dMOvxCPK9qUHTy
X+DRKF3hd6dEE1uAgp+geQFCnbvQJSIPZiQEY5l2hoWtjlMN1q/EI3uUxdPLeSv8
t5xufxk/vfdFkTPvyM8Z469UR+GAtXcfOQt5p37HeFzPYLGWERXwEXP6ReZd9bB6
8mryFLMHx2+/wEj0HNOc77PblE50/5Qu1WJmNmUVmsS95+IyO2Nk46pJc0bT5N61
D+Qw7zaZtWTE2p3zowyi+fs74GhaRQX6sMfaYcaHfmer6JmEvMUA1B6x8iNUmwBD
jup7GPHdBlUDbEyZSL/dKGziHJqPF3BIuDdBjfz/FTzXpqqkb9VYZRkRodUZGJny
UprgzDwH7DgXBvz1rRFApFDACWBSmkPvqBYRokCW/wsIhHk+4NJDF1MyArCjkHlC
hlJ/Hjj7LVKzCQlkzW0J/79DzL7Fs3xC6r/8vQ+ae3Rsba4iDtaqC9I/wmzyMq2R
Tph0EKExvljy77Keewn+nVH9cetyLmFGYKalIm/h9wCTTE1C5FNWBQCDm2eHROTh
BwZxqlYnFmmoUWXhZjdm2E9zUWXdXpaDTsgohLYjXLNTll/SzqH/6hqic5rj8kn7
jTKly63/Y0VxzYgYCOoFyUvV69Ndn4hSJ6kYV6hxJLRSWB7wtYFFspwfc9CpiSIu
lD9L+MXBsWgW+u1qs9p5CakGtaoFsqqmttELf/UTpzqFrGW5TldZbJmBkfSWs+6K
HCoP5SRk9QRXrQ2AOQSZ3DTS+zQwyClkSOOd4GpnxE3B5sGQutMZFqbbpTPFedp2
dOzPaEugYwjc6tJOdHushrdTfVqQnidzifo9DBuNc/497H+WUl053Egi2oeezqi0
HRTDUHbEcWI4X2s+MlDOf1h9WgmB8i6cDmG8WQ09zVKNu83DlGMNZUyvlvckXIoU
/pllUScNF5RXpfd0pO26PUkOznz7bmMdZfwjnOqOwkN6r/v4x+vSCuuvCMxqCYuY
CUi1wIdBOoq2xUMNlXlnygSZnhMy0OwY/Dn8gbwjRwHkVpY08ZUSv1xKVAnKnwkh
Ia8HUGQUXdzJ57rSwa2mbGbtsxa3GW0d3Q+lVFQ6QYyluJbL6YtBZKXjiHLORfgd
eQ/igSrH//qnc/niNBxTltNLI1pTdhpZ2Cd+cXzIFgzhy5cAQPN1GYS8HpWayYEu
IND5m0Thqg9NoNAGE1HrNIjCbqOyJjvlKCmH/asw17fZnEgu/Fr2IJjTxaxam//Y
5DxdSU2q/h1Fzxt0BDfYKveesqa5/+Grf4XAYN19MJbDYmFG+10YQfCQ/PsJwtpG
px+Za2X2Wm1SC3RvvjB1svbtile14+bVs6Nary5fSzM2lKIqcT/v5236H6a/PVvq
9jAf4vaxDAdy3TLtz9mT16FcYGMdaoAc7rIBc+XlEXfUTLvCIpRqUDx8DGPzmLtn
TEAOezXAgnEUVLAhL2iYlhZ3YXOBw7zCLzEZsVnDfKECtK4m5UsjtnLEEApfWSOK
6UI3svMVJGhJFnYRKjs0omMs5x6kRMqLNSRc1MBD6fYDIPGQEnEulBg0gQNi/Vrv
sem7sdbpEuw4CNXrzGc3/GHpkA7SSaAFRsaIXtyo5qRfoU24N2+PoJ+8nMfRbnQ4
E87tlonvddGXD2WBrVC+L9vT+HvASahMpsgugZh3ZKilE/PWWiGbTmovh5HKGrWD
DMi8NPF7s8Tt1PqMIotR+saBwnadWAQ69J4vJGZlxvc76f9RiMIs8OksL/Y6ugN5
X83JzOefEDtDww1iJG1Sx8sRtclXZVpLpEdduipeu6mME4Ypdzvc4lWwCYoj+OFq
F0NPz+O9vzydSvl3qtg9OMfjJDI3ht2cxdtmHRjJPsGRZYQmH2pOGCdJMkFlJpX6
WlhuxVx5R7zevpUEdBDaJ6QbRRqmcagfsCf+S3sSVPkx1EE3BDkEgVsuf72tWJlq
hEwsAEesiSqjcj8PbxvTW+LnPSskz9X3pRuc2vDe2Dl9UlbsClzk2MgP8q0AQ58b
UYf4NNHcQp4v9piISDNa5oifF1VO+Lh3Q+xfnZV/tz7J5Q6D9Z/JaWua/ejcb950
e2GlOMXsAczhPPpJ8fhYOresizbsX8KeddOiocJONvwgFVY7Yj8bwiphb06YnxY2
+vQpM/lU6NXH7EhRokH+iQSQDHclM+K+c9yU46yaMpcQDTPhitAqfDZbyrxYLzqn
qx/KwHM1uA2NL29lPJxQ4Mlpc983DJNlYphhTOk/B+Jdhoh81eww1FC7na/RDnTd
OZDBrvR760e/49AWqyt541uwssFBLBGIsF7ccdDRzlnfuuUeVYqD7p6+yoDTqSU5
iMAOJKbi6465BmcHHZXw9D/kXoOv+XwG4RHaIOXKT9k2562ymxAGLAndBJieoqXi
Muk/lQSU0y/2x3sUsEbrgb2iMbhDteOkajOgjxw7FBPz/JcWSnGW+4HQsYHfiyyk
QAnDfnWFusTyn9tgebeAv8n4XchFQM74/YC7m8vFrrq2TfMqSy6d20l3ZzpMGu8+
Aq45g78PjSK1nuwy5JQKR4VatlUAbt8jKgSu1jYo+w9m/i17jID7qnPUc73uhdpg
XLVbZNt8hIno4QmaFvr9jEo0NsQy0LNbL/t0h47h+JGI1jsvIFWCMTxF4ygTFDKq
ZU+ykSEzKigmpiLgjkUVbBKdFMwcb8lyW7YsfSz8Uu+zs8iUg7mwVSHBXmntUGW9
e1TwAlxGbFdyYMUIODfGr5W9qSgFr5SU0u6ez/4RIEmE2g/3Euz74DNiBPBKcjLg
4O6hMOmC8dDRelrIpzAXcCk/utbMnY4E0ui3qNp1O1K39X3I+vCf2wx8/2US9NNY
C7af9JPbZfEj0N/7jBbUcLN0rwOH+1aTGVKH1R7Yto3rjshZ+W4l0c7sIEZ0kJ4H
NFExI/z3A23C1GhbMCISDacM7ZSiujawvhVEUq7wDcha5GuIzYaVVMCBOFy4T6RZ
Ygdid5+7bcA2bg6RAPFcAHMG1iPezl3z3IgRqtbUJYcpV7MRNm/OhVuJW+tm2Mzd
pgOQo5Ve+lGCBkMfmisVbBD9KJQy2zgQbzLI0hfH4JaS77pTn3/xbZzjyzis5EIS
Cl2870MqX4LSN0YgOParGG4NfKGJW7gYDKjMWCKgbl6xqSaLWlFqBYAahDgSgjEc
19Ruo7yP/nLR5GzWZNTPAzjzY3u0UQvU800uBjucJJJsI3o5M9iC85iOK43DdxGd
Vv7YEb1H1Z8VX9lRlcRniqWdQFrTMCOBPMZu22YMHZc0EPO6smRSYMK5m0xcyyKl
2/icHcxaIIHd0/oTht4KmnIgwOKB0t8KBtQ5Vvkyl1463jrfByjPMC6KByVfeNs9
V0gqRULLpnSvRDBenE8u3kVOKZBCDytZmzTqa39U4Q1MHqHGwjOSmBaAFG2dqxRP
DqenKLwT3IQCsEQG2F81XslGTs83ZNYJoOKO8nnivUhXlqpPxMFITk4CcH2nXVPH
23ZlyQaQVgFrQ5UHiFAGpxloI1zjdn0qGZ3gk0/2mg3z+3JyBf1kMHhB1RUAkR4A
ZgHxRVZId6ekEholda87hK6T48jM2HTXd7puEfre/uiIBv45EIslor0wbkjuELnj
4r96RJqP26x1Ts+PyYmGQ4bJtmHg3fTSxc1tf0Y3uadYx6fztv/StDAarXnCmc0b
KTpzRcqS/V52kQKGrRAPj3gjZP+0Ew55mn/e50IU3UKJzdclKBG7Br20TOqTwYVr
8TVdSFVno2s8rXHjX+vvBU6uyA+0tzpWGSZsNQO0Nm9q9N7vLUOuDMdMPJAUBcAq
iPDOoKtPlRSDpg7jfzIf4jk1tCUP9GmZKtxlTZcvOQLcw+y+onZjvILkMPvyNoK1
vAswMQF+f4Jq21kNXodtn8TGs+UinY6sDWnyBKOWSnzIxcHJeEsan0Nxc4OnAXmH
nitlufpRXGjauPUV+Yw8kweGQWrpPQYbXsTK+P7kqUYjh2xTBWciAraCTqQO/bPs
U1KBgzG+dLlEBQtFd1kh1OILa8nbr87aX/7pzUp+M3YL8Ye3iSfaCKcCfupCR3OH
wJmaNDY7FH6ZZHeWu67osdhAbgDONQrax80Lm/AcoHJKWPea9GOFWvUhcmYuRi4J
j7bENMrFMJhzNXNa7flLoeiab7WcymWtv4vfTKKsXfjY/YSfrmIJLe5CTCSNWFEG
q4CC+1IQOLrcpnJo/DIZlCP68AKi06lE/72TU0zS2AJlz8BOSMn+6gT/aOJnTI2n
qGKTKsiAHwlHgge4JWLw7BLDI4PT1bGBk0ZWmDGwaxepWaxiGz8Glc1Tp1WhLCnp
8VNDtmK/ZLgLEu/BARxEbsViC7lGu+EAYWCO4Tvd8fJ/CuxIkpY+eimzkBf4vVxk
bM6YCL9uzg+j1vOrVBod977CXMzC2rC7ID6u8v05tytRQVJuR5+OaQHM4uWZz2lW
F46PZRrPIYmPB0fBJHt9sWLIYRrIzbM9KnX5kpf7xxRBeHCC16vC90h217gdzuaC
7b0h1TvF5gmUJ0kIbulSrNTacwiTYzE1MLTiB6Z+e6OqceWskHbsN5uudsAm3vhP
zxpqdeX/fDgKQGWedSZO0lNO22v8Dr0IeIbOohB7LZUhTvvl8P//ngXJXAv53vXY
hciH6GXx5rIPJlmg1FqRlrZMGJY1w/A7E++X+P3NCj/atoovdHHV0TWVeBEaA95a
+vEeZK+xnS9X2EVDBuXkQr5cq1KJAQhFqaZXtq+2UWg6VsCHty3TqdylEfYEhguZ
xpekvOT7wpzJ7e9dEyBk1+w3b4xIxSMEePNZR94IsFD1xmCKPkxbDXLNDkLUgim/
V6n/pFHd44aY4+rC75oaJnCSDZxIrjkAr7VSlKoACXdQalzchy5lMLKkJRJYvtsv
+BZfFc1ErPRNpdsmCTGSwvmYIiL/3JKzxSAinBoDMqttMvNTdWq2zOmdtOgJk0XT
MVBnf0bf0v9yl5AGF90pc+7kVkKo9x8uEVSL0xWZ2wmek/OilNqSbvr5WQNGV/kL
FSr2pKktuzFtLX5O32rfu724fRGIqdgp37lOG+jH1y/UGdWaaAfiLgL5ngLhVLGD
HNOzWSGJnOpJcMK+Y9B3DhK2FIsHMR/eeMWzBpsqZIB3KHCru7pnhJQL+tJIPa33
3v8hyNc2Woz8LktASj06IDca4+r+GZmMiniZfIPcdqAPXXRER65K0r/bfZPgFDH/
6/R15iXNz+wv9tNLkJCyBgUJRHxFtcKq92haZJ3HBnS/51P+bPld1XdP/LLa3VoZ
ABfwyNiH3ynZgrF/ZlFacwaw04IbNKvDcsofbTbXsoZ3l/rbULBCQYXTBHn96OVX
tot+nqHn44aMcLS4pGdAEHGdVMhVtgpBMfyWACRAFcX227HHvv0hTg0FrIHaeJnk
DA6X8szqHmEwfshj8jNslUMq75ys9ZFmgxuYkhqwLROdyIgGfGpdNPql5O6zRcE0
5ydts+e+4r6HyBIPs1y3O2ycXRD4sjFm62WzKXzIh30rsyHyMVcxA4VfvrEuCahR
ckpc2qEuUf9hLLBrhWBPZmpLISa1cwxd9NzmynoZTtbL9rqanEhKdgBx3y+GweUR
HIVj2SmhuOqD+JAx9lzx9CYp4W3tKW+6+54sE+MpK0F3IaieAThdS+oMnMSNnfyQ
SblpSLINQ/cNgGiRNMS8LEWcobCulQtcK8dQsZfjX3Il+SvQ7EFxGTiwdPB7E7N2
I06CidCnoYeDW+iqLZsUdl40KoI/QWMRBMpZiWWdkF0OZbLdlhYYsNSyDz9OkqBP
u78FxcKPXkt3xiGN6Qi8w687QWNfVtAkWw1G3iaVkE+uqciQexm6uHKBDY+hEgcN
aY8cr9IltJxnRLg9KiBtgjdZ/iBV0jJPKdGarfsigdbiHP29fvPI+O+QfCfwjkA4
M7AsUfLuuGX24lQ9gW30x1G870Cm1SCRMqNMSAUCPphH/7ZEBcwtiJtKDaC6MAV0
e95Y+zcbg44P7S7oIZy0mEIaun7LPyKV5M+goInHw9oIl+mLwRD48TbTwXW9Bro6
1Jmnbi3f5ktYFBjVGQeEp+eAkRcfBbgh9P+LBKPOgdDM2s9wcZraWrRfhvTI3jPZ
hID+1DGD/gLF6VLE09ecamxSmyywflcweSfy/lR/ZwQmFOSa9Rppb+ivOIZiUavQ
HfkvB8YVVZLV5FcKqVF/auUkwVWkM5bjHiU8XRFX53xJOGVoLBhF3ZbvqUlYqczg
1wUkgmm5tOHcUJOVXl9KCo9+XmKQgJRR7ymhILv7YQqVyikkTc/K6U/doRccYKkb
ggJTi2erTPPs6mZUYa4VmnHQjrJ7dI1bgYi9BP6PPRdt+yI7xdafJrwICVgR9AgS
2yTvlFW4velhMIPKjCFuSIlt+GLzhIuuEC2qoYY8X0Snn/6pbq7t+SEdnP4EtSXx
FltKIJ9Hk3SlklX1C7AFv7Z2LIIbJwX5M1+mzuFLj8NglGN6mlFywoymlNukHwJS
W07UnARoVv8RL8IbbD6qaG4qX2eRG5TLSbXinT9WL4SG+gT5IIB8jCP4HJAt2Fif
vJBNBarH1hQ9h2CkaJLBCQM2/VSoqZjCPzpLsIcSidquXbpT/3/VhQvCUHocn0Cc
gQz6Wg+xV/8VFXuj+ZvARvbDY2zDMkbJQEtTqF6hlkKxlJkZvOI5hKTsuofJptVa
AYG2oyywyEVw0Ecwx0h5L/3hM83F9c9Tuw7uk//nkUY9UvGo/g5VRQwk49AsAs+E
xCRZHUls7tEm8yH5E8Sx6RP8bCLHSTM0FvY6oBKZ8C1C8m1ix7STjjyB8Sd5Aak3
OQ9rIWmNKNB3+FygvpUzjBY/xVpgOfN1aifwk8HEG8ivd9uVb83nPantp9Jx6OgM
nrW0bQaeJ3eFDXiFxS09uuQ10SF8sn++qQBH5SvTJyiYgTpgYxsw+rCWlwueTiOV
OXJocWDVgnw51KXBKNMu46z9CYW0mfVLWO8KFj144rYHddanRHKiEK2Z5cBMD3Hm
xqm5cq7M8BfIV2xgu+YBJtCByaaPUQSRUk3CN//dmTnehsqyxqdIYb4KIQUWAIP8
PQ4m5WhLL9dh2KG43w2gziFeUC00roYW8omu37zwYKtgwMUbdhIvPwV7ZlUlhZxk
1pB7otUQ45f0hlc593C6Mk2vRwSYV0UqPCOaBPsD8i8+4UIqMCHradTpttB8eyxN
wERk1CdrMT9ipG58Su6hl2sOsJFNk/WzBmtwXMvmJ+uE7HcQxV8jFvubhckb0Yb1
QWVP5XDpTZwC1laLqgt3uNlBN13Vq9BBgVYZKFnDoNDbCC0V6QF9Bz+dtZ2XrMza
o3ykO5I8FDT0TZzDvWXtnoqdZmMsOojh+QW31aoyNhYSgRRG23JLfEntCUl5rqzy
4TDvWZ5rCTljI9CkJ+J9SBXxhEoh0Bv69TIlUJ6asZxFbJBAAnhbLypI0UaRog/o
K8DOD6f3JJbmVc4qiPqXYwFXNTk/v/RqkyRt2IUlKHG/YPeIjvGV6EYeQJvOaUdG
4XHC/9ZYGDMlocfeVvfJ0X+5SxV4M+vKNpfSq6SZ+OtuFG7pxXJCyRB7m+8EGQRP
2AXAIZTfO+K8ml6vXxa56g76496clZKtTac+HvoIl9KT3yFWNWWhT4iaX7cq6Lh1
VrCmczQUAgd5ig4ZC8lBJrXZTZQ+l1UOApQr2BBpd9ifBZjAAQPfkPsB0jk115b4
YS9/7FQcVwkf4wDzeJ3D+twJgCL2+JXkg9T1qgD61tu+JRB+M4I9J2H+fA/0p4GG
/w8J7lS3etJzhF4D+NuzEHvMIufX4yWty/QQ6SkuKpTQBfdRUQR9XIlkF/TqijOQ
GOjMYT2AeYREVsxHWsMLIoEt664AAgaLHCJ8DZztoWYXoAOydweaq+V00U4kIeTL
tSQauDLVeZi7kGsIys3+qYDcFinQTWcdmcN4SWP/gAw6sGT45rrJNLnLboJq2keP
A1bPPNeCCIdX4ihkiBOCY2KXKK1zzRosFCNbkfGC2qfjwboj+a80DYAPMEu8+BBX
vGuZlU9y4X0LZyO0u00daS4R6QZU5hACXzjTfAqkXiulnMY6EyANVk3z56v4oOWl
D6IamdDXiqdGbtkjjx3dqQSHowoU3dytHBmozG4cxGk7OCWiPSBm44t0Vq71/QZf
cyAkfyyn8BHurAQez8k0Rsj+/R4aGSCdJe7L6L7G7NqOeXEn8r9iZ8tiVBJ6AehI
23l3ryvguge1MPwD+uFP11TBogGFh/NN3HQaOzQGQzSjPe0cEmjJANk6Q4wkzlG3
jkfYLrn+IJ03y2tZDkrWgJSIl9/X1dIqmcXXxkmqc/IZfoNg6Sswf9OnQjOHwLI8
DTDTCGK8Susm+HNnuKfuL3QT5H/QNUdA/Anrfn7cRpD5b/ovo1tgKRdzz2/4OoGy
6h4YP3fS/j5LMLeS7ZxUSTPL8rtvpHibibl2As9UtfTZqM0S2BCjNS7NfezC4mKr
YvuksAJdZBmOB3kjlvn7lSizmZhJmtNbmUVCaUFePNkarLqfx2jR0b3sZQ+Mc/u9
1xKb/G72jcBcfFvteN2xtuY7wwgLlgmZR/lT+NPUPqvewLDP+FGglj9Cu7n7j/H1
BGcRRW88S9hQtBCxgE5nT14pW0TuTOwY5zptZWiCYzz5Aatv7e7hwo8rwi3sQdN5
DDxgzUcGIcqfuk4ZMKgUGcXciMoOAmOgoYeYKEcJ3QUUASJQGSope2gBUou0lSJw
vOrr0ss10zPhh9uD1ZrL3+9gqjqIemIXExtc967r8W05ZPOyOm4euTUAoh57HYsJ
hFY7hFRiZenPhdZT8ma5T+CHwy1Pns8yorzaSy0vUyLrJwJ5CG0IEaFkqXUUL0Gv
hvaSdAyxiDDcBmnoXN23Vuu18G5ghAX9t/zbV2GR9r89sE0Brh6ihHWBSi5dSsL+
hao0JCICQO8Hp+9yQgPuy0wygc1FhRZpk5Sta5wutCilNFpjN5wJJUsHjw/J6Owr
IcMfcPMvvAIkKoGFQ+qmPsDtjm0OG4w5nFT3tyS1JNVx7vKBaOkqAlm0b4eGZXvq
04c+7I0rhqJeDta4OaAFmjvQtC/hWSWk5U+I2TVty1R9H+5d2ZoZthz9763IR+Xn
bE1v5iz3I70WHlyJj7YYvNbk9miIaaspItZJby+MgyTzXbfvOn/qzMmj9NRMJRDg
hhfjpuRwWJbaLiKJsJkjBvoX0K5plgz/gIDJpkqUSZoAvR/X1hdKB0blX84ud7uh
r6aGisvJZ32Hlxd+V1SfBooInfRy7ipFVUqkRKVAvTllZVo67j4u2ywRSRRs1/Wz
DuRcvsudDxORuP2AQ5WR/BNSjYrVJW1RpICnOZcpvmm075r9y/4A6ftpvt9Kedl4
VMSD6QuXcn8WDyaneBAGTZKCq7N/DFJ7WaZnxFw/YP4qLOe26P6tAMwQlFHa8cdv
vNzDQIRFQUDJvimYZvStcEcpTZnzHwXHc8TFaKSLXr5kK4aCR/AmYpruc/87bQkU
JEpTvIKy7qrrvzwTbttgtA+0pLmIIhDpzhHVujc+ZLBiaIVpZFdWkuGUnmhpUP59
pu+hk6tg2g/OGIrhaOiyu3ZPykAoyRpNAqzwzM5Ecnc3vyMt8ANJb3j6NRXmSwkD
cB93ZNsmoLoDpqLHHZK+ZaZTuIb2GwKZnEGWfiEEX9lXdfjt8+jypx18PqJoZAcx
4vD1WaCf9rUV3SyZaKMEgxT8yA5nyS++656evbBPk/RZ+9AY7qSKWWDzy3hAtlCi
KYpFz6L/plCCDFdPCiSo66eV55zUHi4tnSJJkr3JwL82IcXx5eLYIuMar06SqNUf
ViR4aZS0LDaT1ISxafJQi1D+0EHR0Yo93BLd0apkiNt+rVQIfmDO0IGEHlephYvc
2fVv5FUTBZAmYhLsdKdKe+Vs6YjA53W/M1yP16fxFQUgPAtyaKod+5HUpJc1i59t
abAFHEkeFwAZz+mmG/UCdBq/knEQ5MUzAA51WCyiBC0zlYQMeyKEQ8La6FazAuv2
F2B8PssXSVdFv0cNNiUDpgC/P5sMuRuimMz7/mxqtKSeV4+YeIjUJb+AV9SUrD94
IMRwIo3Ex3l0Lww+BNQYvnAgmEho5Covnpd/RzoLS5N2LVeM6WdCS6DwoXxs8vJ8
VY41CFbGhzMAqVPyCd3IsI06NuD4hDAWGjJvV/uxKeUAAjZ044K7Rzoh2/4RvBZN
ZkflbCCEt3MdzqfAl5cNj6f5dMbaPydI9JfAUkKgv25uykJYToXrZqAsX0vTU8AP
pAj94KslMSOnIOWLuBOB0SlJKnVObKcQGiTqkhYuj7qLEeivbRqdwuqTfE+sTwA4
IrxWB/dYFBBGE1tDCg1pi6eHpFsTR6NTz4mxpnBJz5O4kMf/Dx3NCKNQL8t8o1bf
7G6Fu9PvwXZN4CwDCXDrczTE+y+sdyqdHKAoeZMccFzuG3OnzIJE7Gl7hLFUVNM+
s56kEKFCVVQvUJqgYTZ0syCW0FZUk8eywRonD1QD3z96Q9DcF8pzFI5mwNAgRx8p
SvQl1WHtMznkcjeqcQPJj24TJbWnglmiegYBIrSWfAw8yTievdpz6xI7pgd4pvPH
XyvaoI5tQXro4XpcolynUxXGH8TTTSjmyWUjr1McTLFB7RifIGSrRK4SXCHyldXO
LRik8wZp30O4v1gM0TEOTg/I6I1gl72QvMyo7Wo5TuiCodIvSarHPCaJZ9bNQpWg
MSGr7BwRLvBrGtKJRu8+ggad9QYoPLRA7YmRqYYOmhrY/ZcxQRGFvTIu2O0dh6t5
JYugYEc1fPM9teOcYsLwVS036TK7YArcSgpI4R5eLHsoILjbiM03K0dWn1XLlfyx
muhdjxN6q//njKuaEjPHBHvOTchbPFopTilMfcRqW1OwDXn/6EGOEgqFUt5Aw9EW
RrLFSxkNIDcIJewc8LYYnPoCpwu4a4L4qQL+jHHpla0lCTs2KOIHVoNHsVUlJ6li
JY45+Dh1n8xb4grBOPwR1RBFN99nTEc/38p0XI9b1pNBXIBVk1YlE5QjIy1ALS0C
TK/tnRG3A221j8gRtt9XWEwbtkdfsRFnruIEVtfsWK+sShlCdiVp/NmYozBLUUY7
RP4o6lkqCqs2yhO+xf8AcuI3kROvpllJshKJO/eGxwqGuuKW/O3iEz0mfkc+LwI1
MH3pS+kTnwd2z+wcNMCYiFx25Rg6WK7DO/VWVMI12jAXNtqA0h7QnjgG7uRrO7kl
VsjI2JEbTXGG32hDNZDfucTsuRjKvdttOqfHn3wvWcp5myAp/TTADMn2VGeVSxhO
iJPX1wYPDSzwN6q8Tv477EV0BTwuz9KZK53Fv4KHwAXRBf+0KK4jaDi041Hhi66a
4OKBrhzHv9tLo0TZfFW5MfNfu1jdVJ5bUUI2ILSkyc0li3aITd3XoJq0OMAaNcpx
Vke4zY/zF/jTNLxTJzAhEw83UYkAkXuMPZlK+ymzj5DV2rzoHXaPoAnxN/aMrtzW
oVs2Ed2Al0+Pgq35Z5HZlpK1u/Ohw2vc7HMB3V1EJqRQ+Mt20m1mFgaBZ8E/xrUn
5YLwbxumYACvc0A60Mk1gp+VSMzjJ+O8/vRdJg9a39ZAf9/tg9B/EdAtrAL1oVT4
aOjJo9ZRn2XHKeLQgzzIL7oQM/GW3NGx/eEIzWvn11DEGrUfNe2pzJdPSS9oUni3
EWPim8VVhbVVhEnet67GPmlOGvbZs/26jqi+QBVkQO3jAS21y0rhEx+ZmSkX2AvY
He89eQ7nnniTIVmCMvB1aq/LYUCZdUHbALRfArcn/HszRHBK73s34nu8hgc4JdnL
brTtQQNz2CsB65cfb/tk4BMURb3xZ6C54J8Z8TCnIM9HPxvMYYaqIjTAgIlEclvE
0dRdtFKLa02ZtC9LUdP30N0YX6QqlxKitNtATMrmrCbfl8BWJQ0DUt7QibaVZAdu
csxPbjWo6sCZ50va6FDadAc5aWYXRicquTAwPOPmtVHkBKe3QP0kHMT8Xsj8jBKT
veYxXTPU0oTJZg+56YQFnrWTiMfJDUzKV+L/DdlGHjfGZiMwFvcx7tqKcVWhuBDw
BYIOEeBNnLK8xf3hz6W015FVv2p9O+7yonm4zvMd970oxnXOkCXnQsRpkVsoSvN4
iE50wjMzgOKSBldonYVgeFOYgrBtE63Wvyi75DKi22TwNdVIh0Yta2RjMMQWZYGY
Ar5Pb0Ok48BOLfuFT48ptgpCH1edJwfbfCqWYVdJf/v+XsSMcgMV/NrIFxP6mtp6
0oFTe46squNalVA4WL25xC2dYrBvsJRhM0Qx5xDSrlBbsIPR0FjHMRc2J+gaq/nO
Q+c6g8Zd9Ns+iWiiu7XNAau8XoEivJX9tcWy7XGf6ZCuH5ZTp7JwDVxwcqcKioRj
SvujXXW9fJaUMeIPOky2TTx/ImLIVC+pDDAdJ/mo03QVrGL+b2KcbcMkZj5Vpe78
XaK2NIoUhQijRXfA76BhUb8UrZML7dFD9KzBgYd6PZJAmsr1r1/LDABOAQJ2vkuG
B2KK9x1h7WFR9C63NRB4lbugsT/SKRITXxBQlOWlMIvEyVgboOIjdus5JLvwRvdq
PTJlTdocMtLR4HbvybhkcLJO6NfpflyLEYosFKa8jTt2HxhOsqfRXMcDhFyxgRCk
SBLcpcQwgNAB8vq2NPkPS37mgV31EzgJT172wy3KtgXfNKHY6awqKUzAlB747KBc
7KHyTrQ1oNPH4VHkdrjxgDXHQM4wEPW+dRl9GnB99wlZUoWLvX38CTvWKYxvQgHy
HIuNZETHpWqV74jDtApv1wFm71Z9UjBw7AODCa9BwCYvanIPeS7NCIZn66xifDXP
aKDXnIoJvqePhrQRhbnOaG0bf83YWG/mqFWXRg0+CJh76NmOJyLfU3rivwfHWdf9
VDFDwSoxTPfBn6mrC84qfeaV7Z7yXj/f3k5/zfGMhTsx3N9xuSqEmaURiT/a2PE5
QTLnEF2QgfZXFYlEpQRB11MsiKDEMqGGYHTXO58SWuzjTJPSqCYL+BCJhxR+7sGC
qFTEabHI2izJzVznlSSJRzzxexQk4U9uOZ6XQJzuPdGFZP2ijJlPWeX967ETUIio
KXOWpAClUOyjZvtC2ODzDde+WypML9wvW+s0i5eLfsxMlNimbGaYeSYgr1TRbPoX
/Q+H1IjiCuoczQMMP7wRhMrM4yyHBbxFUBY757GIUJvITU7V3M922wNrx7bdG/5j
7oTipNzvbxHRI1zU5g2o+OcN1j2RLlFiVAAv783H37M/9DR1FLz9eggkOX2p6Lka
HYZLLShU4rLQPM0naAupUAetkWdrxqoPj/5vwNesSY/fP0vSE//nTy0q/ydXqsGN
CLScSM6M5ahywcjFizmTtQLKLMqD5HTurbAlom5G1O7p8acdfyXSi/UHoS9LiBm+
oyNw22cgB0nDtWTB+/gc0XCOyCDWJAGwZv14XoXxRxszCUToilS1EFUUaT72G/US
BQKY+O/bSJtBpEp+BCMiBquzYDLwXEBXg4sZMXmQiWqW8Ve0qbmCjrgdjPtK3EVj
Wp3nuJlRLkzRbh2dKO8OknXAoguI/YSYQ/2DRupKwBp6xcEemBZ2CQbkdcZsVVPk
B3ftuzEv/3gO3HrlinYlLmAeC001BEy5fv7KS9BZDkx0TLw0NPUoAdVjNtjBAI44
0ogTeIiJsmIfhlo278jPPLKFt8PNt/6fDyPjT42D1ACPA9fQEW5pGlpe4Y60Ha+w
CgxcWwHtVTsN4lYfcQaHjEUhbzzD+4FofnjkVN2ahCheH9gF5TPvtsKoviFdce3K
LkmE0dXUxKnWcVcOz/EOwOwdQIJAOCfGmiRM1AipTBpeWbknEmfemrPzAYMr0ltz
CLEnWHuTAPUKNIEBk2TEcbuFrM+cY+bYAjHkKvjV1dFhn4DviKubqE93Yx8/WLrD
ZdHIIl1AyUHzd63Plp1sa9cY3NqgDkoeJgQqWfnAZqy3iarSss7Mgm06hKMhWU3K
7Po8WofsNsYhVnkjrGysitzwwrLqyt3alh0RlR8D5bU99p0qOYqEyQ+NtEVtd/Y8
91Kylyn1EXX/QXqTHZaBN2eD5J/pCev1QSdH6FG/5Diow7kaEUslo7u4ppIIsNN8
YpFhqlm5KnR/4bBImSUPX2lIXkJjnhUS3tuKMst2F19kJ+6TsY9lDU9J//aaY2Kb
K3pDHe/qYwWn+hIuaElwSInuxoocmoPrlHu4+4Yzr2kK2yNRfJ1ZOiB1TG85rvDU
0yX91raDz8ilb72gQ4GuVmhG/csGiuqE9XMPhqHEoGnF4dyUikbrr/t556YVUY79
wV6CY9XV1W3t+WkpGynl6ZERx22f5coKWocuYKQSXGGKw0i5S2i110ouglo5DB/p
HsQ7E7VfHMzlRkClPCAEBET4uw1YNCgcqRL2SRtRV9WT1q1G28DNG8m8OwzQA27H
yCtzf3mF+KyBOjr4Fl3UnVCS+cZIbqXXd5DBkXIsONaPMcFLKlHj6DaO1kPpd8Li
+VQ4DcGOf3nOp4Q0ua9RyGEVA2sJs/1ZhbMXHLbtRghxuBtGduPunnHp6cFn1EqQ
eE4SEBszE8EqTYBSTgqCujE1nfebiPxAVde+oElWTre4z8rAQhXJX7+KYn/8Vkjd
XgINGy/CGpZ33T2PYDaQbs29nu6uSjpXVTH0YHBz6HuajtIbaarzvM+9VXsExujv
2MCIT3GeMn+6fmtJLgQP9WlJuzm2mKQkyRQj8pILOSxmcvSwe4xhOHHxAXjQ/eck
pLcF/y1nqXd2zMbW81VNpV4HDoWvUxiZSCKBkSjdp83byp8wdboYUbHPQY+FPbLc
/SnEnTQ075JJI0N2q92v9Zh/Z1N1HQcYs9vjcN/VUQ3EQW4O6vg+6QhdsvqGhXlM
0DtBdRYCchllT6Rsg0zlcDNwGsE9ApBcQNe6PBVtzlLdCBAgPlaeuLgty1pu+3f2
n5o/9pMQpMdkAVEHyAC2WQQe9sybduIey7PdcS/frebm6c+Mg5Mu2UF+cyu8G60F
GoSMv1nlMRBBa+EM2pxzFY6xXholmHVenHPisEFjCZZjucarEpG2YvxlFcgvG5pR
d/2LJtkSj61X7CeuOxHYDSi+2fhtZpcTjOcFuQQDL7k3S1sZjIwWrvIBUGaYoDRC
J8medSCx6moI/cS5JcXjHwRx0fclkZ0rH3KsFgxF5mq8SAM87T5uGR2jqJ0Ei4u3
antBR5797RAckOMf3j49Jwu3q6KN82zpEI37h5A9PZfTvflJJSuA25pyC3YLf18c
8JGTChF954vbSJR00ktY8g1U9klw4Rdxs9Nr47sSYdB1DuRRbqJXKvNyEass2jxy
MzWD5td2nXySzFs5Q1+665apxfPRT90MKcO1ayatx+EPhPj/fY8xoblhZ7ZXEc44
uOXBzakuGRQy4pdyFGpN7UQu4sAX1xP8v8VSg7H5uAVKWtFb8rHb1KeKTPFrdxgl
/n+Tn4UDpvLH1LXmRrBW4kIOLX/t3gjuNasrj/l9S+EOYBUbYPSmVfejeCwUaSo7
hQYswj+1NUlucBY5i6Mj+w8pJEbuJmC+1QY6D4VJj9ScxsVZXDewmp01H9/GAzFO
oBhoejCODHABAy9//2ulatrwe5BPTC1Ma4aTWjN/8Q3XU8zeCVJ1i2rKDDPKUEp7
jFQetHDRzk9gnE879QRvSwH6Zl/VMXNMYojOfOgYOeqYiPv1kBtlXGQ5Lf7w3TGZ
1L1JNJXRJyXisP5CKk0SCyVRZ2kya3ZsM2DGXcAfSC/5m/ppQq/aAQ/pve6W0eOZ
gmLIIArOVAfe7rROYQ6dbNu6iu0C/TSfS5PrRmUgWQ3WrArfsXqBmet+Bipp6RXw
hmBNw202kPYVEP5zdq3tNZAEpJmTZIiKfI1nirZcqFhlCXwOP/W7wfQbo+sSYqXy
1AkJF6HZs39M3vV+r9oXqlqoSEfOCJfFBY6HeM76Jc83EKYRRB6DjTGYq9/zpdJa
likBRir88R6UdFiskewoVxueIiYGYGgOfxa+ETtPUFmm+gflpcxDt3sp8OPvPX6D
ow4LkwXrH/D996taYIY3VRVsv8Z84llFxuXkCCQkVY2XgFhKqeHmiSSS8+gLlRy4
zOb2BnwV8WXto18HN6NDBr0Kd1xISfilpkwHU7EacUA8EH2yBHxvp9HW2V5bM5Ry
4AyjW63WFcZt9/3aXxqZZBAohj8+CdQ1RwW3B85ve80mBguqPE6p3UDcRE2dHYp+
qXNPVreVK8nTUiAI6rlBtmvz4A+A7WMuecrfADcIG5rbJn90XfPw9k0w5G3mBpbz
oWKxqLXkMnTFwP8nvie21dPT81LMxPFhbrBN43gWcUSH7w61FGVcEoOzzJvIDgQf
mEusk1yTn3R79toEzZsikNh3sb/6/f+m6GiRhHfJVBUU8bj67xGKpRa2f4vCMNLQ
uBaoMZwblbPTvbbR4IAmD5mZs7/LdnkhnO5R1QVn4283NmYMlUFMr8QtoZuvvNQf
B7JT32REGU6fqc2EwTz3pu/ewrVI4yt7ic0gIHu2MHohR+9F2C1y5Yy/oaUPV6gT
CrpClqfTdZ7H4/0ht9VauPpqLCKSdr/9xkn1U0efV+BG8HffoAAqwInCvp4TtrQB
u8lvpvCYQSZrMifqbAJSGtEMLl2g1VC1awclyhnl0qJ7oEm1tZxk4MDn8jNNgyUY
C0pS4OgmgLa9TygiLLMB6b+8voeWk2TojAcDF8UAfm8AJPNjKbIcfQwzwCPwZl2g
+15cIrkfa1CFhpk+AUdDWmskC/uJyP7BOZy5o3Pf6SPEIsll5hHervzoPvu2aeai
VeEgy6YIg1TjcGL8MjzFaf7KcC7CWDyJcS8HvFLOTiZizxIOclY3oHP8E4YOFQvU
1uK5e+GD1n1t5z3JSgBZbFowiJ9AoSpdt5PrhYffjne8O0mevT9qUvPEy79koLiS
B7VLIViMbXqjVLQKswI+AvyNHZj3SxRQL9byXiRlOidIf8RPPfOqF+dDcxSHWcrg
ZX7PigepXgGImkW8zN82gy+eGkH3BTtCACCZPbQC1uGAmJM2Q0lDdHEtzk5pdDLI
mthIpgNs/jA3JPX/B1IIOzIEDnyym7EZi/RUGb+cqA4YvCtdWDHy/Gttf9QwO+n6
GMDP6DoQdSnpmKcXI+LVggwJprNyfOs5cSNMJ73//bnCmb6iIkCIbIAHx+rHiTp2
r8/3dmlJML4O7YM2xMfu2eYycacwzTWdjXIi/VnvT57YcY/bMWqrLEhraEdGBVZw
HM+R/wsr0jjKuc0SuAOhUVyYGYJ06GP6lYYkyMrYQs+M7tVb7Vb+lM6k/GZf+Svd
hNuQoKfpI6Xa4rdWaLbAf5WS3KvuTtLbJCL2desSfUe0rLgkxn0PODp4+V9+TMKc
4dOpQe/vfoLMR+y0D6Ntnl8LDPtXyMhAu5uz7164n0BgHCTWwmPmyHjVHLcrySST
IutfLc0ZiV3xjBgiKefcp4FGT6jglFAp2wqTYHoXRiA0eF1l4sQyJEeZ2dqb80D0
Ma4CD17QRPh8Zb4Rv0wHXdjqvqaHBLuIeaxIiEspTMTlWjYu1LT8Q31CB59FJ1Bn
BrIEabZokPF0/a2Rgae/PzuHkEeev0VXke+0FVTtHZ5wYBDgHiIUuyiQqBAHs4So
DpBk2ipo5pXYPyuD4u7mgsU/maesijn2pZ+vOutpdpCA3kKK/J9HXQDs+YECe4j7
mu+W18uEkAkKxmq/aKfHebkEoLOlILpJnTEDM9ov4LjqvlplQ0jC+3ClM+n6lpf3
fV2SkTelm9GL++vtZte4Qhb0G9fuRWA32qqwB9PuniPM692hi04adVqxdOPZPwwg
1aSblf5Y0De/ggxRUKfIQWGYS/QLyNdweuaOoikFsXQtjErkE3oBa/HeZwBXjncZ
VLPGV685O0QSjgBYxE9820oqzEmu1JlA6S+qakwn1QNuWBFueZwVzXAdppCUkoGH
x1tpCe2iU9J2qVeHMkUBI01R1d3YaYYQuC2mmIqQTt/sWoU8payeeuMI5dTOTrIf
x+zWuL+uddffT3OeXgyHDowcgSeSc8gArGXBWGwqyNOv3MgqxWTJ/wKW8QLAuLcA
qnQh++JkzmOX6ID/QOsZmLB+Q/0BggdnAqi/TUAmMAdWk0lCcUMXWoK/7vZGR3hE
oYW686RVUw9z7yw4NNWhyocmZPpMf8KsxqJN6wVp1yIg7WnL3XGgqJngojk23RCn
kk6sBrGIZL/7eJip2cNyRKvkoeJew/FIFF1JvX971psK44Np5qzn2S66TrSEqH8N
A9oncOYbioezuHAG78l2SFNPP07dkQYEXRN9eI6aEi0JlViTjeksymH17ZBmG4BS
OvyAoxiE495upexCmNXjQjr5SlAFY2ZPVDzofvaOCsmDD+Phe/OK5DnVo8H6Udbr
lDe+y9XhOIH4kQKemVfL6zWLHqnbmHv3tlHngU6Map3CO9dQKsmRGfDARXrcUYAu
XHJnz6uxoukwXSnS2Ykp0JjvxmI3sDgcLpmzvwy880B5Zne64iQV/iGrFKTZ9/7U
JWpfC6U/BtmzmboetyMr097Chy1kbBVSEF83o+M9MrhynH4GR6IYfEsCd1/+Eki0
aL7d8QPA/64a9RA8rYoLxYAOUK+/vF+kkqRQyAiJbYUhvhsQ2/0gZLqcBKZj1+VO
JBO25C7HK1wEWDMmkgd6+VLKX3z0XLydLCMSm0Am1S0RYjxX3bHVhNaEHcFlBhKx
HsaC6eNGKszIOG70DWriHYVPWWxD1863j8H4T8sX5uRYT0LF374HoVK4g4sQsCR2
MBwNOYbEbOXt8VjNb6v4cTHN15hXgEwlrlXEKCOmAsAwpYufLsOhcQHaYyxvmlbj
8MG3ZRGREdmLaeq8w1UL/6smpyeGXKjhAhp23OoRHYXHWFm9768xamzaJ3/g9pIA
jHUb5nhs2blC5+UA2TCIFNCv54RhEeDrcp0vEcK0QOJiLp8FWtndnbmQzFkpeCW/
UbMTKPhgtSvckzKYMABs+Sje/0CyiQU8dNMZrabfI0lMVT/Xq/w1/W9DZQd0wkiC
Qj4f/8E5Qv1pWWkn0BZBVy7oUTIuioWculsQ19KObden6WRTLo/be1h8HEPv/Lys
WMOLPuCN3TFBKeUFJNGalOR8EA7+INkIGCjz8aFR9+HW4QwM6mv3ntQfgJskvQ3n
k2vQ4ARJdJtOaR0VjSfjMIwPzYhzd06ZuiKQYXompedylas8R/1v5M+iE0gio83p
Ywz4TKvAwC0Ap+o1/1tvvR7OJTNcj0UhZBh9hNHupWX0zov7SfFV1GHvxUFAwidr
19CNJxZqS1O7IA+NRDupj4JPJD5rjaNvFOBTaJyFKqThUxp3bpEviGNS0w7QfpIT
aBsQWvG6AoTo3zCSz2GXTRhDXNB5egO4v38aQDZg0OALN3S6ziWxi7crCbgfqSbP
P8/xHFuzgLgCWYr0d4N1qAUnWFUN6z6AYcV7QI/x3vYM28EngpjGZaEqU8VD+Rbi
Dch6oKdlDaIC3jU3p1Zn9DnLBTkkh5fZkZOUT2G/raMv9Q6pzQx8HgLi6lWdYuKX
tNnHQe1nqk/W0sqLRcr21tlwI2kP9cq3JfGQMa7EE0pWaJRtSmf2I7Nq/RZjIA5Q
68pUj/zOE78HKNOUyeodRWV3apCdT0fvxdzS81WcrGv1iGLUL+eV6OD/Aii1Oyhk
JnEpZKBC45PqWFiO770u2Txdpxofq2m6Y9udwI1rU9D8O8p054JQ48uWqZpcrg7r
U4ZBhAw2rgcgskQBmbEi/SJKLF+ojSJwK1/Ra1hRDCOd4+HnzcX4s/c7iI7+AWp3
dmzkt0a4xFQ5o/CWqP7T/l5biFanldIzaf7AzA+RS3AT/YPaxTjLr87tPNhSZcxN
879bxGqvgGmSFENsYMYLlUuahmE9TDKYADlfEMHCynVYMg1U6fgh/zFccZEsiMgS
SM/3goF1fDkuB7lo5bisdmlTX02AnJMZOAbJ0EIzcriLmTa2FYXkXgUreHoz/dtU
9WZJoubs8sG5pEidyKi0olxSychUXTsXUTc8QYtSupIiTwBr0svFjFp/HVWUg16a
5m1ZmlMd6QdGZmzBMM4WEMSwnFZd0BCAGUPzu8iYIQ930fwFRtav910cDgxJHYja
LayoK5lfaZ1C0K9pM3IkP3jXlWUpGak60DxmozM9ycFbWyUZnUosCwBRtOvv8OwG
Viraj/XX0qC8vJkHiu3Ud3sf9hVLZTim3/X09Cxv/ZJlNc8AKc43O7msYkWGBsKn
A4gbeyMLHdJGZ2lrdtNGRAL1Q5y85JwfsEsbrjIkiz6K596R3TygVVGzZVUJRAkn
6wCtOcIpRQ6F6k0SkVDCrQ56F8dxUtqi7ri+HjQsX4/0atOzxnKofMe0l0Y/7Zgp
GlKQvngZ1LJt7QHVyoSmiUkAk3DnRxHmtfN322LqaTuB7xqCKd56z1UbWalCi0LZ
XF+6j8IFE6L4jUFTEb+TxIaRe4jwral5Py96Alqxy+fc3CZkTIpJl6CNFkBevzSG
RQ9oPlUnat+EGAoDSgXympDyn4qfFms3QWreuOY9NWPsGlwFmhJ+78wkU/aJjiNS
bnmYNxLX09kNbb/LfPAF7dDBWgqYkIwJRxfq8ARrWwfstcHSzOXAyAeJXyazz39l
m5g8WDOSgy1i28L5NToba1BGZvsppH9S9Mvy3hIDka8jhs2XR7mGlO3LAvvBSMlo
oEXgfIVCUJ4ceJOvzJmTAjYVwe9zfMv0CvHRv2aPG/RDvy7RiXBNz/bAeg92ORAB
lRJSmDzCaH5K9Km34OIafUwwld5IBSoRrMGKIGDm563417bLVBblGkf1VYQDRNWP
zeljVeAZVKVFSzW30MNG2d5W+PU4xlfS0aLkz9/M3P1HTLZfpJEhyHa1Z0DTFZMz
CUtWAIFml6dXO8i+qmoZzztMzpDPqac41INOXdnpqgUolCgZTImDIL079C+xLVV5
HhExlE78mN+yFn9W54pVxIsCBeO5wmP1QEXio5Tx9/U61X8DNsGuu5yZhVVod2oJ
2+z+3O+fhDjQbS7cMMTBlv0XTJSjGU6IdsHXLVXHkH4wVLjiCuV/b9b53++5VqPT
5o9x29hwL/gNuwsOzJr53tDFRzYSujzbn7v5CxDT9xSAtn0G09WAXwSA0WMU0be/
sO+ye/MudqjyDsREjjdLQGG1sM4Y/OrzeJKsa+5QCuZogVbqJZhM7Ts4Yv9GQJNm
aIzK784n6Fu9QcUC22nc96nYJdedzMSuu6/prbGLmSRDVmf0XiObT+0U0YY+LtTI
QL+i0lZ+gbeG4sVxvPIJH48hkNHUN+NN3zhjlcVQ1xhVagyLMIPSxG9xxpco8ieD
uz+0zwML2CGx5KV9xTvlUdfZZXH1VsMYBF7euozGR3wECYtQb8is11R8bvchW+N5
ywC8Gu8Rvt0txbQQTtGsOZjVybdf3T5+CDCUdtff5f+mQOcZlJOZ+okz6Izean/t
hLMvpJTOO20JISGta8lZFq9Vnk/CBJPoCePmiYDkmIRZDx4Br01m3A6RQJmZqO/w
0681qNTCaLilgXECZ1GNAwQH3yc4K+lBC2Ly4jSSTNL80HdGJwB22IaKJUx9MuCe
Suy21w+Q/Adi8GXHBw3OhzjgTo+kb6GnT3DGfj+H5Z9+OdU3P2KCFni3ZEqme0P6
wm6spLhys7RZ79lXZN/iyJfcNzbs8kVBtYjw8PKNPFcgSH049ribT5tMT3Ogl9z+
cx4C3YUzC90Y3ZX2fTtorBT4M5JY8AQaX7o+2n14Du2DFNkWCPTASe9WdTx64zEQ
nHl9x4ivyzwlFR65dTHj6MoywBXJrxbgTWOkcQySOqdCPPtdllawzHPnmTl/UDup
yXLab7n5K6JSvHBPgnekKnjPBpSUQzM9h9u+sm0YEAErEw76UiCWkTPZwNzlybJy
lTN5lFFtvW/m+yg81KG3a/yQ6766tU9xBcbrDp60etLhEAy4n9iH4GtXCP7Sx/zG
ebllioeIgVQ7dkfaKh9Oo258IMVAQ+B5X5KMeCqD60Z4w3lQmgOfwPt5hlJ95A5I
pDUMFEkbgeS7GQNH1f3PjG8J7JO/Ogh7wwSeW05ixwx/zmJofI8e/sm/qxhdxIcM
XOFGdODgyhKrt0m/i0v9gqNVfeBBvkCxT6khqw1M4G/yb1F/OcFpCfnO/VNtIXq/
I/j0SIeEpr7yZZbxg7JoZkpJgKigKPtsySopYU3aF9exZD30XaeeqbsYBgTnI20/
dpXrnUPM2URCfVef9LNkbIw+qZ9IlU+vdxJx4E2mhIM5iVR3xq5rrXdPiYZzuMF5
feHFQh5CYeWGnU6dy98mpjH9/peIGkd6qHGiGvR8JQ/QI/28T81AtdxA9d7UGrZA
97tg7gq8ko0yYkgwk2K/WyuoOC9TXuiz+5TbBhu88169lE60tNg3LCqxpLBoqFnh
UOWr1eXVI276xbEUErnWNpmmyEnkg3l8NWboeXy3CnlY7gn/LoYwe/aYu2zPVbC0
sTMpkK5eVeX6UXnElEEwSpiWkXw0mGEMVUkSM5WWh3e0vI/2eIDnObTPSsEbAI26
vblmL6c8IFwe4T1tzY8Khi4Mt8vni+ToCKUjS8NmVXH5/+Ck8O2Q5UXKLPf80HO4
1fWw2/mcZ4Evl1kuD38WaIyhtXGEokKQa1qngDdzFFRkB0Aisji/dT1T4wQeXwRL
FS2a/SRs3JIXpRLoki4wajg01EpzRIAaVMgJStecU7IaVPs0DxV3bGShpc7wTfpA
puJ0mjMG4sTNXxEdGC/jW95SSsup/S1WJrpk3jE4A9NgPEYoIXqq6w37l7/J8zTv
/TwZ41r85SYBDRn4qvLR2MMwLuaPXnX3Q+DjRhp76hw9d6/sNaTvGm3ZDeJiWI5g
i1VtFsJ3A40RA1Doj76BJjAGALDgMd2sxNlhCwLywHqffVz8Bo0elnqpsU9c/G/O
JvzPn79xbJr0S35mALkWvgXsTBnCWnXMHWrOOSJMD4FadDM5Vp9J8+PzPAmV+qEk
5RajlbgOS/XRmKML8Q51hQ24p74EJhkInd+TnUHNv5Lxw9RRQ85OmT2amsZx1MXf
RWdcDA0YWRYrXsBpSrl/pbELroyaCXLMRpkKl3cQLdf+7z1uVDjAZ2EExnk0X8qf
rW8riP9ovA8q0l1nVb3S6qBlj3htm9/z6Q07qKFx3K50pXWs3I+rLmw0czu1vgpr
se4Yy/aHbLBBmnTPQVWV67rYYb8VIO5MnnLyJ6v3nLEljv8LMxlnBBCR++EkwRSb
+DqxnJf8DxVIfuShrBpoTD9BmpoPxzpAizf0fx8Teb49+oASD7gMtMP/4phU86Yv
ckEzs2+fwdjODpwCiPuvYFSQx6S4PtzyzbEGQXIradvj6x5JfsPTx/9KFUIlDxGZ
SRtH5FtQk0h1iTquEYw+gyHw8uTYDjtyiO9vz4HA6INwFIwtkh89E/3Anq8n67Ro
Meh5p5xchwzbX+Lhp0R4qJvObqufs2p7uwdAZkfUVcDYnPSpYTLNju7FjTpnq3j8
EgOSLb4AWuSGfo5P0pp19tQit/CDd7JJBkdwBzyuj6TWK6pbIDHlB2vgQiR2PN4n
PtR/xtwyPy3t2yc0RGnqFaWwo/EDyYFNeZzinD6P522XD4+WnOXrgGuIJeu08iEs
f1WaMUG9xht922h1zG4xkTAwUnZokd4u7fSB+UGfgofHhJDLHgv12/A6DGIJMkJv
w2YnkGXo1bf/iw+YJPTK7SR9u3VjRGgWp3mPIhftg4qC2koJz9MAejS/wfzc18Qs
FJurrfRufXb5evcWRopJuD0QzfYuAkSyfnqnL3FXzd+ikDa2RKDWocxy7I6Vime9
YT9nk51lneAqDKjqxXhtxTEswrH+vuhs9aaKuFCs2eesn14RxuV3OFgURfcvNgzz
ZhBiCjK+t6oHIy/Q2l8vsp772nHnszq27ORKa3+dJhxXHC70xFITb9yPgjxJlw9k
OqY+SDCvAKqKsYp4UBE1haD7FT5IUhPdhvzmVQ0j7YX/oLcBcnUjQCYQl8l+CVAY
DHwFfSCXD2XrhGUVEEiFUh7mQPjv+p6beqLGyT3Nj/fs2RziFdsR3IrP4Q977KiL
FNajMKKR0LoNjj0MkNpNh+W10bIw3aduhPDMaCceJCMyDJ5QyD7dsmXFlvfGzIHC
GdFxl4fQV6Yoat5u3Nv3sq3aEmC8iu81o1gSz3JW9YquHy+xQMfXVDa+iZEAhQtg
xfmbgd+InXk+nXs0OOa0HVaASAwZPfyEf1nWaWdUyLTg4Ojqx4XK0gDvk0wxe953
xaUdYyUryhM23OMkVKzomENJfcPCpsNWcZGi0HklFklyBg59CanCxUtknaM9QE0Y
E3+krwTAXnomxXHIi6qNUVXwtsXg2IwUi1XeU6pBhw3FOJg6oRlEF6qQVjNS+RZP
zt+1La24M+vnqyjvO1ag8JXB8RJXQxoWzSLMHRHcVx/A/4Iv7cgHHn8+wifYzQd3
Utpmoybv64EwdDEXiCsHtNBN0rSwtw9csmGaIOGqQB0w9KFcSuLXy6vqySA7KfVe
tlFwMnoHrBlDx/tVHgp9kKC6nR7mUBhirpNHHCsq8JVZ7k4/0ZZT9fIymj5JfhtS
5EEwhPRwzM2dYrUEo8gHZfRsdFz+07/jUeG83ZNCMoSURMhiGqSrX4OFcAwFAa4B
girJIhK4UnZM+dTTK5SgEHU816lVIjg6wSVWaO8dtCNht3evwwFUWihk+wi30cCK
xHmMepouBZiiSEjuwXmXpQfOMMOqEfSq/YkyS86dsmiHBcvC/Sw3L6jaVWt2S7+g
ebjFVh0dhh+PQaXGFMLVx5O38NxBqXvHuOZYca3BVTVlkdMbYqYtP6yrnj+qFjDQ
H/wXxheB8Ohr7rrZyeOKVe4jeCNj32JJkzczZHcb5A0t75ZNnGZVHAHzmrN0a/Kk
JvtkZcpQUY6qHOqVd5yLBvYQqp947QbW7hyK+QxwAmM7bGrWrQwE1c46xjTaucnQ
lAS80+/R1gRJDOgwcWRmuR5CHgyCwvjjMkIOL164iTppW06rVdtqqTIY3YtTUHJf
RN+SQMkbBUrUca6KAGT8UIUEbpHuhReZqjzsBWha/7fk/g9SAjP0rUb1gcllhUjM
1+Gx+moxKKW4WxhbwuY6fB859Lc3MahRR4/nrVR+cA6D/kUlGR3UkJtkw71Lk+/g
SSApbIc46xWxUYnr208yam2f1veyTYZbzCaCYQuMHZSxGocBraL/HKdCi0UWtGEb
LSLgVrKSDO3p44Oy0SlEP+YrCB5W/9AbLDTMRJADQU5y9LmJu5u+vfkATDSi9ip2
EpFjdlJyK404JqUqKthzunkP9Fy+YfVUmmNaX8T9NCnNOuWIr/T4azBtTyL2blrj
YgrfH0c5v2Znd5bfE+9s7bmUoVTGFvVmQZrwBsikf9pYmekEe0KSQVvQfQV3ftPi
TEZXK4oELfWooD1EhzKAZF7weCBcr3hgniiR8od284ogvRDs0hrbfN7+01gUSHsN
8cV3U/l5SZaAn9E1NIxRj87cUleOElqcbo1rHyZ4H7KL9T9P3Qk6sV5YkTH6Nxoo
kFKvbu/kHy6YtWsFJ4KO5gN5Z4BJEO2E+PMpZCFEpT8MmVB+cbpSWYJL4YukWVdF
RetpD67rkohrLobTRrPwHMOb1QcW0MwXwb1DUK53CVo+TejLG9qSz8oVDmxw4qSL
cBGN0gopXRIYD28NzL5JGfJ2Q/cAEIihITqgxDzP4YLa4sWkd8Dkzv48kKREfRnE
6ZCNNbU7dLjseqO+C54dA+jMpT8g1dFWX/BPwCdABafhNv/Q85gWfYL2b+fAomnA
qaiygLrcHL/9ONCNn4irBEqQKSW4pTpudbL8ttenKoOaTh5ftIo9TRk45H/JiwId
XhaKPwScelT3LfN700tG9LnNRaL3/A/dQNR6s8P8Rs+tzcWHc6n4LbH/oRJEyREx
gDy44DLFvrEFqkVDkOGRhQEIZUzFO/73WYOMGVr24x8yTqVnDhRI5RFEzC6426y5
k0szX9KwK80wfyAJ4p8Hb0emrTCccJ3tNYuxGoeG0WtbGpyahzIoDGS1PGQHCZZQ
rJZnzEfbKhp1LwVfMvSSDa4C7RT4UzCG27Uhjx3YOPo15Fj6IayCD0WP6ijU7Tff
uQ+eNUQrIJ7kEq3RwUf8Gwy+SFOLlrBf1RqYAearwoJq3Qiqe+DUYFzO07mxuZPT
EaA1nXT4n86yWMZat8k6M7+brVSqXavcMZaHIAd1CWdFUfsWUjB/9lfpFiXVSFMN
apxFjFBbGJ4J/V2FHOgPfZntOkfdlUVriEMoltQxP8A6BKOTwHqxNLZeZFdAT+pU
WIKKfcgHefu1WvwOXdktfAX1Q4Fhreyp7R2yCuKj8ws9qacH2um6e0ru6nshXCjP
MKcgJ8F73wxMRLQ05BEmR1+HNfTyjw92mViP868sgni+wZyCY+M900JlLU6l1Qjh
NXwYOSdv/KpMzqOVtUp/wBg6xRvdd6tEjt4ElzDhsYqqgCB7J27VPM2Pth95xLh8
FYWWKiUvrDUsLYlKq59wRQNpcPK1QsKNHEPi3d0tUQSpr7FXk+8zNLQwrqpGQ14A
tsCCfX1aF0/hA2JYI+yniYCLBBXlaonKBsqF/7GUM1yjOfd1c+BixlIaMWxq52UW
3C4B+CUHXOi8wdiEotMWiLGsDnTc+i4NgGaCKgggkc89hUEaZeb9/2Nx+Mcie7pU
zCJpbtOfjAo+KxjBdgJ5IO//rI7+JzRVuaFJ6wis9L4YQKyPliL2YjCFMncpzVIv
eY4AjvgczvSGErd54zoe3pkuz0DSH4iE2IqTD5V8NIAxaeJzx1dkpTiy6irkpakm
3oSavNL1rsor44iJBAa1exZ38tZNkGhmlOe1GHItySIQxJvseMs1VOW4B17ZyY59
+tAVEug1lIL0Pf+Z1LpA7F4olgHBTXkPq//X2ZfPwmXwH5wScSKO742bPqDg94vB
NyVlGYzNXFtn+P071BbUZu09UXV1hSUxHZiRTaw8lQ2fQAqBQR3w7g67sI4IgFhZ
YnH79Bz8R5ek2OwifrQU7SwfPFE+t+CUc3+Qw5X5mrSgKz92gJl5LvXaWaPChENK
YNr5B6DY3cXI74RXYP/00z7KKxGVOjELwi/1AfAPY8we8TE5oYzUTs3Ns8RP9m+S
MGxonXow6gJohwHbl8knq5yrtc69WdH3nccOh7+c3wL94yBg3IgHRap+9L9ITKef
3P9q9foN2xb6nqINCTpIazIwm4WGJ4LMHnEnLG4YXFO048UA9JMFv6bHC4GD5RnU
JDZaOUwOFxcT19uVuUqsT8/ahtPRc3JXYxWYVuEWbSEQFDsOkZHyFxPBEiQHlx9b
7teraOG0aILxoLOpaDEBc339HxpoCBUxRSnxQum08GIgi5lwYJOroDLpGnGw+NRx
smKcg9rUa+/9i5k6wPSDq/DVemlc/w7PhYjgwPt3ABWVQrDeJ2XCGQxPnmTCJ0ku
fCVShKxumRWst4jm6IOcjcRaXIZcg/8zN5TBNI84jB+omUHEd3NjAFKqBeQxF8NJ
Ps8GoVoe0K9KAS3PmVbGEQvobyKSbLoXIVS2o2+z47PlBdkTp2j7xSxLQuROKG7j
TgqJOjlamQ2jootSWs7LNZoKGCtKhBXsUfn9cGP7OHkwmVro/yz5yiUAuSqm58nT
NhCu44krpK8MqHQ4OaPrbNXLxylN/QgPqOiBnTnsAW5Q1R5GuiDaacgEi776gRZ+
YKDJ7YRd1Ul+he9XpSlm0AzMpnnwl2RdFlnNhSEK8kS7WObuZe1SsgSQPDRC70Gd
prmkJZBDhBUX5EquQzrkhT5jnDyV0WetnDtCFfFRp94SYKmUY919fhXtaBcBlqnb
3RsTkXFA8uVIVAQWUN37FtYE8HG65sx/FJQ51LBOiodB0iFS0YEarrF8KHKWT+ya
1xoNeiPC0Of/Dhvp+OEuLpCjKkHCZTy9E2mArvwOKHWqPUpAZHPn4q5qimPBcYNI
r0/vvd5oOgX/xwPg1IElJ0YUejqwy5lR07FHBis2YPNFtCnXGpEcxQqgyshIWXHW
/Sjt5ZLitdUCBetyerN/+GXcV5EI+ahHLCAzvJ/VWPlQmOFi9UCo+UQ3CcJ6OB8D
+2/GA9XFLmwhJ1qS134N6KJbWhNLlTO10yMAyI5BTjmaYL0R0kJs10HxuNKGED6l
1sO6Y4qmTTdiy8n+SL8RVmpj2vaHU2lLCkIL0eihCMSWNbTSASPnEpztrxOCvR7d
f/5d2L8sfyjnN4yP7HZq359TvPdt6f5L8DmkJDPSt+nJf0CC6tzTc232NTo+Iwep
aqLY4ZsoZVFMoHkpoGj77O07yVmmmzS0gSsiEdFWVSR0ZnbxgUEb2rdYQzgBNGD9
TmohZYTKp8+x8XiF09wIF5Md1v15Bnhp+Gw0a2i46Wawmror6n0XchokhyjybEou
zR+RFsYQ0aaGFAbPVQib1NY5lw/YNEZ81C8eMVmSt07Wom8D0L/cgf9Wg+8ycgrr
JHlLVoLu3jjkYdFzaJE6ww8lcdW31yyZSVL5kghValOr+W47i1SaIL3dbILQDv5i
V61U8uUKUKEA8HQLuHdjUeGj2V965IgAfiRP5a9Gcunu6w8/ChecC9linrWq45jo
cGwPQyb7JS/BeqbdbTS5lmeLOj6olVa+0kc4DWMLsqIddzMXi82x0aUh5h9KxzxN
IHFrMjJSbNgZxATlnnQ2TYqYfi5YppYGMgt1eu721Xp4onEc2s9Dlrltu20EkArZ
IJBMC2g3INv3M77A2OHz8aXpl+IulBR78uDTCJE/J52sOhTnyvDJjfxmMXEtuyB1
vaA2fG7GaMweH1ZeiJIkDFDEw3J6TqJ4Hdqv6RO1WJHTepco2ulJ6RNKNWpPz6s4
qPjL7e1e3TsEx4tqgZsrvHEMh20ut8vNzm4zFYKzEZ6c/u9IPlqTPFDy7FF2MgDu
ZOIqW1xvlQA64MlnRZILRx03bRntT7DS0lMgvS4npABkLTPxvE/C5YhfKx5v0Hc8
xdMUVzixVpo8vu/yj+kbQ4+o6TbVoTsuCwKZ0NXZbj+CQvzmCI2ZD5z07Z0KCCJ2
y/QdknIisHAGkv6RcqcgrrdUi0pv7XVKmnN1Vc/q1J8J/kDLkEJo62USpCw770VU
nDHbdFICiMyhlByv0Sj0JlgWLVa7tr1wx/UYruIXbZkf63S99Mqp1aLj6JFHqjLd
WRYhuAQ36809EfVQsAKRGL1OW5LOsx8L4OP8tBGTmwe+D0A/AAl328WZuG83m8uc
E24cz9uGUg+vl5T6AzG5+6MM85onrR2/kNXYc/Rbdw7B3X1AXK7OWFqvcB0BujpG
vVzVTK5PrdM9iy6U5pBCXk3zLvmnbHQXaOOJFP5vlsJaNa/L847SLIJNBAHuMVue
3JtYmALYyWd0cnEu7bYxB+Sd19ob1O2nIqmQxjPtVIC7h8Rvirf8B5s/egLItx7P
lPup9P6tiGKuzXbz8eIMTMDkgYLT98LWKhtMgknZIXVaooclf4RfMHAgKXtlEWuk
pIsCPBLNWucI4OQFgq0D930IGnBksSNpdNDiLWFdig3lRWVS5a9e5GOEqO9JzvE0
sGQptw5l3asUZ31ifTkQvayQiskCS4LJRV7zAhz8r4ILAAIDzVxsmq3ClGu0tsVh
rLdneJJFRiCLSht/cdBWUTrzrGx4CzNU73NT8Kd1Ud1IfE8zeBUg6IeuNsL/v5mO
JBUOHgdOX4TZJjJZ8UACtH3O9tRnjxPZRajbh4WiTFKJDqCE+eDgQC/dooSzo6Ad
dpi76onfl7B4Fnk9K5tGv3TxjiFkgP56RkxV7demNle/J5vojhbw4bAubTIVdsyJ
7rte9aV179qIcYVu2styNqOJ59065O/x9qEuE+2H+wZQ0CwbZVBuUnrQ8oNz0UPj
zV+Lr+ZAc9LGSVlzXoC8lb3jUcL0wTw6By6Nz1tCUMmtrfpBxt0YGeMiB3ZG+Y4H
OOtczmyYt87eEuIMMvoUlVGtZ4tjJNfSD41VM6b3Oir7eC/K/slomuhA9DZoN+vA
eTkWAB0TSjsLG++HuL5IIQ4Q8PRCLL2KO8MtgQm9TZdzQA0rxl09Au3r8bjS7D08
JbfzGUTSNA3kGvwu1B10yeWPJcn+XVQVuW3Ge3TZS3rveFiQEEDocOzbTZKvLFHK
zgR24iONkpvcKe1pzhjTMjMKh0hP1WwyC9Vs9iVGJ/bU1jLopdJcAbh7LZNeFlth
AwoGpzt2TKqkTKTqMOswjscLvT2+EFZNQa7mpFiCR9ArbgBq8E7GIKZIH2FYne0d
MXEO3yuurVyOK7wtgnxTozx4IZoBO9QOQHqSK01fuVIwdm5MOSkHVajhuO2xrDX0
iuERRgd2JqXjIf8Sle4t4PX+MeqYTQY1n78MvCrYbOuOLUzf1dWtOZCjZ3ZVnyII
FZ4tMsjhui372PFKq3fBd62vrz8Qwj4RrT36fRW/+7DTUENE848ndxhJ0C43cBSf
Ad1vR7hBN4UUSPZcTYkDPV2KciAoTlrlwn0EFSEqbmTFTFeM8UnBKBlK6V7+y4dl
CQGz40jpnHG9nnwrbi9CZVqL705UFMfUl69CS8pK7YRlxvgmwm+3ZBWZ4HZBdWQ5
/Kl8p62DVVGIrd0A0yR9Fl2O8I02oqIIshRdLT/TDQnCW9fiYMbOf3AIQ6A4O+DR
IEHH00tRpmGMH1Lc/0gyrQDWJzlZOYekwv5Y0HxGL4EIMnODHafy5VL7txXO2ck5
+0SuLinn2UcaVE4pTBZkiJyZe1pcubBiJWc5KO/4Vftej5qK0eMMWLYwk3JwrJRS
ygTHOFGxQLXdF5ZaYm1wxvXHYhlOg36976pZDqBkE5e1J5sH/QY7iR+SF7oN3o+Q
m0OVPIdszYUIcqTXtxOQxQop3V9CYWNuVBpop9FMfiFDrMF1QnWV6boEvHJHSc2c
wAYIRvPk6XB17Ev4bZ+W275kvgN4kaAGM54FY0RcBZwASzDmbaS/Vqup1hhhgQ1n
44EAgHEUEkljc/58mJGcHqEEoRbF1mLbYfCmg696RvmmHCOqslY3lMpkvXTVeQxt
UR/RLs0qXkb5f1Tw8avsNJfhS3iE79SP/O5qnNji/cIRktj/v2KtPM9Rlf8zyEjA
d76HUMGVoys5170ogoPjlxGNXembhzCw/ZXq9xWlcWm1CmpHpETe36/TcgAGHFta
KsMC7uAwJH95U5mFx/zCX3m/g2Nu7RRvrrxbDhALw5kqX9HIBmJCE28vlURUwrAK
fzHl9GVS6WREuVw8kMDWua0+Wene9rBNRtZBI8V3mPD8sa8Xrpz0vkRiKLhgGi4S
hMuUcZ7I1XKMAXqLuPMzFuRAfo9BRZpeoimXBVPFAdLRR9uNreWwpykN0DYbcFz3
jE5KT/fhfRmvQlXAaPXRVO+t7JtA5lEOY6SN7kOu8xaiutqeSSans3aM9kZVFUXa
U+5E/l8WsWZf3iD7vzKPWCeVB39FerlzgSYBKDyfU6ApayVwI/nn9NGh1hOmCCvy
WAKNKxuBz8bGpZNqN9fX8liP8D0BwDsfQ3KJ5YNHZroeF6W0D/eLeinqzOdinsvw
co/j88P1zoBAqWdQIB2k/B633F1s7dOTJukcItxds/5Brej02OIeF03lpTfzTCQ9
eDGOCEoIOAmXHCEPYx3wkZex3uYODdVl11fBgCFAxPhiBT+OLvBAOU/hwLjijLTn
+Ha9z62414rrf1jnACBWyEGL7u3zyju7w/3aTrqihMkRF32WVvZyKKWuyhQt3/vD
CrJPaO6/ChY31oliRTfuduSk1CBQruTUUvAnF7cvcugyMoi+GC65P/4B0lDXHJSY
YLuteRX7NlvtmGucY5TSo+KtJEqQ1md5209p5lvwUFTYtMSgpUuLamgBFJcn+nPA
n0mrYOdnc7MDw4YuVDXdy37Ihtyxk+MJnOmPhA74itwOCMqLoJw2wSpMAq5Xo8Cp
CqPIZ+QmOG/OERcC7R7NADbMiAvJgqRBeifFEEASq/ifgTnGrGFYkH85KvKwxI6K
vzv0L7MkjDlriPwjcgta/L9IdQviefN18atT1sFadNdjoDZwO6kmtOSzCxXA1enW
rO75+qiyZWJPHgi0/C/G1uiagSKRzwz90m1RMQwuAttApwE8ckeDKVigKK9QATUx
C66H3Hw0k4oVatPIJ4a/+mEzPsCyqDvaKHnTey0vdFbmjUVM78HqtnKEXOsw/cl0
UJndYmg5efgtnXBUdxL1KD8sN+SpyUtzJZP2+gLCRudCpJ3/c6pwn2PZa6Zx6NG1
oMgsNLosP2wrupMw/EcSMpZcHKwHyIb8QXZ9BpT9jlh2r8uuzT2SnB8E09EHUu5/
HG5TICGn2N1ciy5NvDg+vAIsM891ys1mZOA5imqkLK6rOWGcz+Ysjug7vxn2S8S5
pNOwc5JrJcb0xe+GmtCiTgWyTNNeA5wxnzVEAe5zZ0ZkR2gbcG6ZkIF1i4tzCZgU
8g5yeQkYk0AJv5g659CKjjVyFtLB1axFyMbUn90ptUEjwJvONaOKvZY/ToGwfDHi
1q9Sk7/RWcxVp2hY5KCleB+KZMVQ5f0c3bkkenLnO8qzr9voZjzUt+577JNNAEnX
jasM7ACb7TnYGHnHbJe5Sgvd1A9hrIh/UWajLz5YpmNGvcnHYc55yusjnzC/bTVw
dCwOCBfBzpExcGPHIcB1FKmz1FEC4zYTN48Nbe7AwVKBphsEnxHScFIIkTqKURXX
I4w6qwHQnVEPeljmBDSlo5VA65HTIZWBJ+0VVTsqWU1IBlGeTTfljQdiQsPFjJEi
r7MmoAmLtbrILJOGE++WSMmsX4G1OnTZARIPl1yKE/wulHGWl5mGHlJJ29E8qyLr
f/eUtJeh9S571thRu2w4oR5esqTQNcQKKKq2U13/X4o5rmqx5ToRtZO2vY+D6fTK
2CNkoX4qTB/KWCZCCJHjfCC33w7LVfSGBl5bTuzb1jTaSrfNfK/AlzRqYz63OKry
Iw0mCX2sLtyv4wWgWopsy3iAJlDnfiPtHEdtEn/VoOJJMf8HC+6jk1PF77gs5U8s
xzgwVD/OAAaDAi6pM9QRGDdKU8X8EoooCJLQ+krBnegAsV6BjYsGRupBXli4hZcj
3+jWttQoobgDGY50LpT1Yp/z1djGauj9OIaJQAk9tsbZtOeeXrKkjQ2B3vJ18VfN
y8f2roUa1id3H2yIOMBc/AuYo7V9FZ8bjrMI0CKXUw3Jsioj1pV6HMbNVb99Lx7R
895ArDsbpGhpwbHYwJylMoqHAkdjsb0m983UVCZu6GLrXkGyM9nqYXK3jvZj4BvK
NoKfnZBImBIi59faaV18/23SESkw2fxXJXGaeXiL+Ki5xvjhsqvufYZTkm2Yuh6t
7qREFFiicQoX3gjW8nT/0hynnPlgmDFNI7xHzrmGlXaT58kVLqwWvRrHEJGfdxSL
MurLaOv3QFFs+HaNYc0iZKq3xzi1yxDduNlSHpYqC8BIiuZ/KiVGiFFP62OK/Y7x
aj8WR13uv23vRbf4Mw34iem4dRnvuENCm+jtcT5vvwj9LRQe1w0udJ0ZQun3euQt
IPB3yFXPMfCEVzezP6evMozXyrwkCWR1KJQo/LcuNy3v4SHVeFB4nxWAYOphHmwt
7AU/VSGDqUtkTSXdacEDq0x5chevwdJr9axY00Cvb+hNSoLbDgWEJSLG1EFHgjbY
Vd85AqBiZoVn727dV7dBK62Mu/m1OhO5mqhsTHGesVUhWewoMxfyByzD7UVkokVU
71H4kl8WvdEDKrXk0JoxE0dBUqEQmPsYca5VDNZvct+k8ey07lYjYFe7n3tOGHge
IvfiSkIfCuWaaxpGBIC1P60tKSQLFc8C4T5yv4J55qxKRUYlV2K/i/vv+ZiWaX5l
IuOMb9Vqf3W9J01D2m6caKMDCGte630ZvxMjE3dVMJo1evO0zFvO7i5rxRqTZYT5
3sp+4aQnAJwasMUwpGY4KalChjGO3RSF2ONzArXGvVyDiFgxxLKzvHA14/UD6q2t
0CYp3BGubH7+gRo3FnxMQTmLK1THDWRN11+QfyIu9fDXZriWniwBWdayOn+06W7g
OBF+pAS6O0dzUYb6NSxmGhOqhGHatlISPqXhpZup6BiUuC9eATFGFtDnCVAYW2EB
Omwmo4o4/BMwfrhIw2d5WCVvE3FIdqs+esndk1gWJ46mrvaF9XTtDGIs1+QPvZVk
4a6SNp1siaUzgAjutXAh9CMylVICwRXPdmCZTjHreWWBZdtZlYqjRrfG+TGN8Z2f
SxUNeaF26xe1rGvWnxqlAW7Sp5HBZZYWuWq0YnmPCCRAV+CFIzi7M0WFL91D00uT
dBY5h/EmvupGTu4cURH5tXiF9y1yfp6BsgOu3fntdyuDC3e4Um56w+MWr8y0Zv46
WpU+8rCvDo3fDfImv1Q2NDyyvttdaOjEjrUNpd7Hx1VNMzm7DhNFOyHOOEcNPheP
JwcHuAJnL4s1BuzT8iJnh4u5ZpJ/dnNgoRjH1l5Os62URl3WmNT6IYm6Gq7gF717
YFQLt8KwtJSjXSzEY9rTkaz+PpC39QsDexzsPB7BHCF+VOoKTskFiNe1XBY4W8tk
SiC9Am8gUzgl7pKeg3N9RL7v+hKUG+oP9dwCyXbkcuVM01AHdWzR5Bn/mu4qZVJL
/vfwfx2q3JUDposTyjTlngGvoqzJJpAPX+E1FWl+JtkF868EbDB2rei8Ik1wFUvX
7pY9msONW62qLmeyOfNcBOhwgUnIY3p7b81/QBV4MOWsE3F+xy8YdUgAkzkyzhUY
9ldFyQLolF2tuGxj9pVNQS6YYbeGhPQOrllKL7jaT3jBAZPE5G9+Q14Jk+sXy8kO
7tKs5B9he8SbNhBOMJFhM5RvhSjFjqDX6gixoViJFLk9xW3YeF1v+/Ry2fuWeJem
xeLooYc/P1qcsxIf/g17r4d0kfPfLOBKlNUTPBTG8mQ8++2F9kSnj0x1pjomkq3z
J4xlf/W/dS4Q/K5bqayY7dRXOuRoJvoxcPN5PNVG9stqm8b5NyBZ7HeMpAeWxd09
Fvfa4jpMyoCAYkov6jZQotbCqu7EYwzYBKGynx6BjfZ+r4UNezZCqsMulxAAG3tp
pD9NXROSJKR4FDzOKY9SQLY5ggmWQQwcFI1RYEZa6ZwJ00B/QcjvioCjs7RQV87b
SLvUMyM1isz591mO1GaLXhBPtztV7cxCaUfh6EyTPYObvfNd9T7pLFwRUWUcP7Yx
nezbpYfdNbEaDs7fjdZ5vk/A1cX1nMS/Fm3hnAbLm+hBz582+RVviCeLpQA91jsD
0Bsh2LbkSMse9NYaePDZQDsj5L/8p5izy1p/IcpS1JfNInmvYUM2i516LjlsdTEo
KVe9y7l124nBTWLKjy2WA4vezrGclWC95i6hE81PYQbfcWLKYEsrVFawTHM11vok
rn9+8nzZOe6mBvWyi/8LeL/175T4R2k7Q77G1Cp8TLNvAPbkL8m/o1kgYk0JfNpk
WU8QmJ58FTHfV5W6Xu6Jk3UpJ06RfS0CKWoou0XE2HCTJC8DbAPVC9qzJHDxvyrD
MQ78eS+DkCw5MaMussV/g5MNEJy0K4qtXDp0OHRNuhh5SzlyMtEqNAABdcwQ8XpO
/erHJWN+BXZvbHix8FEc05Hq+STZcD4/xXB371Mo15RLPjh2uSZ0rLQxa1f7daZe
tYFR2W6c1K6J5G0dmXGnS/Ovw8aHTKoshaja3BEJY2Ks4LN9X+wx7c7ESgZZJ3Nb
Y+mlnQeUUmptPR+bI+nHpgl7yGYqvl4JK/evU6uq6npQN1wCWgzGFn4Z19a5HSjT
cjLZsYH5KCRWE1t6qOm/STonVBdZpsPUEBb0yo10zEqZhkWW3MtogNC3xVoVQOV/
I95tAjSVym6yETQmfk227HxhT5RBmnzPSIplKc/S9re20NuOE+LzzVdWgt/kh2pK
V492Z5FyNW5D1FhIqexUlqObojanYc3r05OBm4GGZNcV4gEOfzVaI/CDq6qGE0Nr
QibH3XQhaq8y22GyUxIJLoKL/2LfXjouUEYyc8edybrohawBCTtIpiHTee8twfF/
aFleOIT0opj0gMEznt4AvB8eA8GbWOQtHFjkvYK2H2OywDmerFj1ZNC/awYf6RJp
SKxc2ZfR0X1eg0oyiayskemOpjDMl4dYAenikA+iyeD9lHcSJHEMGChxqwSOloTp
IYhWig/k024x32zbbWbgDkwBRJv+Z6JJyl3nqTPwUxuGGEDd9NdQI3oLmp8iu2b6
QpQTMgpfK++aoNeqeXSrD4MT0dHqwGKITuFHjn6EH1weyGKBEtLNdeGqcbyFmRlX
h3ZuRvHGmsKgEthZovRKMW7z2uynGg6I/CsFQuckkFV7eGZBscCpb8fr8Bp+VgTi
pB0eap4DXUUjCl/8ADwusFji485zv5JbM6HuSDPaExMjPO38LNqwmbt9fBdH8aXj
2CVbCKk9XbSi5ji+UJu8RFjmzseHYPi84KZXNIVtat5JkQVn0DcODR7jLFGptLbB
UZJ4gUN7xFV+24hz0XXdvnfshT+jdgpd2D+YHFcXbzaGGkw1I9Z8Zl2dFKW8U/BS
Z3IfmcAx8JkPaJe0e1N3fMFYtDlj8RNsEzNa4DEmRJXyRpBPpwPZxO2poW6zlOH1
MnZtK+169BtVBEm8w+m5hnG86sx8v+/gSMgH/tLj3kQoXg86hT+ANjltHwfreFFD
s2YyPPTYHa87l2BmhHzN56j47Po9/ZJQ3Z7GRK4Ve3NGne0LhoRs6UAlhjZNwsTp
Y27lUC43NNVE4dFw02qNLoZd6JmjthGLGDS4s6uJYUvvcgzbhjgHo5qaqELq9V7A
DMz+rFEuEWlG6k4AK5PXOI259POB7J+AULuiHRtylrc9rvUtMx3MtG6kXfF7k+gX
In1U3krnCnG0YIHPnKoZGQdmHh2s+X+S/ZF83wBZBypJSrfpM77AClikju9qdt+p
2np4jcXupRXzQBWyIQytXlnZmEhxp8T5D2IpE9Ir0CB0CZ1C4TgrEo9EALMag6Vg
eoFSiCG+tMAPzVJbC5o+UJXdl5RHXoD3112Cdg8bRibHGY7IOedR9U6Jrff+XacX
/6QzgUF3K9d1uQAqud7nUbg67Yphayb5JZZNN8DzqHOrNsK1PTnRy8Byu7AmjWFx
kEljyzDKtwf/sZdbUhTW4DeD6TkjYU7sLBzulFOpoYR+CxQVylb/5Y7y4C9laYTr
EWNfEkNc9qI/WUlzt1i4o1tZJsay8jvLwYGUUcgUk8WO0XVPLFDDf4Qpa1ZW1Wq0
i+SHBaTzNq66gptNNO25eKsnAk/vYa58B2TFeUh1D0Mtz5hu4QW2fBTAVpF+wQ31
t7QdF3si5wA/KL/LYqFtP0RYZnn7z/2QmeuL3NLFxyLKEKRTQbz5rCiDac/CqOjI
FTQRR/R/ipEO7dBgCD0+fkjjziPtnMkBGNfQgjNdP0Fe8Y951iEJ16W0coHIcMCL
oNAKVGxqxVYilMXYCMMe5EnkCFKUp6SAGHxZpiROdqR3OPQGPm0QwefPqTnmgcGI
SpGmTaIlcI1gJpGr4F/IJ2vw0mF2eUv0zWvcP1uthUCTGlGd8P30vS8VURYcSiwI
4Mz8+BA9U8TPRJOdptY+c9fz2LTHYl+bDWW/cyCryrNPI57amvmQR1X6SDpZFyPO
CbkPftsUXPA39rRdHhrSjSCQOAR8dJDxVkn4Q2r1K0xHaW/ULM3iC5ek+ZItXpzn
8qnAJyTT2pGKMmJOAppXGi4+hXmFwshMYjpmez3snF1ZVPGGk8D/rhegD2uVGAcV
XR6OgXayItG4IUnygADSFinIYXFjh6YB1aviC7cpgSSaYFcNQi/QRnN2xIN52+fi
v0DN+FbqxxGOAz/6VUNtAi8HSltZC77UqQItxw+SBSCvdEGNVK0/swugu23kkYMQ
r+ke1iomi7ol3jnsMO533SJvhtBr+FrnGWhTB3hANhYVNg0UnFkeNh2tpv0FMJm4
09lzgz1Gv+AWydpsPX1fhYe0Oi8TwaVOBUhkx06xfNbOGsdiM3C78vLWyrjTj1+w
gXJDRj5Q5Vk76NseMA5V6LRxdrYcoEFl8DZ0lhmLo2qBNmAt3mNOuC2fN8IYNJNL
ZfLRTOeqo0Av3LNYKhs/6simdbqPVtdQLUreey8IO/Hk0LAkUJdYRdCn3OV0h4jv
a4vzDpBjWfl8eF8ZGg6y3Z4JPwbJjnMLZma8hqcE+S2i+16I7VV6ibMj527JV2cY
6F8wLOt2T3cwzWt5r4zRmAO5OKWdCDiZKFsxgAOSGXILIwIkiJ4Z372fSsNTl+6u
7g3oz5iW0SKCduz3vBLuwfhoXcG0/Yor5KsvEG/ZOycUvU1X4Ck3RJHSq0bRclaI
tKAxQ8FJpyyuCw10jOkD5I+T5yiO+Fd89UzZnjHqtD63Ggc8Psm5sILsuVM4qrBr
IcASURt8HRSjOkv0M9c5kf4JOykQ2AQBUFaZsOqIPnIbAoq0Bm6DDxEHBB47NKwI
bsMvQOex6Z6wYBIoUcL1NSIjP9wt8k4sKo9Unxhqhy8pjLWI2wO7ifgTHK10McRw
K43B4Dc1Nlz7ul26WuQ418NwQc51JozlJynWa3v3cGDwBbDHqpwsorRvnIFwjVFN
+44e4r7TKOlr0q7G5esg0v+8NYaWII9zdGRljUht6GGHCyvSJ7y4F+YWuu9Iej75
VKKMbDcghUlIWyyH7ruxxs/W4pPSfq7lsKTsAUAm5YZC5sV9BZhwVCt0TM/0oB5J
OE+qwX1DfCBG3SHDuvw7ZLraMKQkZwKXp6irFNYFdSprVyFXw1WVMeA5rtDnTOB4
KX7/GBnCSu5pR4had4fUQVwLQkMAgoPJ8iKXRh4+yVmOU7iqOoWmUer4K2uNVU7E
DSD6F70OMO0AqzMJVvkyMDcxgrb3Frrfgh6XGUeHVw8g0m96kR7twsCLwsh+rp4m
p6IsSqK9ZjH7vixkIKyZPKJwb82M1WNDVDo6WKji57Rh5JUwn29/G4vK8/nLYD/H
5z/5w6d8T1g28byK+a4Pw/lrmLo7q9xc5/v/RF7LXQkagChUX0NPJ58g+bjEG1zf
EGPsrG4poP/B6XEg/tiKieLk2TmQSNny+eAnoli/BDonzzmWFh90MaAvtGiM3TMx
DpWDtXfyHe2BCCsGWnGJgj6fnxCs7xLKVFyQ/NaoceAtQdOv6DmLBQ3241qYIwpP
W7Uv6P6MP6c6ny6BWl/TTCm5D5ijY4PYJWk3PbAWRo972a+geo0BLwPi/4qRrTp9
0twnXuLKShTyffkstvjW0Lyw2ir7QvTbqy0wE5zvaedNssbStEFUUFlNj4h1rqF6
aBl9eRdM3EZ9wloDOKX2xFteuc8UKFS1u8b72sK9eTRdWFPy0VXV0tWTE0FxLxuK
SlgaqBqDa325Ozd/S85b56YNUFU19sa3MLG1YVXYPRJmRN7tolrX4/OsY84exUGM
DIou0xnAKsgl1cfX/50RQ/ARDjM024IbBlQRET+rIXZlkS39keJjuWfNHQGuhAQF
UJPb9C7oanevKfPPFwyixBjZ+LHjuNwOiam2K4hmKxxJ5cmvg8t2neENc4A1KxZT
+i9XUHj9Xu+7dN2EhKJR9RlS9BCdyYfI41Qc0XMCTKMKFaHt3Hn8rwF68LQ7Dzwb
sqThwHfDWAeO6UymYHIHRn/OEdzl/zC4IDyNO00KTG5G2R40DdrzQtAlmt4TZ00x
S2VqI7U8S0B1QWAnBLEzagYmpYl84WD+w2E/Wk81cuz2Xh2bup6HiFoURKZlX4Lo
PA/2J0wmE21KDWdzPCH5+WpY9a903GyDiVwaMsgQcGtOt135VCxl7OJGIx9+zIyf
cri7O/Br6H334aaNwFzMt78VOoc3YEkNlZSMWI4Cwx9UUp909GpTTtGy8kUeenyG
GTqA1Cy2OYLClre25uHIaXN+p65PZkna0GLnzlA9Iv6RPHGKEqrclLNeVNQSnr5Y
70yn/wrgCXp9n0FePWzrbICcOtL/+AL3iMPxltTu2xfM6mTqzc+HnH4xdbZtoMJv
aR+Qujy7F6nHccmdhGABUZGlK8rDS/WanVwhp5me3DgXskgx/2H5KHVd2k2zmlrz
eqhe/4O2HyYkQhTToHaF+yvzvtzy7xXkTRBBDwU+dtAPe9mNMk/NjXy47kByMAFI
eQgST98fyHZf+Wlj7Ee0dIuDaB08cB5HHT5O7OoCyxU73BcuFFRkseJ44FNFR2aS
5P+NI7pffVs+fOmq7rAL7Ut9fec701Ds8gayKBb3YuE33TAp4yyPMnSv55QyQ0Vv
v/Rw/t3ClLKwFkjnYfd1ddIakcvCXIN8srN4MEnp75GQSn5fz2Nhga+4Kq/bQ5af
g4WDYkEKck+lxW+Li0AcBqwC8qMZ6pcj0rcQ6nlOGhC7R0jlBCSU5aHX7ifO+8Ii
LGGYtJjn3uz+bWgYMq8nXXiU6+IQI2l6tigPkuJ6eQgnc/xF43Wjbh+47qpmYndl
d212LXjqU0mA9djZcX0OPF2a/Jo3lRB1l2WxUjG+c/oh6LOvD1uAhHsL8VaU5361
R69Y+y47ZFc2bAhTQHTj9UPQWh4tx6r9pviZdTn9sI7edQwe+Nfh/OnEypVFOgMs
C9HSCu44EbzzuiyQauo7UVujvk570+qNTYrKY/eOM9S3HuuDlDFNsGlK0HDx9/7Q
iCeJ3JL4YMOf2dG0UTyRsBJkCrJSHJgGfO1EKrux9MMPbVW6US7iwgk5+Ag844O0
n69nKOTrcdPWn2UdgjAlQeKalFvGXPKPWKm6ZhPzNWi9xqjwB/ubDl5Iv9EzNBPh
3EtLoe4UBVbqbkcFSaPRl+b2v6Ko47NLeuhwV3bs5PKuznAuybOe9YRu5lpRtC2e
+P4AheCb0oBA/1C9r+1iwCePAYvyY6nq0w5eJdafh5MvVDNbSzJwOXKXMDV9pveg
ppm4TluyBjMR1yjj3j+hMit8+idw1W8m9kYGbzahsxeJumE0UVvPCbMoUgFOB4vG
iUapfjz8HhMqabw0vlAkYfA8G+mazHXT7AqPvcqu0WQ3opkm2uLKiYjO0Wgt5WX0
5bL4q0MRYssHFEotpJE8etYX2R0m7lnLXg1UWfdE4BibDADsAgLY+2dG7IynOXuM
PCwJ9OAyv5k8wCIC9b0vPXtLhk7DGgFqOy3lc88YHNsiUyaEjm1ik/D2Y0mFLu9K
DBxLvdq0oWGv4GI7DYCLgDp4jiOXTq6Y8/8WJL2h9dvrAS40vb/9qSROO9FNWWi9
i/e/L7PoY5wLck+t98Srlix3+srvf6qcs0yw/LVSAQusWCiABctLUme2veRXx441
sHum6Pxs/s9lObqpGyaK5/vM0jnXre4UZQdrX2nsJa0UzbKQFK8DBlHm1x/LJ7Tn
2J8aC8FCIWD8zejkODsopTf8rlrU6O7ZYVQQmH2dhhN/QTz4tsLdu078ZkTPAcmp
i/llTt2W6USVAAVR6YlTgKKI59zZW1liBuFOWfBL+K3vftW/ePsjFqSUaIDV3/oP
Li6JxhYc5FPG63ijP/KFwBA5idaFnv3TAMKsWXw8Z+yfWrYfl8tBmCjdTQiY8FLB
CG1uaXgEaJp41Csn1T7BUQvLZBSKIS8EbiumyNV57rfKOoqujlLnQW3fsx6S6QKN
95YXtX/vVEJBJgNgtd0OF6zrz44iVKiHPwpC2yTG92xfMIHoZw8zZtli9CEFramy
O3NLS5TDbqbwkAMo/1HEjfSABdbOL+cUNlcBtLlgq1qIPXij9O+8k2DsV4Afl5kd
HDp371v53ncmy6MCPip5kykR7PIlyaPH5sZ4kb6pO9agbMztpxBHozURA4CTv2Qa
NIOw62zkcvmMtdlC0zbdmrJxAAltF5o0b0bNxlQbmUzLrwKq+0znHocx6BQV/WOP
ysQct8VebeQepHa3loemqtzeUb8Zskgv5QFUx0dFJNA4F8QmPtzavLH5UFam6AkY
wauJ7vUCxyu20T5Q05NxtWqNO0FfPRN2qbQubLDv40DIN76OC9D6iRTC4spH6Y00
DxIGmkiFrPdZEe6+v073YQdvNGM5phmGAEsueJ8GOAA1v2z5CMjsfWE9iXrkNj1J
Y4Z2FoZwbR9QNu3duLALoeOK+kdT4zF2VzdyEnbB1t+iyRTq1sZqgFYK3NYwewj9
Z8ic64U6p6tNY6BDwnbzWxRjXQoL39FHS6K9BwiWh8KIffzRjjYQPsCNvGLUF2hk
2Xr9HwmaRnTuhJTt1+X0yg0ACDi3hH9VsrdvUi6S6ebK3/kwsEZSTQkk90kiG30W
SdSKjtuQP1QR99Mvr0TW2Cgdi5VeVmaS+2aTU3gWUm+oIbzQw1qyxyh+ncD7au51
+Qu8Yt9nSZ9AgIfJ9lWI3WL7B1l7OvTEvvWzubcG5/GUAEfYV7ChDWtounTKB2jW
SrfK5JLkPWLrqMyVNkfo7z7SQPbiaKckw2hfV5dIxauFkmCueS3nHqJ44digPHrw
QHpKz0BZwQQoB5pMNzHb4ODpeG0W1DSj0NbwuBhQM5mCbMx9ATt5PqTCTH+P1iLf
zr7ZouqqPzoKgE7UimRVsTgCM1JI84Pcq4rl7qXbUuNeIsH34Q4QBdvlYj4STcxn
5aIzvMeTFgf+0OEYx5rRidrBfCWHno3NtJXZ37XjbHGcytfdXj9Hsd5pBb03yeNa
Zw5ceIcRC4k9kZs9y0/FREEm6GsB6GhL9I3X0AR5u3Y950LbWifYjFB88WYjgIpf
3Y7hX2iGLZjcq/UDdqkYGBOv4vfG2xU6Z0tKWCcmCE57aA4SB4MEI0IpUX7MpDqG
0h7mQmyjWI/ImSLLZ5UEm624d2Xr9KdxV5KKccQNWBOL5k37VZmEjLEpxvvAEB6o
C7pH9sTddLVtZEuweUwC7hQU+yGSmgOQZcn4cI9kwQqe/yX1RC4Whk9Yly1tW+Sr
clPgUNCNjJlm69sx7tcxQ1R5T5p2pFWR9beTtUbBk0pPyMHhKCLi9UltB5Cbz2II
5zi6LQPtWCONuYO/JsV9qtCRoqcnnuhGoZW4hahOV/aissxTPtP9CL5rcMnGDykO
eBSgEcc8OVyiF9tKvu/kGFrp9lyeGv8aAxf1jwOWrWpA19UeqhDEBbnoQkh8cfO1
5BU0oMx0opVNM+2gnyB9XV4gdUQlU8M/uzJz4hHVLEWF8UCnGz2p6yuQbaqfhQZn
lOrsMGL6Y5pFxOSMHzmkzvrXAhwWRqBEcsdPwmfU9Hgctc7Cf8t50oHpf1Oy2Adl
hFDk+2ZCRu/ZkZuRnT7uQw4eFasEJ77lJjIYYJ4hB965LE9vy47S87GEHotSUQei
/cAzZWbZB58QoVzpJqKkQY+kjwbfJQE/LpoOZ2mBl05Z38JVliaHEfj7w08/toi5
QjxpgtCZxgTrKr6jCvhvHR770+9U+PE7J1IwXeVLjYwIfTDds6gOVzTXBtICo3nk
b+qh3zNV7Hivkgt8A4U7LfxGKmxccr7bKF0J/iuxYlBL50H7pn+0GpdSgLf3Ycej
ycW7UvpmGrtTOLQCP7MOuSldIRy4lZduYLF1kxBj+vx29oCPCEiS7gJvlHhxx+on
7SOSqvkh0+CULmXCMD+HDVgrsdQqb8bXPSoEip62AUWHHtVrwJM4stf00gG6PkyD
QZL3ZdzdF1oXLhw4KOpTljtOshJAoimd2XFIKZ+/lpNiqXEb978oDg7a5Bm3/7YG
IO0UzE+TMV3l2KiFOo1AvfwfPvxNULL6ZM49wbEcb23gOfSokdE294DDiG9Xwx5K
gzsNKnGi6rVBi1Qsthe0YLTHr0IOXD6hEAGGUmkrt2eMFaULHpnv8JRRr3OU3PPx
hdiVtXVX8x5xF2tJD/o1VrVF8S3IEKJwpqKkpPfkJpRXXvp+yRTlSyAHt2dEy4iR
JtiC2rdYez/PNi6IMhbfBSk5ukpha6D3+D3Zd0+RLZ52viXSB2HirB/ppflJTE3u
uHtOsgcX+EPobs9CwdLF4AeIu7cajfeFHqv/V3SSx5pA0J5lkO6cMKgT4FIhW8gv
GhIFMaS4pwZmwQAI8khJ9bLobW7pSwVclxPDH4bixZJ9ZVAiB+DnTueXfW3XgGmF
DuSjOojz6imc1fvniOUuzatRg+EBhTflPscD9cJW1luuMgthovPO/Ca4HehB1+I9
ePRG2uTQRrWzd8/RKyzrmffMjEbXSskFKADTkDesVPd0iY7O1RWS91FoaZdRxkFo
pterKiNjdsWxFpBo2SuuQ6QTuKXTwu8vpnqt7niIVWzAtrRr7FesaqeTyOBAcRCp
u8RdtKk4Wl1KJj31qM/PVPscZ4ML1VS3l+BIvb1gQuPoWqE+Xy3pXL8srlphGN3M
qOS2ui/aMzXkua9X2EkWvb64YxCJg5l5+gtScS469RKfBvRDWtW7qlqKujF9rYsp
Z93uP3ow0/md3XzpCiUcE0fo8D8rghNQq7LePKQy29cVdQzWeewDP9ea35Cz3uuD
IHLErhp/Qay/n0khGbckrpr1VOlUcMSSye2qMJ7xzNMh3lpzap9v2ESAk/WR35O1
v1ceHhtQLUZiKOpwfgFe/lTIzs725LP2vUxQ2FVB4+NR1DpD8Re08LeQZ8b7V3hd
ZU9OgoPVhVPeCKyvJKT1pyzOtPJSlBfhpPmcYBnP6dnHtYnFmvN2ijgmlcyqtokc
E4R4eqzppgyuwkxNZ8EaNtV5BTgmYbyJOFYPqlIU16K/t4PnPNoSJtcgNq/GdDAN
X7b8KvcF42NebqzF9vfvwMyhCOCnJ7HO7CoiBzdtXBSV5ecuU2c95hiF0XmlSZaq
khERxIvvRakJgoiPGdpc2zmKFVjY57nd0OZdqrWC3Z7RO56hqb+58j+7HFS6Ja2v
UC+AfeEsOw93b/nki/NiH56z0HMJgfwk9knB+PvDR18k3YBPH3r2UD0/jP1293yo
kAdTKeIYaiusy1LEuW0jMu7n2xM5tMMjceKgu1OhhwGpIN1VkVR/qaNll8gHU/MC
fxzR7hXWzduM6tMqZq3PImin/8DuBq2brSVzi6LyhYrIJ0A9b+pysygksplKCV3w
ACP33+r6eQCWsilH4hGP8x0H+gQgL1z/xNtc0pfX5cQgoVwNFXc1sKAmCQMRfmi1
xPHE73AdXnFJxpyNkI3pwCMrRV2nu88WLmaTQ7p0pAoVmUq0lo6IOhp09nSrjmXJ
udOiFClkHf1ZCyudCRoqLhIm3Z75FD5kF0IczqdVsCszU/8hSYLbNdHJq3+8R9tV
8uLKLKyeIZTtpi8GTa+3qjBINxderqyctQxess8cIoZLlfAj8JRQQcOW7kU1SLpM
8THBlhzUkQivBj/801dv/kpU0sW61s0WrBG1ww9tc0gyGFN36WgcTDuArFxdzr5L
xn/C9WpCny7WgQBj4JlcBw8S1674XIlSze/GTu1SrJ+uQXMgHI1Gq1bJVuFCCHTb
tnxlM3wEtstkg2z3WEAwL+0f0BDbH2cfBqn/+iYGYSVujNj0lO4yPI07Wz2tH8h9
vcoVeKl6ERJ0s2kJDHRfq8Oac2ZhoHDwIFs88aBHdub9WpSCjc4B0fcWYIZA6hLD
k3LaQoyhFYzlsYwz6wkIgYiJV4Hbui1LzEutUp8kSEHFN7e4o6q0/EZ93n9qQtbO
oFJpvA5X1KlE8xfS+iz/boPU+FUb0d+KroEwIjv0IaQmC6s03uHJiZ3QvNSYvu6t
E860NAizyWoBlpg9pE8lDRYMsXqB2Lp3lgour+llPVnlHV22Q/HQQZmgsU0ieuhh
pv0Gy35UpC5Fv1O7t+csuFHl/Y/k5LkF9MCfObmHJHaah3x/A9HYDQBTh6jS16zl
wsHpRRHd1RszUa+M8ehMnelnqhGUuoZi6zA0eRMDz5Y+VPNdQVL1DmI5Hn28mRqp
paVhJbDyJ4FHoPFjJyeDEAwhlVydvlo5178tGsrc1NN2RTM1XICphnGyy9tcFDFe
UNmqS6TKw+7AP5dB6do9fYKLyS/sYIT2eaxSU+HnN3oAArHzJwsLbZDLxFfac0yl
ckHM75xQGwAe/QYiLj5W0a0SU7qaRgA+S2OhaQewKoJ/FjBhY4ERia3n1XSLJLaK
W4g12qcIGw6EOpWycsrq9DPCHVeq/VqZPiOpLaoZT2w6FJWpIIm2Kwm0oJri/BQA
curtaN+JMdI4GwB6RmCtBEgczVhVh1WedKCbFx2Dx2nWOlC+Lg//omaLz4m4m7VI
1ewZbLi5G4tDil9S3MLwupViFfyy3y7fzTZxDQ597y9bsWM6lkbsflEDFQPRAIGA
OEZ21mBNnmIX4AK3lNKIUev6ErkHtnLxXUyOhgSVpK5jE5Al+obh+PgUAs9vZ5uq
jbRJtgR8MqrF5rf6i8+Qi91mfg2j1U3vsTiqRkl3wSV5XfjFKQZIXSoaZSBUCj9z
G4XGMwdWL+Wv8X8tAAHQmGmfOOv9JZuljkTekP9LiASrsDC/NNGPQsd6u8cDeSje
DEuR59Fl5tQj7ZG1pYJGz5qiaHjq9tlNQvvchYVlkzGbXbzYE8OaDJHsTUO3ESiU
ZtezZdHJ4AyZMPRgO5mLhi/dTxBjh9DmgUAFZTgf8HHi/lrIKWRq3ooKTap3UCRN
FTjeFaJqvY4llLx+OrEH+RUyxPY2YB9rgkmoRTK025K+/IT2hzIQgokiH2QpTdXU
mW9EqDKV3Z5r3WaL0DKQMCQrGXfa+/WT77l9mWzRGcf2Jqt1ZWfGXrY1k7QAmNjM
aYWelGYd8Yfm3qh683q+WUUNWmY01mmm7eUcJbI4XqVJvq8GrgR03+3n0U5II/QS
WIW/Ea7fNVQQ4rAgR4ubI/bKPN8xD9FOZS72yNspx49lmFGdNCcKdV7oCCNnE/wI
OeL4HYTP0qrf9Olkq9Fnl43iQIXHL3JPXKe2Lh9Zaq3cbOKRwSLv95j7GR8nnFEG
CnaUeWYEdms0g4Xugv8/Rd86n5/Y1netrevbuk6022MO5r31JAnJPHvOevmc01y6
xeG7I4IKNTlWWRFDNN8wYulRpjnGqVislxlSrcRb+10/6yftGpe4rro1ODLbiI+D
gTTeaFZiPyxiXkozZ5GJdmSr2sNVUhPA2prynPbO39GdBMsSgJHvZK7u0n0PeqHS
3X4W1VWwqfbSyLWrwNC+h0jqv3rjaC55Q2yCHCn2KLPvz6sWFEtftaiUjjAD8xAZ
n2RSXcUsQZzCqO6D0cXT9qRG44Z18m38FGEn+S9hP9/ry5eAImO6MZWjPg17eUKp
NThHqDx3IDsj+oazLhPQmRLxe75CmqRkYCCH3tP3agDhTGbdRBrYfQ779jU1KMRI
nrkIh+8E7PDa7SGOSE9WCfQWyo1OV7l+Oe69k298Cu8jVCswUdrU1XDbUAP8wGNj
+SsdzATfiG8XJTEN6/rpypyPtCm5cK8HG6prO34WV7++t5NkvBWfXV9R7c7EnUAt
zMvJePIVBz4KDid8qQk0feBQqyMBGR7Y4V0C78PoeA09N6ZyibSjCXbQRO6YmBMF
AnveiXMCyaMN5SYC1/eMbjfe6NL1yud+r3Gnfx0Zi3Ee5WoUFX8wPpwmcT/E4zmm
DBovJO7wJV796Z5wyWkIkNuPvI28dK+bHTOAkW52imwILiXBHS0HmkncT93bcVa3
073NvBtFzNofDXcKslC8Thy7GJtIxZ19sVaXANiLvFRM8gzfhXcYnhZNX6pqU1Dg
AgoziNE/lkub7U6ZT+iDsmyl9RIrfIcTaKvfKFVFEIBcqNcdvLHj0J2KSYmp6iMy
oOyg5ka9jhEXOH0SzW/yOyYv+rMWNj7wiI8oROZPCakbPKoMc6HBoMjlHvDPFisJ
AUqw5kCpc9tGaROibpLNXRK5BlmcmBjjBOk7x6GdkO2pDpvI5FjnGz+QEtA6ydCB
oH2LKyehIA+JAoj8pLsZz1ObJScjH7HBWNmyR1eS4vDuWnBOy1OCRW0hY6L7JNLr
BTQwBU2iJPHI6/HlzxueiG/g1mBeLXihR9vM+92iQAJkTqddMo6FY1HU324Cc3D9
z20XltLIVbB0nxF0qTKh0oJ87s4fs43WVMy4tg2abRc0jH5rCeVIgKuZIWpSRXnz
wbAiPMzLGqRRH76Kj0rw1o3LSMax9x8nbbtH+7vttXG8UOoRjh2GYxpoR2zgEvtd
ijQQypVNZs3C+hT53yIlKhJ3Tc39koVCO1D4gXkhbtAUaCmvv7nqRf0dSyj2p4Dn
y/9Vp81afY9O+ay67GOg4JOSCVIOQ/6g4Wj4OoCDPxzHUy5AYMRX0caeV8e64Ci7
hsLcEWZiofP1DYs13woMTIHS/ONdKO4uIxWDAIZPj31qMN9w6Ryjg87XZTBkApqe
6UAlAygIQKscdph/GGKtLvnhy3U6rXalfaCJaCre05w2WHyPogwRnDogMuiOh7rp
eQ3t5FbNJ5O5D5yu3t6qtoV86s9LkdjjfCZFW6kaf1KCPpYVVSY3Jc5U9W67MpGl
XzVYRUyBQiYKk+eMVUgzHJzwQdS2X4uVyH9aH36FIgpYKpbTzIOf3sjS4DuRVfpn
yDtvUrpWT1401ueQN5BeY3ODO6h0Nw8pYxGTeq9olIkY5y7ACmCtPcDdN1s99IKW
yFlsQu2KZ0P27aMdzjjyrAx/t2AkmGfI4HS6BaabPOhGODZ3oa6AazN+o4UkBXGe
3+MLC7DFTkiDTU1rtYKHvOhFUE0JkHhPa/AvHfE84oA561ajb5VBce88pXXSDE8M
PQjtzDASXZn3ptwwXbptBF09xQQaZ/jBNYDe3qzVma/MTH+Vdxts8pdyGzWspNoT
Xnd9JL1RU6T2vARtx1FPklDKbvgQ1Cn70QL7d8OXz25pMMD9SDmOBMn+vxnEvLeM
f94TNLiEOFSqaWi7vLvWzLsQ90KICVEG2JGXfhZSqJPYh0A2KJz9sl6JPLN5oa9G
KfeHUPx14KO/L1FlYKrmMjOnwQeN9kW9CsLjHGwIhHZA3/Q9oaaw8Y44Z2/AfYzd
RVVktrUa+101oH0Y8dshTLgqIKcAn/lBZahHZ2cNxx3hMZUkxQoGAJrqX2hmNAvF
YM3JTQUIiqlWYHYD13DQ0oKxLZva2e0HAs67t/aZ0PQffJSzRoVOOvUVGcwmtuqJ
SgmyzDRWQ5MT2DIjaO19hOR2M7gGVd2tdUuQZ12OJad1OSpI/Q5hcUVI38tiwiJr
nw10MQKqiKI1VN/NsDXs8mh0ddqJLrJyJWxvpxHvIcZRTzqhQLS/fvfVpF/Kx4Xn
F8j/oarMsi1PUUefwanXqqNMrLpVm2ZkShRwSyOlyjzqdVSBoh0OkLEo2a+nUR8y
SwpGyLS/o9OugbKtyRd4tsH5YtF5dFuuVPnqou2yst/ZcshHhDewYRyJyRvOGMAu
cEfOoHdBmLm3aobEUKUBkjejZy7dO+8Em5q+auSNsO4kyNe/n9HNEIBNcaX/71Ps
DYOgl+eou+0baYeBblPfpogocWo71kNNsmuThUDoFpecKsqRAreemyQD9k78om7I
tE9GW4GsddJ2KA4kaQm8TbbWAH2/6T2NcuUla5b/2ix4o8/5utpuNcaXtdpGHqQE
nfzQLF1LKXtCrsGqC1+eQe5L/pE61jqaBWHppsHct2tgRtk3uQsYB4S7CCYr9k3g
557b4DKn/RCe0XrjJobX04JMSM9IAqgWAptpL1kukEGL5vZTTGaHHQLT++aQspBl
1NNMKTXO/z5Ifp6OD/lUx5e/6KK506mTnkUyzVkOitW6t9bBcJ5mG71M8Wv3MpY5
JV1/B51igIDR+gHqXMYACCpLM6f+VtSaSmnbExbhn36KgWy4k77iXlhOVZzK4qoi
dt10twZRhwUgUueMr2TIDhErRoRbyNMjaLOQeZgdKkELCAlKSzXWb0UER7TFhwOU
HtY7luP4FV+6w/S8ksIlStqbAdHoakjpVkxKM+4zhQ4sebpiPK1a+A//lBMatCsA
jA7uCDlgR+LQbmnhiZHbdhm6AmBtKgPVzvJ7GaDv5hPMKO+lwTeqQ5Ziao9BxioE
R2xP2YRmzv1Z0uHeJ1iOfP9QE9OKxYoye7PNdoDNCwNxtUxSVxkzdTKcM6Y28B4l
L+g5rghHmJjDr09FpdEmxtvJaMCo3GcvjDn98UWjFElZvNpgfULg8lYZDXpCvNGy
4vWBqS7pGw7yYIzWP5gYznzkuWdkS2GS5HPBHd9WpzTlPt7eJnwF7KUWLHJdf8m2
+0nXxCGQuC1fKwpqhfmv8uTIyYviwy0EdFXKF1+oH6SBIouEfXqwP3wyB02nqN8A
4nzAUw06XEnySyCzt9DtRPimMi+lw5mClIlDWsqf6ab9rTYw3SBVdxhQnA8iriuY
P48ab5ACyroF1PiLQkwwC2oO1XwtCq+it4cOUFmUtiEK26j7tDJDYfshCjZnuRvp
wxLbDIwhRndMpyz0G/1g754LXzUw8JQrTDYIjQwzyUMbV2ooD8jkaBC9BoNuHa36
e0RGaplzdO4Ma95Z3kri4mCytZqC3uiR7hB+eZnI6eJDRqBuWjhrj9ZTCFeV0/Wb
1OEerSVmH6vbHPutgBh8Iyl/AfCI2WBQP3sw/5kvVixDovba/2y2IiBWpjQe5EyC
GQy0YkObx/6wWdrgS0bNrK7XV1HnQ8Glp8KyxYIPkx3gL8SdRhiCEpWfWJtVNQkj
nMwhrSDU6hB8NrQvhsJbrSeAe5X/dBUHXMkgNg0WtGJb+8RQ+ouJOvFDbv3FfDZy
sxo1A9qtH/lmt0HnF8PNqzqkF6VxS0JakGAUAf9calxBzWQBsdTD+HOWInVzf/+t
kWacY+EqU79fX+uKbc0nQ6spjv6U+tPoLc4u2fW2FYlVZ8RPJ3KFgLc6hnF/Hf6B
Prjg38j78x4gXViOPh+4OOTPgZP9IBAi+1OMJ3liA2UCrF2954qSywFBubtzHx/M
mdQZB2sEz6lBu5zyV6kfUHDtUUBVQIasExyUv9n+QCQXV/nreW+8ehY6UaMqLyGd
gkCVvF0sB5hwg07ergqgQBJM6pMOwFZeIF79ot4dDq/tOZ5BF1kooee1prDrKeT3
35UjK1cg3eRQSm3KQDVwhx88bUFV/5DlB6EgH00U2dhYMe+NC57ngQFq8PAM+35p
yKa4oNH4svtJd8PxkcuHKXo45j2uJepxR4SBlxrvkNlh/myKtoHxxswRKRfR7sU8
axJTViqcvwsspH/C2UcxjiBsQhsNAio1PewTMebf2VVmbEHfv+cn3khF5me/vS6z
HlWucjgL4dLLqUi9SLbbXPa1MxW1VnF5/5LV19eMfaAIfOUMWKxl8MrM2O41vu2c
iCtyCcv/kPR0oQlZpxdFtPdnhTNYS95EBX7udTMPcGm0AzUajPUhrAZ8QMkmq5VP
j89JvoYEa1KrJyZG5ASbRV1PUKrMdzbE2t1UtaRnZUy2lLWeOZpWut1Z/PFphqFc
K+WcPb0KW/THhPyHUZODwoeIk9OAqQ8DNbs3wS6zKqMpy7jRJsJ4AcgS2cyIVWLM
JmRuDReJ5IqTrKQjLlgK2/kukpYCuphL1h3S5MeOK5lBCmwVg5j2yFcaI2Kjvjot
e2AI04LSZyB1SkxiwBs+I/Z8iLLYm5TBkjnBJpkPpFB7qyQ3jDlJI43ZyYffqHK9
W8VugECWRxPhRxSSyvaqH0kMSVkLTHJUyP3WUYPgm5aP4k0Foh3pgxWGfzqLiGnO
4IOkgk1wSrzpV6bCT2fLe2AD+NOPWXTSPNAUvJz19wRHeyjR/u3C3+X/hr1gjuCZ
4j/Bzg04fR1d41gJzK0EzS23NLNgMdPMw96hQHOUqAigL+u2TRoVwhYAjtJDe1Jl
3yOZX+LkigGMoogiBmJJmITiF5VPYqbFjSfh7KYezV9QDkg6QW6bqKB0sZbX3KAA
6JqAaz+bUWxmWSfdt5DyzNcDx5GmZErAhurU75q1lfoYDsMPz6BFmezO/Dtsgs3t
I3krpvRCnXxhyyad3F8ApInurh3LW3WSfuTAza2C0yUknrvjSVOfhE+Zrp7q23H/
k+XvWdq7ZOmZy1zZhkpTAUooyRWgzP66RD2fyA2AI3/7LhHuQ6tO+RnekKss+buV
QjtPYfGfwMYWfI0eY6iLFC7W/8Wag13ZuGwrduvajhHcD3lisdtHLS8qIzD8qrMT
Dax+Kmd9Me1MkLL17iJkdH3ukHOWwMwRuF0z/xaYY90vvYY9ij0SL+qRGBbVmgph
ZriF/FVgvNk3HPEX2hFGHlMrRS95tCYgQkrogjCAEjBs+jPaJV3Bj9igrHUZk27G
eGqA/FXBWj7Ku+jFORvz76EleXYyYLnxsccm0SElsky7g6f0ZdBzjNziv7cv8//h
bG5pG6p3p9GuYOsVaEJgqpAZYe2skbaWXmkOS9z8QDc7W2q+gHmXOU/nb92f96/2
HIAmkJOaYXUZxD6yAQpTu0/+/PMA8keXHtRkPfDX7pKOXhhTC1GyE+KVs0Y62LHi
lkNqhXuV4XKeRF3ga7Sdd41NGjIdR6wY40FkE3xuts4wnOu4yJoRldr0VRxiSioR
iVVM643tLmLyr4RCIboFkbsRMHkPyvlUmVni5bH4rfJ2CQ+vjJE5eY0tGLvmhSrn
28eu8PiA+OrIDlno0sPqCVij/LJP5NIzrJJujtPVqZuuACcrwvwhciadkFbZcV6H
IUa72WSyrrmaB2qDHIPpfiQXY9UAhtMDa9xYGZ9Qu9kXkmEURE3ZWy6zU72gbRF3
TMhoDlBt90Wjl/gahdrYkTdJNR/VNJXTy6ekKaWNHIDkRopXKnQY4nbUncmJmUbE
F0/7US25rZQ2V/OmbvQQBKOn3oNOidth4LzDKMevVhxUdMNrGbMVay66aRiVc6zI
x1Pd6sHVWszJgC16a8QsOfkEHp4+lo1WDnmU42lnnAKTTuR1xFckHPQMIxTm4fwd
r17XQ2eesTiWBE5FM0fxN308LD/NO4AyKlYOygpwh8dVa15NdYhDxplVn0wWcAnc
uumufsS4nN+gM6sZut2Njah2iq2hNv/YLQZvyBG5FbTHkShOIPJN3ThOom3Z9nbY
nvqCefF3D11aGX95ML00iiLWHfHi682908RbvheTM0u4Dz3NH4+TsRC7NgIZ4pLW
UMrvxoPR5NhVQGlW/fpPeAo6YPHqceuh8zFxfEuYC//shwSgqo7EUh2fXIqV844a
Va4ricaX1CDz11PSjg290tJK5UIvvG8/a8FEb67pTUSIn1gK14BD58XaLyNEI+mk
HVW/i6TkN9txGibhYPzj6aJq07tieaJeMNZcSjU/6a8A7BJGKgJNW6coBzSADO/n
F2i9K707TfYcFoPlgzgbXiR4I2pGeecqQORrJxwb1G6G0/5rtV7nDo91+QQZRMXG
ckdIhMUcFigJpDLR88bbYg+DHlO+aDIbhGl7fwoAmoO4S5Z0Bx8PY/h/wKOR70aV
VHWHF8/7j69Ab6tSMFmhMkzzU8EjcBDKz3Cr0cl1Xbq+StunusZbnImGwxhk/sHP
AwTna4uw6Hr9lE9bEFBx+iElUl7PYAXaqk0VqhjTaOmKu3A77B08w+nr/zfY0w7+
2A8yM3a1+bsenlykwtwTXUd5sW+zYmgTVsD41X2dp6EaCIw+Bww/9MAS47cVfnkT
UC8Hz21xkZTec7EmpyfjlNeGtNY4vOSDD0xCkHXp9SNPqURa9lz7s4J6pkcEwqR/
k155NOX/9mObm19FYwSZmjpO1/xAEOzigcr0VyYAd1OTxqRmFb6cqBNzwgVNsks5
m03wqQlieedgQWC2MmzNWDn7oHViQHVDVYSZmQgnSuIFSINbhEpcqF70n2+dDDBY
Cm3tYRLpHBsQJWKFGIsvQ2m/ljqVFfiNoBW2JD7BFCfGC2q3o61IvaZShzQRdyTi
/Qt+kV0WjLCdji8xgttYsVB08ttyN3bY2TmJWjtcCQBC8QCHfZxup7Pn3CYYvG8b
h56nTaT+dzZc223eS0dMdFTAGWVE4Nq+zbKCNDRSamOlvu9bl+my5fy5dlaNXTEL
PIkQJA8/1/C1LZup3KRwRkMN009oKWGYmf1AtMYysIlXDS/XAsopiEXzu9mudATx
6ochjd92yl//JPfRWoGMNmyK1vhKsMLJ6pvUR0gS56Hjf32p5Bytkpbqj8QhWm0i
3HSxBpKUWKcIsuX4IRxM9bpPuhVZDJQrS84klON3aE04t/7xPcktJFmV2ZVTLkEb
K4QQpPoMAxeEyHyTPS2AcsSJUbaECQudzQpYit588VvYHdcCN/9ZQNkzy0LvWVgD
xAKXnVJMrEuskRiuG/RpIJj4Re2fW8pBRBtH29UOgKKfycLKFumVdCIP8OMjF3ky
BEhVRp9Ix0tHws6OjFdm0fumgj5f7LJpPIkuyOumGpunsvT3mr0Rk/K7krYw3DAy
o3IcoKBg2AHZOSZKAJhhfTPZjQ3pfX3s9ZgCTx04qK0v+5G1B6Q5ZWdl1DCylDB9
LSMW3M/9ljhFTPb+rolH4+yVucErOa4AQrX1dUy2z0X/S2N9MzRWgNXRx/jq3raL
60rbnQNiiJgIXOMFtDxIFSVjWapZDlH/TVmzHimS9Et7mhoMB6MUKaJe+nbOpFs+
3xtGaZb91eZQq1d1tX/166FKOAukh5cKdGZvceTgv3trEgxhGqfXkjIhKa7da/k6
EtnzeNI/mWIacMJs1lJA/RhDOmq3GzODke62Vy4SLu2fFDeA42f/Evx7NVPbWqpe
Qvrtii5TP2E63AoMeG3WwxKKeWouaiUrR5V7p9k+cz2qP9GMaKsJMVtysD7lWlz4
gi2ldKHLo0C+5Wr+Yxz48n8Cz9dAyXnKHmJ/a5WQ1bf3K9R4YoKrqh8XZjdBMONK
XvxqBLDJWpmV/jTZ4E7nYKUemk/uViCqnc3yOE3UNI/QCuJQOMqbhQmScpBocXh+
4FDb1MDhUJNOYW18om38X/JlUkMKn6tujV3on+fUqRze8CoRos2GTBLEur3zrR6a
AH1HzxlWGKz0ImypcgENjKUffs610o/Rd/wE2cKMFmkAfPhDs2D3syPzbk8z88o9
G8x3bEl5feixFJd0xvE6kWtFRUJ7IwQvTwrnJxCZR+8rV0/18dv9uYWtylJGFdbW
RdalT2InkyngjkAoPyrlYC9+C4WdHoAD0bR0mCzj0oE5F9fNhBTJEpMT9Vj9s1GO
tw60Cmm5Fe3obluVbhD0JAUIP0tq6wVo049Pr/fsc2PF4t61eCie7y6QslGZdOlJ
mjF8t19NHMT7tTlYyIe1cMwaMr2TyjfqjcPme1XwgoWdLti+5ubMLpzxpoGzlQWp
Gutl+hQC1CPCXvcmAaVVwSgwfwvB2/8wnJZ/WQw0jFGGJEBSPvRWt2wiKnrGe/rw
Xr6ZoV/Xg1UuEM9DdGGGyi1tpRIPLxGkTD7kNY2SGGuQowzsR14jKU/82gIpIN33
9hgirKM9IV+9RUt0RTEOQLld6jW2IZgYMfsNOblmZ5zisEr58ythLr7EdsXTvCW+
7oN/uCWK8iYNMu4tziZOb51xz6F6/QbmfC4lajIUjWmKGwTARIrQk0gzGQbhNwZb
lZibuO5/ADbjxJNXswIVaCRyAGVTMzZzaLWPQu2NrafdyLrajCaUTC0LpMSO3GmK
Vh9uH8GnwN2M1QtXiyNkVo6INP3MJ/oxLiJ0E1WXjyjYMcDPP0lyan7ymBZ3oWFz
4Ywriy8+dEQ0oCQtwmiJejkHlAqaVdKBdLlyWwmxKZPk7TGTR8vb4zany638nwbH
eBdhjPd+ZeYSrkNYA8R+U/0jVmvXHvsnbOOFrpS2IgJ3FPot72XK+L/GzHjd9/td
80lfccj8eRjYTwJmb5Fc0Fnl7yFkLFlEiaXT1IqBKuo2BfifekewlOeOnZlxdLug
xBrwXhePbCZ6M5jnqYDVSMYOVhRNo45v1uFNp4oRaWVj/TUndsU3Nyry131a0ArB
QFQ5zyBqG3jzW1YpdHMgx/Tn+iJgFTBNUGDJnxw81nFVmxSnMH7w1uas3yaXq8kf
jfjR4bXpjGLUrFQQe+wybPRuqfVSJAhsMRbn3d1dM3VLpxUcndsa6HkjxooCL0Jm
/MMyE1rNBVShwlYu8ycC58r+HvV5H6rz22rTvB05JRgI28+rPNle51iD4IZDKK5B
BF19nFBv0jiockDfK6498ng78obi2fEgSM3ILSmfOEGbpxAZdMz00HLY1PBJP/XJ
pP9b78goZtBtDw1bNT7n37pkdjQZmslYIBjDmJOZ+U/D4hpgfYY/o6fkxsUaXD+b
VyYiVURFCNsmA8nfipdk0rGB7hx1vHvTRCjfKIL8e7qhtlYgwyaobRKQRTGm4v3I
jFKecHXOasIXD7O2MNEclqqb+5zj9Q/qouOhV4firVH8GNQYf5UmZXfRkn5g28Fs
3Rf2jI8NQITQrcJ8GAvmsUI4esZdIjSEQw4nzXGRK5FWeaGc7syJewjrrU/NVBsF
Tqz2IuuuUMi2ArtI0hCsZDlrFi3zZK7br2WHMliiwRIliBityIWvU/4vMDlozDQY
jWJ294MsL+7o99UhCUbJWDqB1wBDD01TM4ButuS3+GrZ4bHkqJepbHsSsqLO6Gk7
kxI0NEQPUA1pf+GQ8utCWTB0ugD3MFlsoD8WvJvBj/a7oYLryexVZD4DqWPluKlS
AV/0Vv5LVKdxao49V+EEN1nLJfay6uLpLRG5UGz9d+khr7QGMbynsYPxQ/S+QZsm
c9IH/bSoEsGIULMQnvQYOE4f8uZnD+KfiAPsAMH9oWlvjIeFfX+4LbfgtYRDKTub
uK/uv0iwLQInTb3hOYr3JAgiXXkwQzjtMNllcFtLUAbAPOO/vG9GsMtOLexS9csx
tts1Wr14FxDVKpnuK6W9CiIerW2B/RvnHcHdjpIPLRconuAALA+CNMhHsg0BSqRE
sm6u6EpKpSwEJTgWylvBpfGoK+TnRniDr3XWOFEiWGLp2J5Uhsgoac6qUOzLPcqm
7mYuUEsJ6EgvvUPmUO8A02jfPbvA1cCSKOgY1a+7QJaPR+mMX8HcCYuu8zJjwjUO
bVhidWOi6nc/ksBqRJq0iqtiUvhKECWJcGzjPb47lj0MWbvSs1Fy1effVXNMGlEy
ASZx8NQ6Oq4r9l10X5ea4KIhG6FjBw7yuy/yb1dE4o84k/fh2I1Rca58+dpf7X2/
V4bKpW7zv4++kmlmBNs1QeJpPO4b4ZMceLtNGQx7CSUe2cAe5oKExsA4EVvHBcpA
ei7ucbyf6Y1nnvGJL8tK+HueadK85Waf8srEyMeQBlVpaa3i2MjLxnXh3VkYCBAX
d5UOBb8GGdzbGlcycnxKnV3YrH6Mdb2k17bFeg/aWlsno91+4vbcwLvflpflGOeR
F2bi1wS9+mAhW5xVrENnGUaWtbdVqc6yWPzz/2RlvPOt6vsxb0px0j9IJYYqMgDi
IL87S5xSCf15uYTV4lwcS/zJ6Px8DdpzzGkrOLEMmLCx792KmWewnlo7MOU5aYMG
zsIYTClPwtrrOyxJiYLbucmLlBSR2M73s+QzkSaKVfZrD2vbBk1oa3UkPb49CoT+
JI2H+F9SH6vJe4ekNIJEJbWeJL0LZksmsBJqLxD1qRFB6AJzvntUUiI4atBHzOVn
md+YicMyHxr12TBAHz6GxomxXeUYH3j98Xyfa2NdeXqTjOkz9VfdMtZvrDU0Mtj2
pLWBf3mkClbBZG3M+hN0pbcQp9DgPPkA4RnUZHWBQCyh9bbPADZA9ydEy5QjrNQc
wBrVHoOjKzJqQFo2qr08gkFORkPG7wHFGyk5uncag/CQZhWtpdRhzE/kxqjPVxMb
IPGDkX8jGbnj6najRpeT30SgqZUsu+mL3tAgTYZYEv0KGly/bWnC20zVkI5ZRsXQ
hp+GhrRkPPuKOw4RONx40fpIVaa1O7iXMGJi/Ya4HxODWlEhBO8d+ALoi8kFl4pX
Vlj0513pIZ6k9dptTYQy+uXXz2HuxazW/e+0QGi7jFcLPOwc6qTcB8vTXPblu5yi
OFPVqnF3iGlfWiC9uXuDikA14YmzmE1rd0umz/TRjwMypoIm07C3iXCETEc5oz86
QJBMt+C7C19JiRsm7+Eo4lIJGy/0c5qf8SpLNqutuIPGX1SZF3BxpEEdlSogBaAj
kFwud2DhHc9xKYA0ku94ET2HCeXk1Wv2cLJTRRay66IVI4J2Losm7mCwsIcaHtvQ
UB6+osFTN+KrKagdH7+7SLzUYZFHLSW9q9Mh+5w2ze8zWNVzRTh32U9Uq8BMTcAO
PM79tDTfD+RBizkxknB4mkbpzrwm+7FxUOyLp9uHj/YhuC3w4uOKYZ2Z+2RoedoD
ksq6fMAf3xoIIp+Z+eI9i6J0ymlGrXpGusJucB3Vg0l/nHmeI3Td/Es/C2ngxTlP
tC6P0g7jXwYXobH66/CwuLbbp6nmfq4TUa7ynZiR+Vnt6iJqOf/upCoBf5264Moy
3d6miOh+kwFFTtYU09HPHm98E0HfjRRylKma2BYT63Rek7oA9djrLZCbX76o105T
YEvEPHE7kpd8w559RYLKnoQ6OKDjP66/lTpxb48cykSyKwWCVDazZd7E8KcrBDV1
zU/EAYLMrQDszhyGYf6yfqWBndsRJsBWhlzaRORTcBT4CylnE+3pi2bdnZFQQJbS
eVyifU4H9ypGjf7B72JgGw8yRppTaOIkhsnLBFX8MBOQDl9zRvj7R9bqqNrdVtIi
PlCbVdKY0m2mbbBfnLZlF6oW6c3xSUNnf1ehdXKL6OizM1WxppRRaU1plXXRhYyI
evGt2Pxgo+BjNFu7kIA2+BrjJy8uc/0vvp0BIc+uRA0zhTrWy9+dEXTyg6+8LfSx
KElN3ixuojHy6wAPLspQC1AsCH1vbbqbUQVM1QTZYAZu0jD7S8YOeE3W1cfFWTmz
rFtPNkig9e9ceitCn52aG474IvX3dIcTzbSTGdr+kGuzKEljT3HXUVVpWoV7PqO0
hK/fUWKdvKeMEfa1w3SlZNAC7wGYMvcgLPj/GqyrC0kADinkpBJR1NPTdGJIcvU7
onVXo8/CH642zN08LWjTUkuaoZqTqPnyClYw6zCvwBM1PW0gAVqlPLXGMtMdb7zR
ojHPLdpOatMLdCrLj3bl9mAftJuteouxW6CJUAa5rdFLzZWhgZ0lw9+ZFE6xxyjM
gy8aJzeXGeAlCcNELbzSZfUAdj5y3I/G5aw0NcagmLW7NcO7kfpY7eI/2+0tNKjU
H9geQTZrT3VFanqV2B6F676bnr4Ib/giAxy3oru26genNA2ZDA3NksS1xjuwXasw
88tmeZJ3BzFHd9mjXWJOeWfw5kRUDbDP2FNUtuCsmGuA7cP8a2o6hkuApv3+WayO
oGmVrL6e02p4kvl9uC286yLj+0fcC5V+s8wJ9zp1R5qWAtp5s4JqEds1tClw322i
T5USp/J249Wp2lQbKgXCzQg/rjIVA5mJsZj9JZfTm0uBPFSvQ7/Gn0WI/+3nxw2i
YzZVx3H2Hz+/vqQoEq/WlrUFr22b0/IKtH4mqrr4qBtgMiLwFkZKjbAsSLxkO2Br
Hr5WoT41HEm7aCJ+6f3JCTxNA6CiRtoRYteLKIRN8knjezrYu3dFsnLtOSEHkLmA
YTIsizkrzSqlgKOvbIxKpDqKwJXuXK8t0UwDNjFqjXjDK7q+5ITOzsqRYo/E1Ngp
tTCsb94GVKut1uUloPvluwPkoDRxmyskSEGyf3eh5Ovjcaecb6D2dbto4TTaSvSo
PXD7pc2iwueXTj72GTl8uTyk/HRABPh6s/AeprFOkhj82S/V/DVlgHsDqT6US4fI
ZQIgq13nn+E2daVfIxsp+vi/36g4sXgbXwRHB7NlU8ylDg0e9BAUKb695Rz/ulMn
7fDQPO7SXjz1oPIILuDDi8oNxqzUxtel8iruazb3YubOunpubigxErXni72Rm4gH
gRfaeb8Aj5uvUTwZcAGEzKp/PUYNYhb1Ls7NlubkpjwA+/pCrPF7nGobIUy71tF2
j0FacYMu1fVUj+Tyyvm6liftq4dXqSTINKpDqnV3VJJgQQBU0nPmt95/CMnAy7+9
k8Qk7O4+AeseUaneeRbfqIkWcqPE43CC28ZT81ez9S7ihlk7UAUCZyvEWaB92cAC
mpz4QBGf+AWvHHAiADOGlGztl4vgsfR89imFAOltrXcGQ6UxvHFmK3Uh4d5Qrdu3
r01Fcd6pt6P8ZTsMJK+t9hAh3c8ZtzMGC01Lsbtx53U9Mw2UK5CBHgNjPrf33YbK
geycjm6i3L66wOkHMUQGk0ndKIYatrEJ+U30TgeIStHpe6vzIl5q3SUiMJy0mbI2
4atSqAcRxnTjt3msVDIsx7gA9sJQedIqqRc93AIXjy0jtdtV44aHaKR0HDA38Uav
1aeHSPzbp5PL0lI748lYCFRbzD44rSrkozRXoiCcOdJlH6zI1/IaCWlJn+2rrej0
JLscPQbwnFhYFFl0nPyorpMiIrOd37WFz1C4gX6arukJpxOEwvsbrZlwu+7hbzRl
BkPEKxxwvXnoK7OOwiCX868qXmwADQwA7YrJsTLoRBHL0VadZ88L7wffzOs/LGhl
/PL0s3vXHqibN3dqFjni4tARUq6n/VDR8HbNHUWUT8aW7iWKZmk77+xqWLafCkoi
fNjEh0Q7YA2s3YOOCIYoR2mlcyqB9Q4cIN3EW4g56J/3OUeM4T9BAdTLAPFf51SW
ZBswUhXxlJJvB1gWCL72VpsdZ1Srpo7Rsfv82s3bRUk9kDYpf+B2y5ZGQM2X2i0d
BrGFNdUmrxJhJmhoYeRpqTQLZoQiZLTpmTUZ63Bymz911W1ku3FTmolOTQNxW2A3
7sue4idvF8ngaBHSqe2XFo+sUmeWbQVBr3mlZ5KK/OqVj7RTmLWKvVry09kGmjep
8mImuZLihH5Pv/EpHX4Z2Mwx2zFZMMZAjZ5lOus1fy6VOJ+vTaY7NT432E50Z2Eu
wiNCtp9h//s6n7KRE5D4w6f9GD3yKR5uWSQuzEwlhB8jCoVZT6tYdDWncxAsZdA4
tnYmPMuF4AuuaDI+z8yilmHR/xFcOFx+1Ri5zH+zDllRLJzm5xziYDOKEIvp5H4Z
I2XsGa1OqR+tOQ78QrrXzJxzbaKd/+Zdvr/HsP+xG8aRUFVveVSEtsCfLp6mT7EG
5rFeXlpXXeah9w1Jasz76WXIuQRG3sjC4pzxKDq0SkuUVCekOWOa1bil8rNQDfN4
5eXLoOyJs4ZuOnuwmdPyl87x4pqYslUNa/YxFRfShDy4KCGzD5s+F8I/E4U24MVw
Xl6rUjiDSJfiLlSdbxySUzLT1qeQr3V1tlP4HWXqlbxPbTMlT3gMRT7xhHWeGbgA
pb2aUuuiiCqffgK2JREri1PNYj/bQd/2zb5nzaAvpGtxLHFGX79XeMB39UyMaHLt
960x4yNbh5J8xf4V1r0ZdfVpxxeDnhBAkxVOKiPVX4tXd1Hm97FHdNUGjq2QnXNy
69z5csjpyM6tzmpRj2P7gwK3kOhmoQxkc/5tQhGJ8t0BGRO/o+6I6LYhNIb/EPS0
yVBhj9wJ/1a7X1HJpceOt5Pu4ToRELSdA6+kYmlKOBFVlTvZrDzP9Ei6uNPaDp8l
aj1zHUlKcR+hAY1grmH9rBBWE1Y80EUzOA+sSil/yKBxOH3LX8+wHpqFeqsX0zSv
Y4GikCvBm9X+qUtWZoBxHpXPPmjcGqCAqlusyHJ91LgaXUEN8d/aexMpdce6PNzv
Jg5abD5FAKuXhasAv/l43uFG9KFLOwGrkfpekYYCPWRDNSsnA+58ia8mjNB4K6CK
FUE5ObBHY7pLKPFi97gRvemVbyqw95f1s7f+1Zb4Ji2cxzFHS1udLu81Tz6bGt2f
XaW2UrusyWOratEEZsrNcaRB97cF7s9ubf9e+O88amsaUBRr8COLESQUUbqBy/ls
PL/VPyiS0Tzu1ZFRgp4XDy3gVESEIC6lATiErfpzjF9UBNZI7rp70KQwQSohGHTU
kQWqJrPLRVh+ZMlEVPCP7gOm9vyoJdZNISyPySBnCkjUjCSvKfQWO1PgaQjEq3b9
HyuWu58+hbdmBi32QzwG5IzZN1i4RISiWurWhK7s680LMxl4LuZ8S83VNf8WPEQ4
HgZpDLcesF52I9eLRR5EUx6GGORcwotZarw72bPd5tARpwYCUP4qgacrrbloADvZ
f83eub6zarPiK2XSk9TdiwIXKmer9tdoMmQN1EEBFrgExzIFTJx1+XGY/FXn3VGL
tJOdakpq/L+/PIFMqLYnEUWbF0grEmxXdgUHA1xAIs2QM7fTeHNQ2rlfzL1NueSS
3YB91QQUDJRfzznsQPzVb5ycO2olR8yZfRZCAgyVvNaPov+FmZ28Ifr7e4yvxWJy
jK1HRMkcGYaJmqXvmBD837VFiSvBKsRNl15Wx0V2dOzkrSe/KFJbrY0j7+mPQjG5
abx81UtfyIEFZXNYEbZ+F62+3cyqc+LffJsf82pDHWFxuapn2r12Epicr8rCeVFm
N63ly931JZ/jA5niNYnxhJdsJ1LPY5tKLX6Iri/fZE56HWftl0pTOTUy1c/ZceNo
zgoTrB0qiYLp0UxGWu3PkAG2LrcCbStUuLPFxkQwvA02XMUZab4lsB5jCdCz7QEb
0/48IoozPyb7sAqtT3++FvUj1WfNpsSDT2qBeJsfI95KI0xC40eQANfH3tiGEtJZ
KyT2u4Lb8Gfx4yrY7FDKxdiiK5maZfCKvo4v0qokhT+xVDmvY/XZB8XjKuheMaaR
VyL38mYzOzoG2oJ2rzVM5X3LJgCtCsJuAmbHlDtfYyWyzMEAxtT88cO6ZWPQhNVd
SSS2OaOTqHvuELAmDk7dcwm9htRlDWmBviCBKjhKwHXmEz0XfMQLtV0owm4gy+QE
1+pSiKOTVHmwQb6f/g3IGBzIAVJ9zbcp2MsOZLK1A33FPfrpekd6zGIgpkT56685
ExtWrQlAulJKPOHvh8qdpMfBE/VTyZ5HoK6jwcrN3YjWciLIYnIMpc6aT85tJNlK
i3MEQ3P1k+Qe0Fd+bBdUkkPr1hOfvdtDiXyQqDugLzOLgzjO+7n4HudH3qog1eMg
wAkBxDcCRxmgB/FdkEAcoaLDiFX1E3yjm3cAy4lXv6OHmfffw7U5cRHYVxD9+E2s
GOeryWWnHLDvezHBxLySee8afNE5juwG2z45xlT689HLisiy0nj58uQHCLJcm8JP
yVnDmQz9XJspyEXq5nvaVrEbvNEXwz42lF4udDnna6H8FvA1cu+h8F/nX0TyP4Bx
anDa/Cz+Vx2Fqy42iNWyppOzZgGfJOyzNCBsb3qiujh52yBGACwmhyLQq3wM7SNZ
xe3pN0JzQGRPXMG87ee50s95AJTyq0cxkqQM/pJcpHVtX1wYQTEyB/WCdzwWYFqR
y9LWUm3+VCjaQ41vJW5eZt6spmwHZRsJ1HxgmYqLGrWG0fYjoGHsY5fc9VaiWKgr
mc8Zum613xuWtE1r6AA0q/Zahxtw8ZR7tGWDkVHT7/2Ida48CbwMi/br7oUHQjmz
lGCHEUHQqzxH4Qcb43nuPyzNO+qfbhWPoKAdZfpS2CxyHy4l75Az68qCIsAkNzR+
hsYi4QhuhArIiT9R3EADsKxF8mZFVK0JOz7uMXWGmyxKz3pLObQNHLTXMHpxUMov
pkwX21TjnV5aNeP4U4Bfmtzg39m80bOwqL+l4HmF95Vlaad4OtSHj8ML4+p/T1zB
p4tmqc8ZRe90WQ2HxS6dowyeE/ycWY2A0cxODMZimI0KOiYJWd0j+4FynTI5cwor
YxrZN67Y6+gcvUshWwUq0uZ4zdMQ5rdHrxw1n/jtH6NmTVNFNuvi9sRmn3oAcJ+C
dif01oW4wp3uUsGsxCIkzUE8DVxaQ+vXOz1o9RPhDrJMK2IN1vXWxVAQTohIKN66
Osi0uk7Xlxg4Ulwb5cJcCV5tt9OcCc6770JBpkFJcTS3Pe09qGjy+3eihzxD341I
XhjZYlJTfp33i/NQCYkk8RfypRUAQ26y4W0IIdERO37SbooKak4j8HnwI1TYx8O2
SoxZiJ5gUMcVTqdvMP0ip+vuGci4XFE6UB1upwAQ7TBICTcbvTxTyoTIYD7ay62l
L90TtbpqA5YcVQRiZImpKbKZFRjVvZeuipLfpq7x8Nt6qy/vvRA5yJgzQuqzydqD
2UuW2cYka1EbPAlYisnxO6ZFoxQoIafzNMwU0BBymXxxfsPPxRaQyY4XFX4TTZXt
7Fk9La2Oz6sixTIVOyKYlcFTImYp5k4T1J6IV4/7OEL4cToGDIUzExHdY2CZq1eW
l5Wmri/l8/1jxXnEZcKAMNlpAW+f2+wzSrrpPNDxa1LQ5eVYr+4ejebQl/5O4rVH
Ftt5tVXAfOcbzXMM84Em7sf6qSHRQk0v+C12fM25AS7YVqQZkQTq+xvEITyFl61k
8AJ7nlcOuxbYtiHsqeWTY7lrlooHZiCyMX0cLT5qnpj3rAJ1+vzs6Kcn5Iw23gji
x0SwVmlLPhdO8AEa8H3azwXSG2+3/L3LFhsf4mfyKUEQfFrmN6CAGs/Z2eg6ztdA
7F1V+wjmate6QsByxZ1ZavkHkcf2WqWv48hgzTNVK4w1fYRrkzruHJTmQ+0wjZ/Q
DRqg3ZNKOMc2EFuNK1lWGiAPe/AAglGVu/dnvZiOdwWykUPskQrx5pu9LZGDvSO6
CZx2s5Ge96Z2hBbJKz6HVY0wW8QgwdCmtWTgCLRfItbxlLMxdsxic66FyRJ10afu
MmvaTUJkDJydnfgXEKwbstoSNPiz0VVjA9lpWYtN+eV7b1/S37omvHPjsVWDWJMc
xgPjHQxCi0BhaQr8/bW0B1LLZL5CIl+I1tlglx3fBvwd2zPehRd8eM14Ot0bWi2I
e3XzFTTaO/7SehVvpj3ScsbnOarxH5CR1aWSXpVIXDN4yczKMvG4rGFybuuPLyYV
jubX5W2cpiQCvW3ERuB/acwph/WiRALpaz7TamatdoJQx5UDcn7cdUm1d3dq43m6
v3sLJ+EBt9T+vZ73EC43vKax48LTYUolnqNl2f6OJY/3RoWHFG7kQiB4Mj378AFd
CuNFFVW6MGWx3i1V0XbwYKBO2PhB5RL0n0tJeRn6N4RUF4hS3Gh9Mkz/5/iZ8ZP+
+uFzG7ZPyAJLKoH75VaVNDQbXvXm6wEWmq/aR9web+NXY/forxHnJnSchZrUIK+O
F7uugAEbax3k+IvKN/LJN90bCilFybxHHydUB4GH1YLzUS0bb7n4WSUrb9J3aQei
iPxfvhlfpHcbkzVl97ZJJiilkSyGt5D2BOL+6fnMMnGDQr6xnol3auBETToNVEjS
KmdUlY4HjNzb06fIgalfcpKNc6NZgH8dUCGHd5HUF8JQ0DF/6Kp0YjlblX2rqT+j
PpREtrza6GeZLoh9LMp0gevtkZ7KbqCk81rQ4vi/hOPo8ufthsOyvfcHL9maOpC0
ase5WNFkUazfMDCau3UIYBYp/0NJ97j4U3SIYRSBVze6cTU1UWjEVcBioi2AcTun
0OTuiZowsZeamJf1VYy6SbpuhKLuC3EZVMbqypXotojqZZb3ZnsOrFgFRjsCTe4s
EnwHTD28k9wvXtV/a3np2zH/SekyeO8SsArUS14di2Tn8boVW545XkDwIOZXZalS
hfxp1mW374EJ0YS6305Ovb2LVCSC8qpla3L0tB2HeeJ79IsMo+EMr5RIV35MJN0R
bufCdEaEPg08QEXrz7R6/guqxS/kSIOWh/2H7mKF3fQJd5rWv7WS9L79h5yVrDv0
LrhVfhBhAIOQn03Jpb6QFQzxjLfqOTJqWtGpBl4vhg/CbAGefUFotiAGGyVloEyq
Zu1as9BPAv1Z18GBBLryNgBRz8AXZr8b5rsy6+D0RIA173KfpL2E7laQQ/g7wjaK
s2uNoMjJw4mQ842VFnJ2Y0COiFyXeEcm71wycNlCaBxfyymMTLZ3Hlor7Wct7o5f
CSaoWD1hbQYJvetiEAwTb8V+gDUq8xcCcvkuE7tOnDrbwynX5IqwZPxtRTUVpo9o
w4NSFgNxwtY2sBpHitvep+lUEshqz3VMdVkO14B9DChjT0gk3gkY3ZQVLAPphzUh
qMHUXc5h+3G1XlJVbxzyvnl2H+0f6nzhpqQagI0Oy3LzG676UjVk2nDecHQtIAm6
cjoGhsjd25O6qLFBmAyPFyoJLWVniHABAQDx2v7tnKZthQpZBkLU0h0/vz3dpzSk
pLP7coI5qEirNJkVZKqW4YXXRc8ViqhZMytC+HuW/HSyWvmmQlzqa5oJVUHiGsQQ
e7Wj82S9r1e/0BURlVPP82rTsFbDlDQsSK2TLshoN/jFj1O2PC6vnbjDjV9QSlqu
sPvkI65bD+aHUiFCvlsENX6lNuvuXN+Z2IF9+rgPYhh46JC0cQ6ayLdST6aZe4AT
4ea5G/9WzZwaG7WfeUwSzjmkA9hHRT1AA3V5KOLH+BUkswewu2vBcYx1noCTnvvp
LYLyvH85+fd8FbIHy3oGxHqaMKNI4kq6hlAUoTumv485bYLCtMsIHPmLZXlgS4W1
ncArDqmvkjtftPo1GZuiakslreGoL7GfOJ4B2AlC+O28cmEaV+hTm4LlsmVSDjl7
FNii1nBISW4rV9BtirXm6zS+u7efypUJFiERtxPn3FLOedNPJAxCiwXunNOLv4o3
vucJWNsvDshjTMKzztUNCPY57wDanmgD7x3/+je2tyZNUTbPfSjTsTXqTYQRPhDw
1yda0Ds1QuUe7OGVuI3NCQSZUNYfOZMP1I1S21KRQQA+/ku5dQfQz4niKyLWHspC
lwtaB5ROXW9RmFnbg12rFwTsz1FdAhD44ZEau5dq7rYF+FvNvzY5g1Z+DveS00Su
bXvLixEsUa5ddFg/gs9h/pQ3F4w6e6kvYuxHHdW3N1cIKLzntrQyFjdvnqYz85dV
xwwmVvJbiXENijWjuEM1x7ICvugLw6T0t6B253RapoBG+h43Nkzxp+zsOWB0I0Ds
eU32aYIy5X5zLZaDYiVlk1oC4GDL46QvepPSSoLG1+ugLNSnkxoFxI0N1h/OW5s+
d0UnLI2UYLcYicPEpXPKCwNUh3dFJMgIQjFwWioI/DDLbJ0pdmRdd/w5Vo23niE9
IKaJrySnxdpBMXDUd7mQU6YkXTBRydq5Zr9T1CEG/Qu7nw53Di+K0wYLO/TuY4Va
1tw7nqi4X4tccQXd9OUvypOErk+/6oYVsmmP4oGlXWKp6MIJCC5M9GUYD8i3SO/g
div2OtcBKQQTOkEt/wSsqBy40Q39Id6tlR4FuUN9UCaMIX2ljVj7wmliueP7n4zY
Sp/S71nPw8uzSuIGTWuT8MFwKVJ2Wa0C08EaSQap3wu3mjyzA+w8W61oF2kFb4Lq
O3C8fx6/On9tRgYHjD44wpfcI5ItD92csNZI1C6HZQBqfYdq40MicVGe9KYh10P6
qEpZOoD2Gmxdz7f92DpIaY0TVbZJIkjawP+ubUwF1w7ZW6xd9/X23/7BQpo8CvQJ
9avJUkQLdk4dgSebLMBeqV/oLDvrt8ppXxffAAZDAU9/jTnzlPBK+dTVZKYTiqxb
UiQJA999rDsw6R/hzGBBgm1EJ/F/r20XH83oKdbFFCB/p3H9ibeP7fY+aHyUAwYW
w6i6JTC1a3axAxv4RmMGSFXQtmlDM8oPSsvwqNr7JFGcHolJCYD/K1NcMZw7o/4w
AlbyUQrvtRem+1NbH2VbF1PMjHFfZeoJ9Cv6eC3Hb+Zawl9EUUUXXWUKo+Ldn+7M
q20CAtVxHWkOmB5BjJwAuMIKoJziLSa6CvDTxj++ao247z3wBhlgLmrlFE0S/loz
6gm6Ic1vOBEzadK6dDsYmw8pzd0+ZIdO/16TgJqUv/1JUYjWZ5F2hQsprsKZmGkd
p3S9q3QThgHT+QIxwLZcznHNnUgOIeIXhaaG0jFV4OUi9qSa51fbsTbn6F2zxAg5
RiMYhnsGJfNUdWVTzIWRdDSJI5w7WIflqt70Var+EgYF9jiSbU8RJt4IICq1iPwv
T+Om4zx6/Ixgp5Kj95Egsh6SienTLU5DzNM8gNfulp8vIa6K+hMR/MXa1M2EfUKI
t4qkcW3OYXaK3tWL9D2jSwqYgPWMizozM9sMKiZ4Cm99szvDh6rTTeBDjz3e4N0x
5ArdWDTiiojT2gWaMwPc7T5W1niiiNje6DqZrGQ20RyXaQor1SYw2MHSfdhs1nou
C7ZLZaCUj7fWlMp2t3qIwUSxI/Pa2gSV/zoTr3Aqlnzwc31ZhGhbatRZ964kyS8F
qPazHQxxFll7/AR0Rd+JsLmQ5mW2vtfh2YlSIlvmKrWI2kHAmhvo5BnLPiqnPxaa
J8iTnasRdeMgrGMeJuwlJ4r8YhSepm3A+G1cQucaOgeFrlN9/Z16LL+mSpZ9MEmH
PUDr8KnwYweSgKNczSAoyGZU0pb7KTYJpuXKYS13bUBCs1vNfDKPyyIEfMslESXu
5IdGSbxz1HVyv5/OtvXbVET2wKF8rtUgqb+fj8wQdHTwbS7fQv2EWVL4vwQ6CGU+
AhRbJU1TD922FD/cdm4QOzVpWlI2P83QG8zycu1Hh+2FJB0qFjjXfwtyskqW1Waw
c4X0Ec2gjgAUQ6iLJ0/DoBPEqzCygt1PWa6j/ShAiwUvL8FZvrkbuEeReZo1gC1d
gwSZ0a6OynN7jr63qyMmGKP3PbCu/1/aQAlweGp3tSmp4G11J0mP882zgoW8uG5W
O7TvxGpb1P5xv0I43tubznuEBMKP3atdH10IHqH8F+3ILW4BLADRWdS5PcYQzO8x
E4RPqZQFTGV1VkGIZqo18qXQhPGG67A1MqKhrPI0LbvGiGpj7FEywNR2Kcm/SW1q
+mCLisY8BlAnFx/SxYG5XqRcQxwJ0azovA4BTe5An8tDdcgBbkMKLH08uF9k//Hm
g2ObpLEs5F+Oz4Lz5v3yIfWyvrmJ0KZaaGE1Ca86O1T7U88/IUxgLAyB7j8+t/Bv
IVIzsxQcYtGmttjazmr1Ok2NmGCr9v0TciyrU2IsSQxta//kQMDYMsiE/wUOmnbm
5Php9naFVhBtoc/ZVzmhLHjKq5yO++LQq6qwRp0ZKddyTidL/E4Fo3jFzqWr+bjx
YlfR5dy/CsPfor7hm1mrupDLOFnQ7pOcGL1LsKY5vK/5fnHTWoj7PucARiML/Wm5
bauFvuDIiOwgCwob+ipYHyIf3bTmucRkhP1WumtQFCLc6BQgXK+Ty7XFgpOq0wIs
SysdLf2AUjNAs+EmtqEwzjBnaKVYNF+aIHTD5wlyyznNCF79eTLiPfJp31YnPwQg
PbKfA7gJ1F86WvA5y5fhEk3nqqhMEiqP01xnEhQcMHbRQQMz8Z8SrF8Ibn/EuXx/
aAlshaz+0PU4mzajVhrt0PDSRWjolXBHTcFVh462T+rXjNDHvVxXPEfoEK+9716d
DbZKqKQPN5Yv0FAdJ1Gm+rC6cTwuMG4Hsgq6v/LS+uq6JgAHY9v56+sbWcqDr0Ei
q5eDs7u7NPiYHDATqoL0Gu5HLqy5DgWskWGAgnp4wrhvuF3bYc7KMyvBNibRQ277
+rQgdrMn0thIIQTFaXHP/mAkNli6bsXqSDDDLTL/42TntbeFKOISznddi/qPg1e/
nzomaf51Tse70iUmVCr1Z28kRjVVurgY+a4lwKw7kKVPFqpqP0LTrBTkCfa+c5Zb
QE/m6vpgHVMTEgGaNJxHCH5j1XQUvpCDB5Kza+hHnsbuIjXbOUjFVG5IrLwQwA3U
Y2tF/Ii4tIoAka7VnHMogP4vBBngCREBAqeSDrCXSBFhuZLkm/DlemHGqzmyUdgV
7NXR7YsHmL+Y+8BULRm3dCGcSGXdTwfdO6PzOTr0MAlzXH6MKzI/3Z2nIHK2UEGU
h7+f16DgvimggV3bLrb198t/4qydHNfOvSychbM0+fl/KLnRTHW6Dex1NXENyTrc
ACAOuY9gFTGorCNtvYhp7NUDS95RY7JDajNc/jQAsBRnLz3mA9iBVxhJfNzfdKYj
djdACuGq5Q1OCRBybBPf3e7HRo+ioUp545mufNX/5zek/m0o0plCQw5nNBlwS3QQ
TZwJg6du7KlbNKIkWifDm7t4VTQEAkqT3AbNr3s9Ipf7TmnssmrCh0ZDVyVT/Cfz
f59muff05po6409u8vgpKVoacr1okTjlDynOQkXoJZSA7p0rIu+Bp5RQ63QYn27V
pIWIZtBFcdkBTfAvhEDSXHAKmEnP7jhhrGWCVt8LQ8pYifNEQZ6dyABkR8Sep2Tu
2lbCHN6hFp+tV0vNGv9xr6BwBumuUKSAstCry7SuJ98JHp+o+DIojCsw+A3xDtMw
BWSB68mE2/EJeadUmIILFoNe0o65e3vX5Ns4gXLxSXqUBbT8mV2MPD+IQbd+bzxt
E5LTRsKeiaFqpBLMUuGXhhe7rW9flSad4KrJytMQyp/7rD+BCXWSXLSf5McApfgB
egzJ2yqwa7qxCtq/Vyl0PMAD5EySYhNYfifc1llVy/ecQ9xT9IxSZgdFih3yepKw
GNe/DdHG7VBB9AuXgIi9MCFskx5+IAYBdoVhBY1OzCf0heT9cvE06tKtHX23kS33
G4576jN7icxLHrpPnaOk18hc5A6z/bKAFVzWhm5l1f41+Ju2XwXMHJgYXJ5DODBi
LqUmGMuvLq6oxmfRyMK+0TXEc1hcNB8bQ41G09bSSVqisxqEt77MN5uZFaAIcpPi
bkGllB1Yh3w3dBOFOOUA9EVw8sGk44QbGRkRUe7E+PSTz2GRJPhMOyLCVQEFdUT1
R8qUJ0mulTljzzZNdEibuPwlENObKlqCQ8tYyemrNaoBbvwc8IF5P2pyDUc+i9Ck
iTZsGjLFWTF5q+P8d2gjyyJeS2/LDWu0VrWtZvrXsgWAFiAtqEVRmy5GAllD+MNi
dnRpbYkR4nUktz88GMegWV3s3p7+m7XNIpgtP4/xYKmz/6n8LX/7ixC02nXJH2Mc
lgBno8+WOnkfUoSdTsSekTn0uIIHgwVHDQRKrpII/XSidvuT3LxbgmKrRQtc08W3
4Gy4ukjBbsdUfBTE1NJGUFsrJyrSV+09uOimQVPskfC+x8VRTqXn48f6jWNUpLnE
xfpeIG80JaxUsce2KjJLKdyNPgvkKIrZ+qH/uNcOVLBzVul+MnU5LwOkSkPm2DFV
5JExTLMnPrFypFWM64B47+5SKBp79Q0fsJtdI97+ELJBfphlPZcy4Qp5BvibqNvn
ZW3wZlVSffi/EgLyzv9hqnlSPPvv8sbb9p7cSSqMJzr4CTJjjZ65V2Vj8kpauNPE
DRENhvy1H8HJMcYlmMhbUrLuyXHf/h1y2UepFC51ugL0HpAf+XUqSVUwzL828lVc
XKhHaTfiuBYEBmA/4ybuzFn/qhvqpgqt072HkaWrpOLdIBJ6ugvV4NDS80T7zly0
fAJF7v0hPSvDUQ6M9dHZmQBs2oUJ66eWyueYHdb4CQoarYWJa2mWFUpfrHVa1D4T
azpuxBpU07Okanm3hFFEidFEteg7H7kWa6oIxBVDc9dX5kCpywke9D2TbOvi22kH
lIpUjhgEz6WwiRpYh7sOg6OnyyPFMttbP3jvoZTqItMWcrO2GC/bpty2fOKyoy3Z
dk9Kkpa8VTWVno3lFUhUioRvdN797UHK6X1AGV9iSJDr8/mHBH1zCvuUJdrYvDRX
ORUbVKnKS5RpIBO+iPnQuPQfj8x5okn7pFJY7p2jEA/nThpjLPe3ucO9s8i+TRuR
qLmXuUISRQn0GBIjgXzGYZfuNYsvcbOGF/fde1zNozwRmOCz14+N0uU18Ntkia+T
J8r6DN2sG6axWT/CR2bs8N4blqrr/LJEDYs6AN8Z+vQed8pJ8pLj4bzWW0cjbPmt
b5/Edg2Qmob0RxY9hrzYlfVeKj8EgGsEl/7+lmbWNbGSr2Og6dH/03HPiZY9GCtO
Y8TeatklMdtO1OUvy/x3WNPwXnV5bDg4HZ+IbCPEQZG2oSZQ4sd+B9bgOlNjclUn
`protect END_PROTECTED
