`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tHUfsWA7hq9wMdvRJTOpT7yHPLwiGGS2mHgMRvz8H5H2Wmba0FT7ko1u3shAXHZY
rjv+eCZYrqHgAslY2wlYkftgnjxImpbWXxXpvoQ4dWGP59vkf99MricQFwG+qw1T
s3B+dk5fB5quce3+VqOdZ8WxUdf5NkKkOKjW7wemk3oXMj8eEYfIJCgVrjg45hPW
7Z4nWUVpR7VBUikfxhfWL4f6BG4toPdhxLHbJP9Z5yN44dlWP1Y88dhvfuPDXUAq
OLlUwXAbKyVUzQux54f8XMraDCW+5qW+iylhX33izDw992qQGM22J4YeqfltNzNj
zzCjjh0039xa0WyfD4NQzx2JJ89vHEtp1sdr7FieGMAHcMjI1FckZD/8lAtaYpkL
qVLa6TuY/y7/FufP+Ocpl5uV0ZOe/cK/7O3rxMnwNM7rybIQEjFGTJydoN6B2TKO
owkX8Daf7+60wZLir+tKos1xFKx6HRt0Kpq2cw/QOvjmCh/uoVujpMiQVT7I83z+
dCdTEf5ufKmv6+bRi7eeKg5hyAZj8GI51YarcwDtCOhFaXDvlw8he+C0SAG6jxrh
C3Kf6g8v3jtgcuhHZiFbtqTAKuvCrA/aE5k8hCuBZUrXHwe9EK2RlitpRkQp2LUu
bsie/tQP2SYS+KzCLeMh/XUfZ/iWYSpApBfRhXPEGqU0h0Bx6VjFZgZrjrimzEUQ
/q/frtc9ouLviQyjz5waIlDas9J8C/reqwCFvtqlqkTB649Eq13QvOnXp2fGjpVN
eYlSsc8xifNkONj/89vgBoYzMkpRGTON4tPPg2D0t0JwRMEKtAeW+SQPb43DRCdP
fVxYayErEps2uIxx1D3BLFxKWjwp34m7/FQAVWfU2hVbav1uDAxCWJkpa1uKigsC
KO8OWItggyg96QMUP9i9BvtvKdJPyJokmkBpKS46/wE1yyZwEIzT0esc5thM8sPw
040aNNaj+O0dk+0izFrhX3x2J6unNolsTRBChJIklbD68wWYyd5dz9ISq9WEc206
nf5cUyenpKH2+sOTmNM8/72hjoBJVBcGZTsN5cd1sehzZ7uYr0Lnt9TGpJTQL8m6
k7lJLz4VPxO/P3v9Pqwn+dgrcVRgjWJbMitr5hHwzZNey4klHs/Uwno3CiEurkb5
zjMxeD77wsS8YdyrjM9CX9MSADrBeFTULyAQv7anVhSsTpHQQ15Fp+LCsMiHEXM5
JiYySo7xxx4jkagYQhqp2LLt0Y13fA9IpSBTzxV1T6Oeh5p+UiJyBYkxNeo2gJ3p
e3W1sGfNsh6SB7Y2e3NK0e1hUXpOB01x5AxdV3Zhxb6FHGaW4aZf0d2h6subzQbn
DJjplujmV9n0DdpFkcbz9qKwcs3sB0iz3VnH84EC5tKLVBRJuJSlk23NfiXksvck
uod/F5hjvnddife3IHLS7++udCRbJ/lEFFFB7pPS9WRmodPXgBWSHS2Pm858xJE4
r4WU2b0hBW/tqUfTSsENkoOSVhZ8oT8Zc05uchvoAqOu7Nbdh0xU+MZzhQnBSXkU
2+8GxucOBbbJBLvXEzKOpWOOmTbqmjvv5YyWY6dUGbkX/lWUkrne/i+JRpCcOCJO
d7aVOFz6wjbDQUsCATsfMdw9Zp4GiOSyQLZ8iiihQyXNWVUnNtZAU5xKBaPXw+rz
A6aCpG00GRiP77nFgQjZjEbrY8Fn+JqHKPvq1oK5v6B0GcZy3a1RIOuSU2/4aJ5l
QjmXuX5cDQ8F2GFZrcdAcI0wEBrg7d2lynP8ZaL3CxqnkKcxoIZjNWKrI3Gf0cxK
mcC2jtCZgci4Hqo246J7WpxEapFeNTAHMoLeAsleI+zc00Vnc1bEzpC+2hasRzlh
O+a7KbpXuoCZLKrKYG3N7XKVrfrVvmBdgHnwRafeHh9pHwfRQYV6xNyGdmmdL5Ql
0aZLFI/I4cpn1ebXWbBJLhuVDR2XD0Z6kpvY/gKIlrGKju6sUbTwxpuvXF8I89Ak
YuChRPkp3SSfDWs0EAYOe0SlXEAkWFNl4qyUD1aYxd7NLg7yuVel+A+ZmYAslhO8
vWb0SyNDstfwdhJlL8zTGPTCt1IK4NJzoC4gX5RP1AWdiBGJOkApLt/xsPqeucFq
sX2uAG5sSAhtwdw5idPqqv2r4om0kBF55dWs8h4blUjr/RYzyZ01UEjcutX60Xn+
P3bpTBoiRki/sKnmbZMBTw/QlBHA+rQEtwt3+ubVxfAmaWOIXeX6KqrlBLe5XDmO
LQjBMSSGuO8sICNKFl2MU9siK3WurLJ6mZx6al+KL6RPhF/L92868Rfo4vVCjYdd
SIl2IXIrDawuv4CEGH8x/mp7buAoXn6eolHW9gp4fFu4gsL5onsRBWhNiv5oN8IG
m2F9+xnq9/2NO6+m2HAaaOiEMF4POopTtuKPaeQDU5gI1t3tBmflANOGAoGvQxUX
Kz4v7V66zz/RguR75cB6l1QT3fJweUfBITwKbqbnthzoEvWq72zLeyzVeYKo2x12
OVTm6g6v8HpCkFfvkU6922HpHGP2J6xGePEl/n4kwKyBSruLNfU5+lnDbPc2x+AZ
pJ/Jj5Ywmd6WWE8rQmPFbIaqGsmoGxeiVA1M35Aq92n5r7FYd/6VXSwgIduz2hUC
kR09QH2dfjtxNR2hnxSRB5jFvDVI4iwjjLlcS0TPKjeEQ6d+jx+c0m2G3Io+5z0Q
c8Vr85rOXSbGlI4qje8g6puJW2ZNmZ1HpcnGEWvrR68+YoYsYmWjuYPE5FESnxOV
pZpBrL+ZKsct9+kCPe8MJJnH9TlhWVCdwTVNnA87m4upC6pgfkvs7Y8ynPMLOqo2
dV1VYmGfPPwDwH6ULFgs29yw0CXHHWf27XtlkzoC0b/T7Wz8mjTBXxgiHVQambUB
nrQ9ugsgZd2K24ovCs9qz01o0Ch8ntjhjCoS5XEPjwXn1+llMJamvAOV+1uEDL+p
eSzDS/0CSKTg5X4LtxPJRuiO8xfcssQ2z8m16lSxcVscc0fPvm5h552+Kv6QTktZ
SKTQ86jFQJDZVbjnIqHX6PMN7brC52QK2lUJzr3q6KEwtqRiVXTl7CW1JR9D3h0y
Mach5cZ/jDIdB7ximNOURw4M5/5cKqjbR1n0SPwB8fs3wnd01Olb7cHnKD2dE9YV
ud6EDfnrgFGwRTwl+K8sa02IuvujF3gVClmcU7jRwcso3pFZ30Y5rwQCydszsp6U
DBrpi2KLkq+8yeiAnWJt4NOcWyTWqL5W1T8LWFZQa36+lajiOf0JvRHQHckfQGBf
/aApNSvPpe5BKHp6T8kjfe+VGBIv8TiuuL9sjwaeIBDXa4vk+aIUt6mjTzcYsF1v
VzWibQwJw4UAWgUNb2dDwQKiWqpGM9vVYgYVg9fgNzN1bvKCjQ4DKjeCTEKrSNrI
NF4KBHRbnkv52tEdSRzVB4rMkst+L0giGtUPMqPglKK9h9uGed1P3ySex9AWwWZM
E6KP8QAiROanHYRmmkiKmoa0CVpxqtheGh6Zy/FYrNt9p/LGzlph+ARN8VI0o/88
j4V0hCzdTR3G0jtw63Fsf6d3p9MTxMrsnatZkYml78w2UiapztZWB6rGP4iAEtoP
VXKHNlDikDeW0O79ntesM7VFACRLzY0/AuZbyGt6IYNSEfiKvSaLLaCwpXVL7cMs
o+oQ3AbNwjKdLKUkD38qU0QXeyVJYGiRrP0jtu6QoY/EyoqLCcO8xuTZNUwWTG+h
duVbEzK9Ra167Pi34mFcGQ==
`protect END_PROTECTED
